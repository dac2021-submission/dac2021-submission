module IBuf( // @[:freechips.rocketchip.system.DefaultRV32Config.fir@215163.2]
  output        io_imem_ready, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@215166.4]
  input         io_imem_valid, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@215166.4]
  input  [4:0]  io_imem_bits_btb_entry, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@215166.4]
  input  [7:0]  io_imem_bits_btb_bht_history, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@215166.4]
  input  [31:0] io_imem_bits_pc, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@215166.4]
  input  [31:0] io_imem_bits_data, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@215166.4]
  input         io_imem_bits_xcpt_pf_inst, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@215166.4]
  input         io_imem_bits_xcpt_ae_inst, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@215166.4]
  input         io_imem_bits_replay, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@215166.4]
  output [31:0] io_pc, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@215166.4]
  output [4:0]  io_btb_resp_entry, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@215166.4]
  output [7:0]  io_btb_resp_bht_history, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@215166.4]
  input         io_inst_0_ready, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@215166.4]
  output        io_inst_0_valid, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@215166.4]
  output        io_inst_0_bits_xcpt0_pf_inst, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@215166.4]
  output        io_inst_0_bits_xcpt0_ae_inst, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@215166.4]
  output        io_inst_0_bits_replay, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@215166.4]
  output [31:0] io_inst_0_bits_inst_bits, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@215166.4]
  output [4:0]  io_inst_0_bits_inst_rd, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@215166.4]
  output [4:0]  io_inst_0_bits_inst_rs1, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@215166.4]
  output [4:0]  io_inst_0_bits_inst_rs2, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@215166.4]
  output [4:0]  io_inst_0_bits_inst_rs3, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@215166.4]
  output [31:0] io_inst_0_bits_raw // @[:freechips.rocketchip.system.DefaultRV32Config.fir@215166.4]
);
  wire [31:0] RVCExpander_io_in; // @[IBuf.scala 86:21:freechips.rocketchip.system.DefaultRV32Config.fir@215247.4]
  wire [31:0] RVCExpander_io_out_bits; // @[IBuf.scala 86:21:freechips.rocketchip.system.DefaultRV32Config.fir@215247.4]
  wire [4:0] RVCExpander_io_out_rd; // @[IBuf.scala 86:21:freechips.rocketchip.system.DefaultRV32Config.fir@215247.4]
  wire [4:0] RVCExpander_io_out_rs1; // @[IBuf.scala 86:21:freechips.rocketchip.system.DefaultRV32Config.fir@215247.4]
  wire [4:0] RVCExpander_io_out_rs2; // @[IBuf.scala 86:21:freechips.rocketchip.system.DefaultRV32Config.fir@215247.4]
  wire [4:0] RVCExpander_io_out_rs3; // @[IBuf.scala 86:21:freechips.rocketchip.system.DefaultRV32Config.fir@215247.4]
  wire [1:0] nIC; // @[IBuf.scala 41:88:freechips.rocketchip.system.DefaultRV32Config.fir@215179.4]
  wire  nICReady; // @[IBuf.scala 42:25:freechips.rocketchip.system.DefaultRV32Config.fir@215181.4]
  wire [1:0] _T_4; // @[IBuf.scala 43:19:freechips.rocketchip.system.DefaultRV32Config.fir@215182.4]
  wire [2:0] _T_5; // @[IBuf.scala 43:49:freechips.rocketchip.system.DefaultRV32Config.fir@215183.4]
  wire [1:0] nValid; // @[IBuf.scala 43:49:freechips.rocketchip.system.DefaultRV32Config.fir@215184.4]
  wire [1:0] _GEN_1; // @[IBuf.scala 44:73:freechips.rocketchip.system.DefaultRV32Config.fir@215187.4]
  wire  _T_8; // @[IBuf.scala 44:73:freechips.rocketchip.system.DefaultRV32Config.fir@215187.4]
  wire [1:0] _T_10; // @[IBuf.scala 44:92:freechips.rocketchip.system.DefaultRV32Config.fir@215189.4]
  wire  _T_11; // @[IBuf.scala 44:85:freechips.rocketchip.system.DefaultRV32Config.fir@215190.4]
  wire  _T_12; // @[IBuf.scala 44:80:freechips.rocketchip.system.DefaultRV32Config.fir@215191.4]
  wire [63:0] _T_19; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@215200.4]
  wire [127:0] _T_22; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@215203.4]
  wire [5:0] _T_23; // @[IBuf.scala 121:19:freechips.rocketchip.system.DefaultRV32Config.fir@215204.4]
  wire [190:0] _GEN_3; // @[IBuf.scala 121:10:freechips.rocketchip.system.DefaultRV32Config.fir@215205.4]
  wire [190:0] _T_24; // @[IBuf.scala 121:10:freechips.rocketchip.system.DefaultRV32Config.fir@215205.4]
  wire [3:0] _T_31; // @[OneHot.scala 58:35:freechips.rocketchip.system.DefaultRV32Config.fir@215215.4]
  wire [3:0] _T_33; // @[IBuf.scala 74:33:freechips.rocketchip.system.DefaultRV32Config.fir@215217.4]
  wire  valid; // @[IBuf.scala 74:37:freechips.rocketchip.system.DefaultRV32Config.fir@215218.4]
  wire [1:0] _T_39; // @[IBuf.scala 78:63:freechips.rocketchip.system.DefaultRV32Config.fir@215228.4]
  wire [1:0] ic_replay; // @[IBuf.scala 78:35:freechips.rocketchip.system.DefaultRV32Config.fir@215229.4]
  RVCExpander RVCExpander ( // @[IBuf.scala 86:21:freechips.rocketchip.system.DefaultRV32Config.fir@215247.4]
    .io_in(RVCExpander_io_in),
    .io_out_bits(RVCExpander_io_out_bits),
    .io_out_rd(RVCExpander_io_out_rd),
    .io_out_rs1(RVCExpander_io_out_rs1),
    .io_out_rs2(RVCExpander_io_out_rs2),
    .io_out_rs3(RVCExpander_io_out_rs3)
  );
  assign nIC = 2'h1 - 2'h0; // @[IBuf.scala 41:88:freechips.rocketchip.system.DefaultRV32Config.fir@215179.4]
  assign nICReady = 1'h1 - 1'h0; // @[IBuf.scala 42:25:freechips.rocketchip.system.DefaultRV32Config.fir@215181.4]
  assign _T_4 = io_imem_valid ? nIC : 2'h0; // @[IBuf.scala 43:19:freechips.rocketchip.system.DefaultRV32Config.fir@215182.4]
  assign _T_5 = {{1'd0}, _T_4}; // @[IBuf.scala 43:49:freechips.rocketchip.system.DefaultRV32Config.fir@215183.4]
  assign nValid = _T_5[1:0]; // @[IBuf.scala 43:49:freechips.rocketchip.system.DefaultRV32Config.fir@215184.4]
  assign _GEN_1 = {{1'd0}, nICReady}; // @[IBuf.scala 44:73:freechips.rocketchip.system.DefaultRV32Config.fir@215187.4]
  assign _T_8 = _GEN_1 >= nIC; // @[IBuf.scala 44:73:freechips.rocketchip.system.DefaultRV32Config.fir@215187.4]
  assign _T_10 = nIC - _GEN_1; // @[IBuf.scala 44:92:freechips.rocketchip.system.DefaultRV32Config.fir@215189.4]
  assign _T_11 = 2'h0 >= _T_10; // @[IBuf.scala 44:85:freechips.rocketchip.system.DefaultRV32Config.fir@215190.4]
  assign _T_12 = _T_8 | _T_11; // @[IBuf.scala 44:80:freechips.rocketchip.system.DefaultRV32Config.fir@215191.4]
  assign _T_19 = {io_imem_bits_data,io_imem_bits_data}; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@215200.4]
  assign _T_22 = {_T_19[63:32],_T_19[63:32],io_imem_bits_data,io_imem_bits_data}; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@215203.4]
  assign _T_23 = {nICReady, 5'h0}; // @[IBuf.scala 121:19:freechips.rocketchip.system.DefaultRV32Config.fir@215204.4]
  assign _GEN_3 = {{63'd0}, _T_22}; // @[IBuf.scala 121:10:freechips.rocketchip.system.DefaultRV32Config.fir@215205.4]
  assign _T_24 = _GEN_3 << _T_23; // @[IBuf.scala 121:10:freechips.rocketchip.system.DefaultRV32Config.fir@215205.4]
  assign _T_31 = 4'h1 << nValid; // @[OneHot.scala 58:35:freechips.rocketchip.system.DefaultRV32Config.fir@215215.4]
  assign _T_33 = _T_31 - 4'h1; // @[IBuf.scala 74:33:freechips.rocketchip.system.DefaultRV32Config.fir@215217.4]
  assign valid = _T_33[0]; // @[IBuf.scala 74:37:freechips.rocketchip.system.DefaultRV32Config.fir@215218.4]
  assign _T_39 = {{1'd0}, valid}; // @[IBuf.scala 78:63:freechips.rocketchip.system.DefaultRV32Config.fir@215228.4]
  assign ic_replay = io_imem_bits_replay ? _T_39 : 2'h0; // @[IBuf.scala 78:35:freechips.rocketchip.system.DefaultRV32Config.fir@215229.4]
  assign io_imem_ready = io_inst_0_ready & _T_12; // @[IBuf.scala 44:17:freechips.rocketchip.system.DefaultRV32Config.fir@215193.4]
  assign io_pc = io_imem_bits_pc; // @[IBuf.scala 82:9:freechips.rocketchip.system.DefaultRV32Config.fir@215246.4]
  assign io_btb_resp_entry = io_imem_bits_btb_entry; // @[IBuf.scala 81:15:freechips.rocketchip.system.DefaultRV32Config.fir@215243.4]
  assign io_btb_resp_bht_history = io_imem_bits_btb_bht_history; // @[IBuf.scala 81:15:freechips.rocketchip.system.DefaultRV32Config.fir@215243.4]
  assign io_inst_0_valid = _T_33[0]; // @[IBuf.scala 107:24:freechips.rocketchip.system.DefaultRV32Config.fir@215259.4]
  assign io_inst_0_bits_xcpt0_pf_inst = io_imem_bits_xcpt_pf_inst; // @[IBuf.scala 108:29:freechips.rocketchip.system.DefaultRV32Config.fir@215260.4]
  assign io_inst_0_bits_xcpt0_ae_inst = io_imem_bits_xcpt_ae_inst; // @[IBuf.scala 108:29:freechips.rocketchip.system.DefaultRV32Config.fir@215260.4]
  assign io_inst_0_bits_replay = ic_replay[0]; // @[IBuf.scala 110:30:freechips.rocketchip.system.DefaultRV32Config.fir@215267.4]
  assign io_inst_0_bits_inst_bits = RVCExpander_io_out_bits; // @[IBuf.scala 88:26:freechips.rocketchip.system.DefaultRV32Config.fir@215252.4]
  assign io_inst_0_bits_inst_rd = RVCExpander_io_out_rd; // @[IBuf.scala 88:26:freechips.rocketchip.system.DefaultRV32Config.fir@215252.4]
  assign io_inst_0_bits_inst_rs1 = RVCExpander_io_out_rs1; // @[IBuf.scala 88:26:freechips.rocketchip.system.DefaultRV32Config.fir@215252.4]
  assign io_inst_0_bits_inst_rs2 = RVCExpander_io_out_rs2; // @[IBuf.scala 88:26:freechips.rocketchip.system.DefaultRV32Config.fir@215252.4]
  assign io_inst_0_bits_inst_rs3 = RVCExpander_io_out_rs3; // @[IBuf.scala 88:26:freechips.rocketchip.system.DefaultRV32Config.fir@215252.4]
  assign io_inst_0_bits_raw = _T_24[95:64]; // @[IBuf.scala 89:25:freechips.rocketchip.system.DefaultRV32Config.fir@215253.4]
  assign RVCExpander_io_in = _T_24[95:64]; // @[IBuf.scala 87:15:freechips.rocketchip.system.DefaultRV32Config.fir@215251.4]
endmodule
