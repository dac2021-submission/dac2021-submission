module TLXbar( // @[:freechips.rocketchip.system.DefaultRV32Config.fir@4792.2]
  input         clock, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@4793.4]
  input         reset, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@4794.4]
  output        auto_in_1_a_ready, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@4795.4]
  input         auto_in_1_a_valid, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@4795.4]
  input  [2:0]  auto_in_1_a_bits_opcode, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@4795.4]
  input  [2:0]  auto_in_1_a_bits_param, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@4795.4]
  input  [3:0]  auto_in_1_a_bits_size, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@4795.4]
  input  [1:0]  auto_in_1_a_bits_source, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@4795.4]
  input  [31:0] auto_in_1_a_bits_address, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@4795.4]
  input  [3:0]  auto_in_1_a_bits_mask, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@4795.4]
  input  [31:0] auto_in_1_a_bits_data, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@4795.4]
  input         auto_in_1_a_bits_corrupt, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@4795.4]
  input         auto_in_1_b_ready, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@4795.4]
  output        auto_in_1_b_valid, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@4795.4]
  output [1:0]  auto_in_1_b_bits_param, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@4795.4]
  output [31:0] auto_in_1_b_bits_address, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@4795.4]
  output        auto_in_1_c_ready, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@4795.4]
  input         auto_in_1_c_valid, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@4795.4]
  input  [2:0]  auto_in_1_c_bits_opcode, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@4795.4]
  input  [2:0]  auto_in_1_c_bits_param, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@4795.4]
  input  [3:0]  auto_in_1_c_bits_size, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@4795.4]
  input  [1:0]  auto_in_1_c_bits_source, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@4795.4]
  input  [31:0] auto_in_1_c_bits_address, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@4795.4]
  input  [31:0] auto_in_1_c_bits_data, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@4795.4]
  input         auto_in_1_c_bits_corrupt, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@4795.4]
  input         auto_in_1_d_ready, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@4795.4]
  output        auto_in_1_d_valid, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@4795.4]
  output [2:0]  auto_in_1_d_bits_opcode, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@4795.4]
  output [1:0]  auto_in_1_d_bits_param, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@4795.4]
  output [3:0]  auto_in_1_d_bits_size, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@4795.4]
  output [1:0]  auto_in_1_d_bits_source, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@4795.4]
  output [1:0]  auto_in_1_d_bits_sink, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@4795.4]
  output        auto_in_1_d_bits_denied, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@4795.4]
  output [31:0] auto_in_1_d_bits_data, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@4795.4]
  output        auto_in_1_d_bits_corrupt, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@4795.4]
  input         auto_in_1_e_valid, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@4795.4]
  input  [1:0]  auto_in_1_e_bits_sink, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@4795.4]
  output        auto_in_0_a_ready, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@4795.4]
  input         auto_in_0_a_valid, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@4795.4]
  input  [2:0]  auto_in_0_a_bits_opcode, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@4795.4]
  input  [2:0]  auto_in_0_a_bits_param, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@4795.4]
  input  [3:0]  auto_in_0_a_bits_size, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@4795.4]
  input  [3:0]  auto_in_0_a_bits_source, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@4795.4]
  input  [31:0] auto_in_0_a_bits_address, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@4795.4]
  input         auto_in_0_a_bits_user_amba_prot_bufferable, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@4795.4]
  input         auto_in_0_a_bits_user_amba_prot_modifiable, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@4795.4]
  input         auto_in_0_a_bits_user_amba_prot_readalloc, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@4795.4]
  input         auto_in_0_a_bits_user_amba_prot_writealloc, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@4795.4]
  input         auto_in_0_a_bits_user_amba_prot_privileged, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@4795.4]
  input         auto_in_0_a_bits_user_amba_prot_secure, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@4795.4]
  input         auto_in_0_a_bits_user_amba_prot_fetch, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@4795.4]
  input  [3:0]  auto_in_0_a_bits_mask, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@4795.4]
  input  [31:0] auto_in_0_a_bits_data, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@4795.4]
  input         auto_in_0_a_bits_corrupt, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@4795.4]
  input         auto_in_0_d_ready, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@4795.4]
  output        auto_in_0_d_valid, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@4795.4]
  output [2:0]  auto_in_0_d_bits_opcode, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@4795.4]
  output [1:0]  auto_in_0_d_bits_param, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@4795.4]
  output [3:0]  auto_in_0_d_bits_size, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@4795.4]
  output [3:0]  auto_in_0_d_bits_source, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@4795.4]
  output [1:0]  auto_in_0_d_bits_sink, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@4795.4]
  output        auto_in_0_d_bits_denied, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@4795.4]
  output [31:0] auto_in_0_d_bits_data, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@4795.4]
  output        auto_in_0_d_bits_corrupt, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@4795.4]
  input         auto_out_2_a_ready, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@4795.4]
  output        auto_out_2_a_valid, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@4795.4]
  output [2:0]  auto_out_2_a_bits_opcode, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@4795.4]
  output [2:0]  auto_out_2_a_bits_param, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@4795.4]
  output [3:0]  auto_out_2_a_bits_size, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@4795.4]
  output [4:0]  auto_out_2_a_bits_source, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@4795.4]
  output [30:0] auto_out_2_a_bits_address, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@4795.4]
  output        auto_out_2_a_bits_user_amba_prot_bufferable, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@4795.4]
  output        auto_out_2_a_bits_user_amba_prot_modifiable, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@4795.4]
  output        auto_out_2_a_bits_user_amba_prot_readalloc, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@4795.4]
  output        auto_out_2_a_bits_user_amba_prot_writealloc, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@4795.4]
  output        auto_out_2_a_bits_user_amba_prot_privileged, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@4795.4]
  output        auto_out_2_a_bits_user_amba_prot_secure, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@4795.4]
  output        auto_out_2_a_bits_user_amba_prot_fetch, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@4795.4]
  output [3:0]  auto_out_2_a_bits_mask, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@4795.4]
  output [31:0] auto_out_2_a_bits_data, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@4795.4]
  output        auto_out_2_a_bits_corrupt, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@4795.4]
  output        auto_out_2_d_ready, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@4795.4]
  input         auto_out_2_d_valid, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@4795.4]
  input  [2:0]  auto_out_2_d_bits_opcode, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@4795.4]
  input  [3:0]  auto_out_2_d_bits_size, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@4795.4]
  input  [4:0]  auto_out_2_d_bits_source, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@4795.4]
  input         auto_out_2_d_bits_denied, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@4795.4]
  input  [31:0] auto_out_2_d_bits_data, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@4795.4]
  input         auto_out_2_d_bits_corrupt, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@4795.4]
  input         auto_out_1_a_ready, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@4795.4]
  output        auto_out_1_a_valid, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@4795.4]
  output [2:0]  auto_out_1_a_bits_opcode, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@4795.4]
  output [2:0]  auto_out_1_a_bits_param, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@4795.4]
  output [2:0]  auto_out_1_a_bits_size, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@4795.4]
  output [4:0]  auto_out_1_a_bits_source, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@4795.4]
  output [31:0] auto_out_1_a_bits_address, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@4795.4]
  output        auto_out_1_a_bits_user_amba_prot_bufferable, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@4795.4]
  output        auto_out_1_a_bits_user_amba_prot_modifiable, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@4795.4]
  output        auto_out_1_a_bits_user_amba_prot_readalloc, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@4795.4]
  output        auto_out_1_a_bits_user_amba_prot_writealloc, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@4795.4]
  output        auto_out_1_a_bits_user_amba_prot_privileged, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@4795.4]
  output        auto_out_1_a_bits_user_amba_prot_secure, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@4795.4]
  output        auto_out_1_a_bits_user_amba_prot_fetch, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@4795.4]
  output [3:0]  auto_out_1_a_bits_mask, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@4795.4]
  output [31:0] auto_out_1_a_bits_data, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@4795.4]
  output        auto_out_1_a_bits_corrupt, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@4795.4]
  output        auto_out_1_b_ready, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@4795.4]
  input         auto_out_1_b_valid, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@4795.4]
  input  [1:0]  auto_out_1_b_bits_param, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@4795.4]
  input  [31:0] auto_out_1_b_bits_address, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@4795.4]
  input         auto_out_1_c_ready, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@4795.4]
  output        auto_out_1_c_valid, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@4795.4]
  output [2:0]  auto_out_1_c_bits_opcode, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@4795.4]
  output [2:0]  auto_out_1_c_bits_param, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@4795.4]
  output [2:0]  auto_out_1_c_bits_size, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@4795.4]
  output [4:0]  auto_out_1_c_bits_source, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@4795.4]
  output [31:0] auto_out_1_c_bits_address, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@4795.4]
  output [31:0] auto_out_1_c_bits_data, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@4795.4]
  output        auto_out_1_c_bits_corrupt, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@4795.4]
  output        auto_out_1_d_ready, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@4795.4]
  input         auto_out_1_d_valid, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@4795.4]
  input  [2:0]  auto_out_1_d_bits_opcode, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@4795.4]
  input  [1:0]  auto_out_1_d_bits_param, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@4795.4]
  input  [2:0]  auto_out_1_d_bits_size, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@4795.4]
  input  [4:0]  auto_out_1_d_bits_source, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@4795.4]
  input  [1:0]  auto_out_1_d_bits_sink, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@4795.4]
  input         auto_out_1_d_bits_denied, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@4795.4]
  input  [31:0] auto_out_1_d_bits_data, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@4795.4]
  input         auto_out_1_d_bits_corrupt, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@4795.4]
  output        auto_out_1_e_valid, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@4795.4]
  output [1:0]  auto_out_1_e_bits_sink, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@4795.4]
  input         auto_out_0_a_ready, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@4795.4]
  output        auto_out_0_a_valid, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@4795.4]
  output [2:0]  auto_out_0_a_bits_opcode, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@4795.4]
  output [2:0]  auto_out_0_a_bits_param, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@4795.4]
  output [3:0]  auto_out_0_a_bits_size, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@4795.4]
  output [4:0]  auto_out_0_a_bits_source, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@4795.4]
  output [27:0] auto_out_0_a_bits_address, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@4795.4]
  output [3:0]  auto_out_0_a_bits_mask, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@4795.4]
  output [31:0] auto_out_0_a_bits_data, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@4795.4]
  output        auto_out_0_a_bits_corrupt, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@4795.4]
  output        auto_out_0_d_ready, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@4795.4]
  input         auto_out_0_d_valid, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@4795.4]
  input  [2:0]  auto_out_0_d_bits_opcode, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@4795.4]
  input  [1:0]  auto_out_0_d_bits_param, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@4795.4]
  input  [3:0]  auto_out_0_d_bits_size, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@4795.4]
  input  [4:0]  auto_out_0_d_bits_source, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@4795.4]
  input         auto_out_0_d_bits_sink, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@4795.4]
  input         auto_out_0_d_bits_denied, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@4795.4]
  input  [31:0] auto_out_0_d_bits_data, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@4795.4]
  input         auto_out_0_d_bits_corrupt // @[:freechips.rocketchip.system.DefaultRV32Config.fir@4795.4]
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
`endif // RANDOMIZE_REG_INIT
  wire  TLMonitor_clock; // @[Nodes.scala 25:25:freechips.rocketchip.system.DefaultRV32Config.fir@4804.4]
  wire  TLMonitor_reset; // @[Nodes.scala 25:25:freechips.rocketchip.system.DefaultRV32Config.fir@4804.4]
  wire  TLMonitor_io_in_a_ready; // @[Nodes.scala 25:25:freechips.rocketchip.system.DefaultRV32Config.fir@4804.4]
  wire  TLMonitor_io_in_a_valid; // @[Nodes.scala 25:25:freechips.rocketchip.system.DefaultRV32Config.fir@4804.4]
  wire [2:0] TLMonitor_io_in_a_bits_opcode; // @[Nodes.scala 25:25:freechips.rocketchip.system.DefaultRV32Config.fir@4804.4]
  wire [2:0] TLMonitor_io_in_a_bits_param; // @[Nodes.scala 25:25:freechips.rocketchip.system.DefaultRV32Config.fir@4804.4]
  wire [3:0] TLMonitor_io_in_a_bits_size; // @[Nodes.scala 25:25:freechips.rocketchip.system.DefaultRV32Config.fir@4804.4]
  wire [3:0] TLMonitor_io_in_a_bits_source; // @[Nodes.scala 25:25:freechips.rocketchip.system.DefaultRV32Config.fir@4804.4]
  wire [31:0] TLMonitor_io_in_a_bits_address; // @[Nodes.scala 25:25:freechips.rocketchip.system.DefaultRV32Config.fir@4804.4]
  wire [3:0] TLMonitor_io_in_a_bits_mask; // @[Nodes.scala 25:25:freechips.rocketchip.system.DefaultRV32Config.fir@4804.4]
  wire  TLMonitor_io_in_a_bits_corrupt; // @[Nodes.scala 25:25:freechips.rocketchip.system.DefaultRV32Config.fir@4804.4]
  wire  TLMonitor_io_in_d_ready; // @[Nodes.scala 25:25:freechips.rocketchip.system.DefaultRV32Config.fir@4804.4]
  wire  TLMonitor_io_in_d_valid; // @[Nodes.scala 25:25:freechips.rocketchip.system.DefaultRV32Config.fir@4804.4]
  wire [2:0] TLMonitor_io_in_d_bits_opcode; // @[Nodes.scala 25:25:freechips.rocketchip.system.DefaultRV32Config.fir@4804.4]
  wire [1:0] TLMonitor_io_in_d_bits_param; // @[Nodes.scala 25:25:freechips.rocketchip.system.DefaultRV32Config.fir@4804.4]
  wire [3:0] TLMonitor_io_in_d_bits_size; // @[Nodes.scala 25:25:freechips.rocketchip.system.DefaultRV32Config.fir@4804.4]
  wire [3:0] TLMonitor_io_in_d_bits_source; // @[Nodes.scala 25:25:freechips.rocketchip.system.DefaultRV32Config.fir@4804.4]
  wire [1:0] TLMonitor_io_in_d_bits_sink; // @[Nodes.scala 25:25:freechips.rocketchip.system.DefaultRV32Config.fir@4804.4]
  wire  TLMonitor_io_in_d_bits_denied; // @[Nodes.scala 25:25:freechips.rocketchip.system.DefaultRV32Config.fir@4804.4]
  wire  TLMonitor_io_in_d_bits_corrupt; // @[Nodes.scala 25:25:freechips.rocketchip.system.DefaultRV32Config.fir@4804.4]
  wire  TLMonitor_1_clock; // @[Nodes.scala 25:25:freechips.rocketchip.system.DefaultRV32Config.fir@4834.4]
  wire  TLMonitor_1_reset; // @[Nodes.scala 25:25:freechips.rocketchip.system.DefaultRV32Config.fir@4834.4]
  wire  TLMonitor_1_io_in_a_ready; // @[Nodes.scala 25:25:freechips.rocketchip.system.DefaultRV32Config.fir@4834.4]
  wire  TLMonitor_1_io_in_a_valid; // @[Nodes.scala 25:25:freechips.rocketchip.system.DefaultRV32Config.fir@4834.4]
  wire [2:0] TLMonitor_1_io_in_a_bits_opcode; // @[Nodes.scala 25:25:freechips.rocketchip.system.DefaultRV32Config.fir@4834.4]
  wire [2:0] TLMonitor_1_io_in_a_bits_param; // @[Nodes.scala 25:25:freechips.rocketchip.system.DefaultRV32Config.fir@4834.4]
  wire [3:0] TLMonitor_1_io_in_a_bits_size; // @[Nodes.scala 25:25:freechips.rocketchip.system.DefaultRV32Config.fir@4834.4]
  wire [1:0] TLMonitor_1_io_in_a_bits_source; // @[Nodes.scala 25:25:freechips.rocketchip.system.DefaultRV32Config.fir@4834.4]
  wire [31:0] TLMonitor_1_io_in_a_bits_address; // @[Nodes.scala 25:25:freechips.rocketchip.system.DefaultRV32Config.fir@4834.4]
  wire [3:0] TLMonitor_1_io_in_a_bits_mask; // @[Nodes.scala 25:25:freechips.rocketchip.system.DefaultRV32Config.fir@4834.4]
  wire  TLMonitor_1_io_in_a_bits_corrupt; // @[Nodes.scala 25:25:freechips.rocketchip.system.DefaultRV32Config.fir@4834.4]
  wire  TLMonitor_1_io_in_b_ready; // @[Nodes.scala 25:25:freechips.rocketchip.system.DefaultRV32Config.fir@4834.4]
  wire  TLMonitor_1_io_in_b_valid; // @[Nodes.scala 25:25:freechips.rocketchip.system.DefaultRV32Config.fir@4834.4]
  wire [1:0] TLMonitor_1_io_in_b_bits_param; // @[Nodes.scala 25:25:freechips.rocketchip.system.DefaultRV32Config.fir@4834.4]
  wire [31:0] TLMonitor_1_io_in_b_bits_address; // @[Nodes.scala 25:25:freechips.rocketchip.system.DefaultRV32Config.fir@4834.4]
  wire  TLMonitor_1_io_in_c_ready; // @[Nodes.scala 25:25:freechips.rocketchip.system.DefaultRV32Config.fir@4834.4]
  wire  TLMonitor_1_io_in_c_valid; // @[Nodes.scala 25:25:freechips.rocketchip.system.DefaultRV32Config.fir@4834.4]
  wire [2:0] TLMonitor_1_io_in_c_bits_opcode; // @[Nodes.scala 25:25:freechips.rocketchip.system.DefaultRV32Config.fir@4834.4]
  wire [2:0] TLMonitor_1_io_in_c_bits_param; // @[Nodes.scala 25:25:freechips.rocketchip.system.DefaultRV32Config.fir@4834.4]
  wire [3:0] TLMonitor_1_io_in_c_bits_size; // @[Nodes.scala 25:25:freechips.rocketchip.system.DefaultRV32Config.fir@4834.4]
  wire [1:0] TLMonitor_1_io_in_c_bits_source; // @[Nodes.scala 25:25:freechips.rocketchip.system.DefaultRV32Config.fir@4834.4]
  wire [31:0] TLMonitor_1_io_in_c_bits_address; // @[Nodes.scala 25:25:freechips.rocketchip.system.DefaultRV32Config.fir@4834.4]
  wire  TLMonitor_1_io_in_c_bits_corrupt; // @[Nodes.scala 25:25:freechips.rocketchip.system.DefaultRV32Config.fir@4834.4]
  wire  TLMonitor_1_io_in_d_ready; // @[Nodes.scala 25:25:freechips.rocketchip.system.DefaultRV32Config.fir@4834.4]
  wire  TLMonitor_1_io_in_d_valid; // @[Nodes.scala 25:25:freechips.rocketchip.system.DefaultRV32Config.fir@4834.4]
  wire [2:0] TLMonitor_1_io_in_d_bits_opcode; // @[Nodes.scala 25:25:freechips.rocketchip.system.DefaultRV32Config.fir@4834.4]
  wire [1:0] TLMonitor_1_io_in_d_bits_param; // @[Nodes.scala 25:25:freechips.rocketchip.system.DefaultRV32Config.fir@4834.4]
  wire [3:0] TLMonitor_1_io_in_d_bits_size; // @[Nodes.scala 25:25:freechips.rocketchip.system.DefaultRV32Config.fir@4834.4]
  wire [1:0] TLMonitor_1_io_in_d_bits_source; // @[Nodes.scala 25:25:freechips.rocketchip.system.DefaultRV32Config.fir@4834.4]
  wire [1:0] TLMonitor_1_io_in_d_bits_sink; // @[Nodes.scala 25:25:freechips.rocketchip.system.DefaultRV32Config.fir@4834.4]
  wire  TLMonitor_1_io_in_d_bits_denied; // @[Nodes.scala 25:25:freechips.rocketchip.system.DefaultRV32Config.fir@4834.4]
  wire  TLMonitor_1_io_in_d_bits_corrupt; // @[Nodes.scala 25:25:freechips.rocketchip.system.DefaultRV32Config.fir@4834.4]
  wire  TLMonitor_1_io_in_e_valid; // @[Nodes.scala 25:25:freechips.rocketchip.system.DefaultRV32Config.fir@4834.4]
  wire [1:0] TLMonitor_1_io_in_e_bits_sink; // @[Nodes.scala 25:25:freechips.rocketchip.system.DefaultRV32Config.fir@4834.4]
  reg [9:0] _T_882; // @[Arbiter.scala 78:30:freechips.rocketchip.system.DefaultRV32Config.fir@6856.4]
  wire  _T_883; // @[Arbiter.scala 79:28:freechips.rocketchip.system.DefaultRV32Config.fir@6857.4]
  wire  _T_180; // @[Parameters.scala 55:32:freechips.rocketchip.system.DefaultRV32Config.fir@5462.4]
  wire  _T_383; // @[Xbar.scala 173:40:freechips.rocketchip.system.DefaultRV32Config.fir@5931.4]
  wire  _T_164; // @[Parameters.scala 55:32:freechips.rocketchip.system.DefaultRV32Config.fir@5446.4]
  wire  _T_374; // @[Xbar.scala 173:40:freechips.rocketchip.system.DefaultRV32Config.fir@5902.4]
  wire  _T_148; // @[Parameters.scala 55:32:freechips.rocketchip.system.DefaultRV32Config.fir@5430.4]
  wire  _T_365; // @[Xbar.scala 173:40:freechips.rocketchip.system.DefaultRV32Config.fir@5873.4]
  wire [2:0] _T_892; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@6866.4]
  reg [2:0] _T_898; // @[Arbiter.scala 22:23:freechips.rocketchip.system.DefaultRV32Config.fir@6876.4]
  wire [2:0] _T_899; // @[Arbiter.scala 23:30:freechips.rocketchip.system.DefaultRV32Config.fir@6877.4]
  wire [2:0] _T_900; // @[Arbiter.scala 23:28:freechips.rocketchip.system.DefaultRV32Config.fir@6878.4]
  wire [5:0] _T_901; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@6879.4]
  wire [5:0] _GEN_5; // @[package.scala 226:43:freechips.rocketchip.system.DefaultRV32Config.fir@6881.4]
  wire [5:0] _T_903; // @[package.scala 226:43:freechips.rocketchip.system.DefaultRV32Config.fir@6881.4]
  wire [5:0] _GEN_6; // @[package.scala 226:43:freechips.rocketchip.system.DefaultRV32Config.fir@6883.4]
  wire [5:0] _T_905; // @[package.scala 226:43:freechips.rocketchip.system.DefaultRV32Config.fir@6883.4]
  wire [5:0] _T_908; // @[Arbiter.scala 24:66:freechips.rocketchip.system.DefaultRV32Config.fir@6886.4]
  wire [5:0] _GEN_7; // @[Arbiter.scala 24:58:freechips.rocketchip.system.DefaultRV32Config.fir@6887.4]
  wire [5:0] _T_909; // @[Arbiter.scala 24:58:freechips.rocketchip.system.DefaultRV32Config.fir@6887.4]
  wire [2:0] _T_912; // @[Arbiter.scala 25:39:freechips.rocketchip.system.DefaultRV32Config.fir@6890.4]
  wire [2:0] _T_913; // @[Arbiter.scala 25:18:freechips.rocketchip.system.DefaultRV32Config.fir@6891.4]
  wire  _T_929; // @[Arbiter.scala 88:79:freechips.rocketchip.system.DefaultRV32Config.fir@6913.4]
  reg  _T_984_0; // @[Arbiter.scala 107:26:freechips.rocketchip.system.DefaultRV32Config.fir@6990.4]
  wire  _T_985_0; // @[Arbiter.scala 108:30:freechips.rocketchip.system.DefaultRV32Config.fir@6991.4]
  wire [1:0] _T_20_0_d_bits_sink; // @[Xbar.scala 282:19:freechips.rocketchip.system.DefaultRV32Config.fir@5123.4 BundleMap.scala 248:19:freechips.rocketchip.system.DefaultRV32Config.fir@5172.4 Xbar.scala 317:28:freechips.rocketchip.system.DefaultRV32Config.fir@5180.4]
  wire [49:0] _T_1012; // @[Mux.scala 27:72:freechips.rocketchip.system.DefaultRV32Config.fir@7028.4]
  wire [49:0] _T_1013; // @[Mux.scala 27:72:freechips.rocketchip.system.DefaultRV32Config.fir@7029.4]
  wire  _T_930; // @[Arbiter.scala 88:79:freechips.rocketchip.system.DefaultRV32Config.fir@6914.4]
  reg  _T_984_1; // @[Arbiter.scala 107:26:freechips.rocketchip.system.DefaultRV32Config.fir@6990.4]
  wire  _T_985_1; // @[Arbiter.scala 108:30:freechips.rocketchip.system.DefaultRV32Config.fir@6991.4]
  wire [3:0] _T_20_1_d_bits_size; // @[Xbar.scala 282:19:freechips.rocketchip.system.DefaultRV32Config.fir@5123.4 BundleMap.scala 248:19:freechips.rocketchip.system.DefaultRV32Config.fir@5227.4]
  wire [49:0] _T_1020; // @[Mux.scala 27:72:freechips.rocketchip.system.DefaultRV32Config.fir@7036.4]
  wire [49:0] _T_1021; // @[Mux.scala 27:72:freechips.rocketchip.system.DefaultRV32Config.fir@7037.4]
  wire [49:0] _T_1030; // @[Mux.scala 27:72:freechips.rocketchip.system.DefaultRV32Config.fir@7046.4]
  wire  _T_931; // @[Arbiter.scala 88:79:freechips.rocketchip.system.DefaultRV32Config.fir@6915.4]
  reg  _T_984_2; // @[Arbiter.scala 107:26:freechips.rocketchip.system.DefaultRV32Config.fir@6990.4]
  wire  _T_985_2; // @[Arbiter.scala 108:30:freechips.rocketchip.system.DefaultRV32Config.fir@6991.4]
  wire [49:0] _T_1028; // @[Mux.scala 27:72:freechips.rocketchip.system.DefaultRV32Config.fir@7044.4]
  wire [49:0] _T_1029; // @[Mux.scala 27:72:freechips.rocketchip.system.DefaultRV32Config.fir@7045.4]
  wire [49:0] _T_1031; // @[Mux.scala 27:72:freechips.rocketchip.system.DefaultRV32Config.fir@7047.4]
  wire [4:0] _GEN_8; // @[Xbar.scala 231:55:freechips.rocketchip.system.DefaultRV32Config.fir@5083.4]
  wire [4:0] _T_16; // @[Xbar.scala 231:55:freechips.rocketchip.system.DefaultRV32Config.fir@5083.4]
  wire [4:0] _GEN_9; // @[Xbar.scala 253:55:freechips.rocketchip.system.DefaultRV32Config.fir@5106.4]
  reg [9:0] _T_1054; // @[Arbiter.scala 78:30:freechips.rocketchip.system.DefaultRV32Config.fir@7185.4]
  wire  _T_1055; // @[Arbiter.scala 79:28:freechips.rocketchip.system.DefaultRV32Config.fir@7186.4]
  wire  _T_188; // @[Parameters.scala 55:32:freechips.rocketchip.system.DefaultRV32Config.fir@5470.4]
  wire  _T_385; // @[Xbar.scala 173:40:freechips.rocketchip.system.DefaultRV32Config.fir@5942.4]
  wire  _T_172; // @[Parameters.scala 55:32:freechips.rocketchip.system.DefaultRV32Config.fir@5454.4]
  wire  _T_376; // @[Xbar.scala 173:40:freechips.rocketchip.system.DefaultRV32Config.fir@5913.4]
  wire  _T_156; // @[Parameters.scala 55:32:freechips.rocketchip.system.DefaultRV32Config.fir@5438.4]
  wire  _T_367; // @[Xbar.scala 173:40:freechips.rocketchip.system.DefaultRV32Config.fir@5884.4]
  wire [2:0] _T_1064; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@7195.4]
  reg [2:0] _T_1070; // @[Arbiter.scala 22:23:freechips.rocketchip.system.DefaultRV32Config.fir@7205.4]
  wire [2:0] _T_1071; // @[Arbiter.scala 23:30:freechips.rocketchip.system.DefaultRV32Config.fir@7206.4]
  wire [2:0] _T_1072; // @[Arbiter.scala 23:28:freechips.rocketchip.system.DefaultRV32Config.fir@7207.4]
  wire [5:0] _T_1073; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@7208.4]
  wire [5:0] _GEN_10; // @[package.scala 226:43:freechips.rocketchip.system.DefaultRV32Config.fir@7210.4]
  wire [5:0] _T_1075; // @[package.scala 226:43:freechips.rocketchip.system.DefaultRV32Config.fir@7210.4]
  wire [5:0] _GEN_11; // @[package.scala 226:43:freechips.rocketchip.system.DefaultRV32Config.fir@7212.4]
  wire [5:0] _T_1077; // @[package.scala 226:43:freechips.rocketchip.system.DefaultRV32Config.fir@7212.4]
  wire [5:0] _T_1080; // @[Arbiter.scala 24:66:freechips.rocketchip.system.DefaultRV32Config.fir@7215.4]
  wire [5:0] _GEN_12; // @[Arbiter.scala 24:58:freechips.rocketchip.system.DefaultRV32Config.fir@7216.4]
  wire [5:0] _T_1081; // @[Arbiter.scala 24:58:freechips.rocketchip.system.DefaultRV32Config.fir@7216.4]
  wire [2:0] _T_1084; // @[Arbiter.scala 25:39:freechips.rocketchip.system.DefaultRV32Config.fir@7219.4]
  wire [2:0] _T_1085; // @[Arbiter.scala 25:18:freechips.rocketchip.system.DefaultRV32Config.fir@7220.4]
  wire  _T_1101; // @[Arbiter.scala 88:79:freechips.rocketchip.system.DefaultRV32Config.fir@7242.4]
  reg  _T_1156_0; // @[Arbiter.scala 107:26:freechips.rocketchip.system.DefaultRV32Config.fir@7319.4]
  wire  _T_1157_0; // @[Arbiter.scala 108:30:freechips.rocketchip.system.DefaultRV32Config.fir@7320.4]
  wire [49:0] _T_1185; // @[Mux.scala 27:72:freechips.rocketchip.system.DefaultRV32Config.fir@7358.4]
  wire  _T_1102; // @[Arbiter.scala 88:79:freechips.rocketchip.system.DefaultRV32Config.fir@7243.4]
  reg  _T_1156_1; // @[Arbiter.scala 107:26:freechips.rocketchip.system.DefaultRV32Config.fir@7319.4]
  wire  _T_1157_1; // @[Arbiter.scala 108:30:freechips.rocketchip.system.DefaultRV32Config.fir@7320.4]
  wire [49:0] _T_1193; // @[Mux.scala 27:72:freechips.rocketchip.system.DefaultRV32Config.fir@7366.4]
  wire [49:0] _T_1202; // @[Mux.scala 27:72:freechips.rocketchip.system.DefaultRV32Config.fir@7375.4]
  wire  _T_1103; // @[Arbiter.scala 88:79:freechips.rocketchip.system.DefaultRV32Config.fir@7244.4]
  reg  _T_1156_2; // @[Arbiter.scala 107:26:freechips.rocketchip.system.DefaultRV32Config.fir@7319.4]
  wire  _T_1157_2; // @[Arbiter.scala 108:30:freechips.rocketchip.system.DefaultRV32Config.fir@7320.4]
  wire [49:0] _T_1201; // @[Mux.scala 27:72:freechips.rocketchip.system.DefaultRV32Config.fir@7374.4]
  wire [49:0] _T_1203; // @[Mux.scala 27:72:freechips.rocketchip.system.DefaultRV32Config.fir@7376.4]
  wire [32:0] _T_26; // @[Parameters.scala 137:49:freechips.rocketchip.system.DefaultRV32Config.fir@5308.4]
  wire [32:0] _T_28; // @[Parameters.scala 137:52:freechips.rocketchip.system.DefaultRV32Config.fir@5310.4]
  wire  _T_29; // @[Parameters.scala 137:67:freechips.rocketchip.system.DefaultRV32Config.fir@5311.4]
  wire [31:0] _T_31; // @[Parameters.scala 137:31:freechips.rocketchip.system.DefaultRV32Config.fir@5313.4]
  wire [32:0] _T_32; // @[Parameters.scala 137:49:freechips.rocketchip.system.DefaultRV32Config.fir@5314.4]
  wire [32:0] _T_34; // @[Parameters.scala 137:52:freechips.rocketchip.system.DefaultRV32Config.fir@5316.4]
  wire  _T_35; // @[Parameters.scala 137:67:freechips.rocketchip.system.DefaultRV32Config.fir@5317.4]
  wire [31:0] _T_37; // @[Parameters.scala 137:31:freechips.rocketchip.system.DefaultRV32Config.fir@5319.4]
  wire [32:0] _T_38; // @[Parameters.scala 137:49:freechips.rocketchip.system.DefaultRV32Config.fir@5320.4]
  wire [32:0] _T_40; // @[Parameters.scala 137:52:freechips.rocketchip.system.DefaultRV32Config.fir@5322.4]
  wire  _T_41; // @[Parameters.scala 137:67:freechips.rocketchip.system.DefaultRV32Config.fir@5323.4]
  wire [32:0] _T_44; // @[Parameters.scala 137:49:freechips.rocketchip.system.DefaultRV32Config.fir@5326.4]
  wire [32:0] _T_46; // @[Parameters.scala 137:52:freechips.rocketchip.system.DefaultRV32Config.fir@5328.4]
  wire  _T_47; // @[Parameters.scala 137:67:freechips.rocketchip.system.DefaultRV32Config.fir@5329.4]
  wire [31:0] _T_49; // @[Parameters.scala 137:31:freechips.rocketchip.system.DefaultRV32Config.fir@5331.4]
  wire [32:0] _T_50; // @[Parameters.scala 137:49:freechips.rocketchip.system.DefaultRV32Config.fir@5332.4]
  wire [32:0] _T_52; // @[Parameters.scala 137:52:freechips.rocketchip.system.DefaultRV32Config.fir@5334.4]
  wire  _T_53; // @[Parameters.scala 137:67:freechips.rocketchip.system.DefaultRV32Config.fir@5335.4]
  wire [31:0] _T_55; // @[Parameters.scala 137:31:freechips.rocketchip.system.DefaultRV32Config.fir@5337.4]
  wire [32:0] _T_56; // @[Parameters.scala 137:49:freechips.rocketchip.system.DefaultRV32Config.fir@5338.4]
  wire [32:0] _T_58; // @[Parameters.scala 137:52:freechips.rocketchip.system.DefaultRV32Config.fir@5340.4]
  wire  _T_59; // @[Parameters.scala 137:67:freechips.rocketchip.system.DefaultRV32Config.fir@5341.4]
  wire [26:0] _T_210; // @[package.scala 207:77:freechips.rocketchip.system.DefaultRV32Config.fir@5492.4]
  wire [11:0] _T_212; // @[package.scala 207:46:freechips.rocketchip.system.DefaultRV32Config.fir@5494.4]
  wire  _T_215; // @[Edges.scala 93:28:freechips.rocketchip.system.DefaultRV32Config.fir@5497.4]
  wire [9:0] _T_216; // @[Edges.scala 222:14:freechips.rocketchip.system.DefaultRV32Config.fir@5498.4]
  wire [26:0] _T_218; // @[package.scala 207:77:freechips.rocketchip.system.DefaultRV32Config.fir@5500.4]
  wire [11:0] _T_220; // @[package.scala 207:46:freechips.rocketchip.system.DefaultRV32Config.fir@5502.4]
  wire  _T_223; // @[Edges.scala 93:28:freechips.rocketchip.system.DefaultRV32Config.fir@5505.4]
  wire [9:0] _T_224; // @[Edges.scala 222:14:freechips.rocketchip.system.DefaultRV32Config.fir@5506.4]
  wire [26:0] _T_264; // @[package.scala 207:77:freechips.rocketchip.system.DefaultRV32Config.fir@5546.4]
  wire [11:0] _T_266; // @[package.scala 207:46:freechips.rocketchip.system.DefaultRV32Config.fir@5548.4]
  wire [9:0] _T_269; // @[Edges.scala 222:14:freechips.rocketchip.system.DefaultRV32Config.fir@5551.4]
  wire [20:0] _T_271; // @[package.scala 207:77:freechips.rocketchip.system.DefaultRV32Config.fir@5553.4]
  wire [5:0] _T_273; // @[package.scala 207:46:freechips.rocketchip.system.DefaultRV32Config.fir@5555.4]
  wire [3:0] _T_276; // @[Edges.scala 222:14:freechips.rocketchip.system.DefaultRV32Config.fir@5558.4]
  wire [22:0] _T_278; // @[package.scala 207:77:freechips.rocketchip.system.DefaultRV32Config.fir@5560.4]
  wire [7:0] _T_280; // @[package.scala 207:46:freechips.rocketchip.system.DefaultRV32Config.fir@5562.4]
  wire [5:0] _T_283; // @[Edges.scala 222:14:freechips.rocketchip.system.DefaultRV32Config.fir@5565.4]
  wire  _T_286; // @[Xbar.scala 422:50:freechips.rocketchip.system.DefaultRV32Config.fir@5584.4]
  wire  _T_288; // @[Xbar.scala 422:50:freechips.rocketchip.system.DefaultRV32Config.fir@5603.4]
  wire  _T_290; // @[Xbar.scala 422:50:freechips.rocketchip.system.DefaultRV32Config.fir@5622.4]
  reg [9:0] _T_416; // @[Arbiter.scala 78:30:freechips.rocketchip.system.DefaultRV32Config.fir@5992.4]
  wire  _T_417; // @[Arbiter.scala 79:28:freechips.rocketchip.system.DefaultRV32Config.fir@5993.4]
  wire  _T_299; // @[Xbar.scala 422:50:freechips.rocketchip.system.DefaultRV32Config.fir@5650.4]
  wire [1:0] _T_423; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@5999.4]
  reg [1:0] _T_429; // @[Arbiter.scala 22:23:freechips.rocketchip.system.DefaultRV32Config.fir@6009.4]
  wire [1:0] _T_430; // @[Arbiter.scala 23:30:freechips.rocketchip.system.DefaultRV32Config.fir@6010.4]
  wire [1:0] _T_431; // @[Arbiter.scala 23:28:freechips.rocketchip.system.DefaultRV32Config.fir@6011.4]
  wire [3:0] _T_432; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@6012.4]
  wire [3:0] _GEN_13; // @[package.scala 226:43:freechips.rocketchip.system.DefaultRV32Config.fir@6014.4]
  wire [3:0] _T_434; // @[package.scala 226:43:freechips.rocketchip.system.DefaultRV32Config.fir@6014.4]
  wire [3:0] _T_437; // @[Arbiter.scala 24:66:freechips.rocketchip.system.DefaultRV32Config.fir@6017.4]
  wire [3:0] _GEN_14; // @[Arbiter.scala 24:58:freechips.rocketchip.system.DefaultRV32Config.fir@6018.4]
  wire [3:0] _T_438; // @[Arbiter.scala 24:58:freechips.rocketchip.system.DefaultRV32Config.fir@6018.4]
  wire [1:0] _T_441; // @[Arbiter.scala 25:39:freechips.rocketchip.system.DefaultRV32Config.fir@6021.4]
  wire [1:0] _T_442; // @[Arbiter.scala 25:18:freechips.rocketchip.system.DefaultRV32Config.fir@6022.4]
  reg  _T_496_0; // @[Arbiter.scala 107:26:freechips.rocketchip.system.DefaultRV32Config.fir@6100.4]
  wire  _T_499_0; // @[Arbiter.scala 112:24:freechips.rocketchip.system.DefaultRV32Config.fir@6105.4]
  wire  _T_500; // @[Arbiter.scala 114:31:freechips.rocketchip.system.DefaultRV32Config.fir@6106.4]
  wire  _T_291; // @[Mux.scala 27:72:freechips.rocketchip.system.DefaultRV32Config.fir@5624.4]
  reg [9:0] _T_568; // @[Arbiter.scala 78:30:freechips.rocketchip.system.DefaultRV32Config.fir@6251.4]
  wire  _T_569; // @[Arbiter.scala 79:28:freechips.rocketchip.system.DefaultRV32Config.fir@6252.4]
  wire  _T_301; // @[Xbar.scala 422:50:freechips.rocketchip.system.DefaultRV32Config.fir@5669.4]
  wire [1:0] _T_575; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@6258.4]
  reg [1:0] _T_581; // @[Arbiter.scala 22:23:freechips.rocketchip.system.DefaultRV32Config.fir@6268.4]
  wire [1:0] _T_582; // @[Arbiter.scala 23:30:freechips.rocketchip.system.DefaultRV32Config.fir@6269.4]
  wire [1:0] _T_583; // @[Arbiter.scala 23:28:freechips.rocketchip.system.DefaultRV32Config.fir@6270.4]
  wire [3:0] _T_584; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@6271.4]
  wire [3:0] _GEN_15; // @[package.scala 226:43:freechips.rocketchip.system.DefaultRV32Config.fir@6273.4]
  wire [3:0] _T_586; // @[package.scala 226:43:freechips.rocketchip.system.DefaultRV32Config.fir@6273.4]
  wire [3:0] _T_589; // @[Arbiter.scala 24:66:freechips.rocketchip.system.DefaultRV32Config.fir@6276.4]
  wire [3:0] _GEN_16; // @[Arbiter.scala 24:58:freechips.rocketchip.system.DefaultRV32Config.fir@6277.4]
  wire [3:0] _T_590; // @[Arbiter.scala 24:58:freechips.rocketchip.system.DefaultRV32Config.fir@6277.4]
  wire [1:0] _T_593; // @[Arbiter.scala 25:39:freechips.rocketchip.system.DefaultRV32Config.fir@6280.4]
  wire [1:0] _T_594; // @[Arbiter.scala 25:18:freechips.rocketchip.system.DefaultRV32Config.fir@6281.4]
  reg  _T_648_0; // @[Arbiter.scala 107:26:freechips.rocketchip.system.DefaultRV32Config.fir@6359.4]
  wire  _T_651_0; // @[Arbiter.scala 112:24:freechips.rocketchip.system.DefaultRV32Config.fir@6364.4]
  wire  _T_652; // @[Arbiter.scala 114:31:freechips.rocketchip.system.DefaultRV32Config.fir@6365.4]
  wire  _T_292; // @[Mux.scala 27:72:freechips.rocketchip.system.DefaultRV32Config.fir@5625.4]
  reg [9:0] _T_722; // @[Arbiter.scala 78:30:freechips.rocketchip.system.DefaultRV32Config.fir@6526.4]
  wire  _T_723; // @[Arbiter.scala 79:28:freechips.rocketchip.system.DefaultRV32Config.fir@6527.4]
  wire  _T_303; // @[Xbar.scala 422:50:freechips.rocketchip.system.DefaultRV32Config.fir@5688.4]
  wire [1:0] _T_729; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@6533.4]
  reg [1:0] _T_735; // @[Arbiter.scala 22:23:freechips.rocketchip.system.DefaultRV32Config.fir@6543.4]
  wire [1:0] _T_736; // @[Arbiter.scala 23:30:freechips.rocketchip.system.DefaultRV32Config.fir@6544.4]
  wire [1:0] _T_737; // @[Arbiter.scala 23:28:freechips.rocketchip.system.DefaultRV32Config.fir@6545.4]
  wire [3:0] _T_738; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@6546.4]
  wire [3:0] _GEN_17; // @[package.scala 226:43:freechips.rocketchip.system.DefaultRV32Config.fir@6548.4]
  wire [3:0] _T_740; // @[package.scala 226:43:freechips.rocketchip.system.DefaultRV32Config.fir@6548.4]
  wire [3:0] _T_743; // @[Arbiter.scala 24:66:freechips.rocketchip.system.DefaultRV32Config.fir@6551.4]
  wire [3:0] _GEN_18; // @[Arbiter.scala 24:58:freechips.rocketchip.system.DefaultRV32Config.fir@6552.4]
  wire [3:0] _T_744; // @[Arbiter.scala 24:58:freechips.rocketchip.system.DefaultRV32Config.fir@6552.4]
  wire [1:0] _T_747; // @[Arbiter.scala 25:39:freechips.rocketchip.system.DefaultRV32Config.fir@6555.4]
  wire [1:0] _T_748; // @[Arbiter.scala 25:18:freechips.rocketchip.system.DefaultRV32Config.fir@6556.4]
  reg  _T_802_0; // @[Arbiter.scala 107:26:freechips.rocketchip.system.DefaultRV32Config.fir@6634.4]
  wire  _T_805_0; // @[Arbiter.scala 112:24:freechips.rocketchip.system.DefaultRV32Config.fir@6639.4]
  wire  _T_806; // @[Arbiter.scala 114:31:freechips.rocketchip.system.DefaultRV32Config.fir@6640.4]
  wire  _T_293; // @[Mux.scala 27:72:freechips.rocketchip.system.DefaultRV32Config.fir@5626.4]
  wire  _T_294; // @[Mux.scala 27:72:freechips.rocketchip.system.DefaultRV32Config.fir@5627.4]
  reg  _T_496_1; // @[Arbiter.scala 107:26:freechips.rocketchip.system.DefaultRV32Config.fir@6100.4]
  wire  _T_499_1; // @[Arbiter.scala 112:24:freechips.rocketchip.system.DefaultRV32Config.fir@6105.4]
  wire  _T_501; // @[Arbiter.scala 114:31:freechips.rocketchip.system.DefaultRV32Config.fir@6108.4]
  wire  _T_304; // @[Mux.scala 27:72:freechips.rocketchip.system.DefaultRV32Config.fir@5690.4]
  reg  _T_648_1; // @[Arbiter.scala 107:26:freechips.rocketchip.system.DefaultRV32Config.fir@6359.4]
  wire  _T_651_1; // @[Arbiter.scala 112:24:freechips.rocketchip.system.DefaultRV32Config.fir@6364.4]
  wire  _T_653; // @[Arbiter.scala 114:31:freechips.rocketchip.system.DefaultRV32Config.fir@6367.4]
  wire  _T_305; // @[Mux.scala 27:72:freechips.rocketchip.system.DefaultRV32Config.fir@5691.4]
  reg  _T_802_1; // @[Arbiter.scala 107:26:freechips.rocketchip.system.DefaultRV32Config.fir@6634.4]
  wire  _T_805_1; // @[Arbiter.scala 112:24:freechips.rocketchip.system.DefaultRV32Config.fir@6639.4]
  wire  _T_807; // @[Arbiter.scala 114:31:freechips.rocketchip.system.DefaultRV32Config.fir@6642.4]
  wire  _T_306; // @[Mux.scala 27:72:freechips.rocketchip.system.DefaultRV32Config.fir@5692.4]
  wire  _T_307; // @[Mux.scala 27:72:freechips.rocketchip.system.DefaultRV32Config.fir@5693.4]
  wire  _T_987_0; // @[Arbiter.scala 112:24:freechips.rocketchip.system.DefaultRV32Config.fir@6996.4]
  wire  _T_988; // @[Arbiter.scala 114:31:freechips.rocketchip.system.DefaultRV32Config.fir@6997.4]
  wire  _T_368; // @[Mux.scala 27:72:freechips.rocketchip.system.DefaultRV32Config.fir@5886.4]
  wire  _T_1159_0; // @[Arbiter.scala 112:24:freechips.rocketchip.system.DefaultRV32Config.fir@7325.4]
  wire  _T_1160; // @[Arbiter.scala 114:31:freechips.rocketchip.system.DefaultRV32Config.fir@7326.4]
  wire  _T_369; // @[Mux.scala 27:72:freechips.rocketchip.system.DefaultRV32Config.fir@5887.4]
  wire  _T_987_1; // @[Arbiter.scala 112:24:freechips.rocketchip.system.DefaultRV32Config.fir@6996.4]
  wire  _T_989; // @[Arbiter.scala 114:31:freechips.rocketchip.system.DefaultRV32Config.fir@6999.4]
  wire  _T_377; // @[Mux.scala 27:72:freechips.rocketchip.system.DefaultRV32Config.fir@5915.4]
  wire  _T_1159_1; // @[Arbiter.scala 112:24:freechips.rocketchip.system.DefaultRV32Config.fir@7325.4]
  wire  _T_1161; // @[Arbiter.scala 114:31:freechips.rocketchip.system.DefaultRV32Config.fir@7328.4]
  wire  _T_378; // @[Mux.scala 27:72:freechips.rocketchip.system.DefaultRV32Config.fir@5916.4]
  wire  _T_987_2; // @[Arbiter.scala 112:24:freechips.rocketchip.system.DefaultRV32Config.fir@6996.4]
  wire  _T_990; // @[Arbiter.scala 114:31:freechips.rocketchip.system.DefaultRV32Config.fir@7001.4]
  wire  _T_386; // @[Mux.scala 27:72:freechips.rocketchip.system.DefaultRV32Config.fir@5944.4]
  wire  _T_1159_2; // @[Arbiter.scala 112:24:freechips.rocketchip.system.DefaultRV32Config.fir@7325.4]
  wire  _T_1162; // @[Arbiter.scala 114:31:freechips.rocketchip.system.DefaultRV32Config.fir@7330.4]
  wire  _T_387; // @[Mux.scala 27:72:freechips.rocketchip.system.DefaultRV32Config.fir@5945.4]
  wire  _T_418; // @[Arbiter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@5994.4]
  wire  _T_443; // @[Arbiter.scala 26:27:freechips.rocketchip.system.DefaultRV32Config.fir@6023.4]
  wire  _T_444; // @[Arbiter.scala 26:18:freechips.rocketchip.system.DefaultRV32Config.fir@6024.4]
  wire [1:0] _T_445; // @[Arbiter.scala 27:29:freechips.rocketchip.system.DefaultRV32Config.fir@6026.6]
  wire [2:0] _T_446; // @[package.scala 217:48:freechips.rocketchip.system.DefaultRV32Config.fir@6027.6]
  wire [1:0] _T_448; // @[package.scala 217:43:freechips.rocketchip.system.DefaultRV32Config.fir@6029.6]
  wire  _T_454; // @[Arbiter.scala 88:79:freechips.rocketchip.system.DefaultRV32Config.fir@6039.4]
  wire  _T_455; // @[Arbiter.scala 88:79:freechips.rocketchip.system.DefaultRV32Config.fir@6040.4]
  wire  _T_461; // @[Arbiter.scala 95:53:freechips.rocketchip.system.DefaultRV32Config.fir@6050.4]
  wire  _T_463; // @[Arbiter.scala 96:67:freechips.rocketchip.system.DefaultRV32Config.fir@6052.4]
  wire  _T_466; // @[Arbiter.scala 96:67:freechips.rocketchip.system.DefaultRV32Config.fir@6055.4]
  wire  _T_467; // @[Arbiter.scala 96:64:freechips.rocketchip.system.DefaultRV32Config.fir@6056.4]
  wire  _T_470; // @[Arbiter.scala 96:13:freechips.rocketchip.system.DefaultRV32Config.fir@6059.4]
  wire  _T_471; // @[Arbiter.scala 96:13:freechips.rocketchip.system.DefaultRV32Config.fir@6060.4]
  wire  _T_472; // @[Arbiter.scala 98:36:freechips.rocketchip.system.DefaultRV32Config.fir@6065.4]
  wire  _T_473; // @[Arbiter.scala 98:15:freechips.rocketchip.system.DefaultRV32Config.fir@6066.4]
  wire  _T_475; // @[Arbiter.scala 98:41:freechips.rocketchip.system.DefaultRV32Config.fir@6068.4]
  wire  _T_477; // @[Arbiter.scala 98:14:freechips.rocketchip.system.DefaultRV32Config.fir@6070.4]
  wire  _T_478; // @[Arbiter.scala 98:14:freechips.rocketchip.system.DefaultRV32Config.fir@6071.4]
  wire  _T_482; // @[Arbiter.scala 99:41:freechips.rocketchip.system.DefaultRV32Config.fir@6079.4]
  wire  _T_484; // @[Arbiter.scala 99:14:freechips.rocketchip.system.DefaultRV32Config.fir@6081.4]
  wire  _T_485; // @[Arbiter.scala 99:14:freechips.rocketchip.system.DefaultRV32Config.fir@6082.4]
  wire [9:0] _T_486; // @[Arbiter.scala 102:73:freechips.rocketchip.system.DefaultRV32Config.fir@6087.4]
  wire [9:0] _T_487; // @[Arbiter.scala 102:73:freechips.rocketchip.system.DefaultRV32Config.fir@6088.4]
  wire [9:0] _T_488; // @[Arbiter.scala 103:44:freechips.rocketchip.system.DefaultRV32Config.fir@6089.4]
  wire  _T_497_0; // @[Arbiter.scala 108:30:freechips.rocketchip.system.DefaultRV32Config.fir@6101.4]
  wire  _T_497_1; // @[Arbiter.scala 108:30:freechips.rocketchip.system.DefaultRV32Config.fir@6101.4]
  wire  _T_503; // @[Mux.scala 27:72:freechips.rocketchip.system.DefaultRV32Config.fir@6111.4]
  wire  _T_504; // @[Mux.scala 27:72:freechips.rocketchip.system.DefaultRV32Config.fir@6112.4]
  wire  _T_505; // @[Mux.scala 27:72:freechips.rocketchip.system.DefaultRV32Config.fir@6113.4]
  wire  _T_507; // @[Arbiter.scala 116:29:freechips.rocketchip.system.DefaultRV32Config.fir@6116.4]
  wire  _T_491; // @[ReadyValidCancel.scala 52:33:freechips.rocketchip.system.DefaultRV32Config.fir@6092.4]
  wire [9:0] _GEN_19; // @[Arbiter.scala 104:52:freechips.rocketchip.system.DefaultRV32Config.fir@6093.4]
  wire [9:0] _T_493; // @[Arbiter.scala 104:52:freechips.rocketchip.system.DefaultRV32Config.fir@6094.4]
  wire [40:0] _T_517; // @[Mux.scala 27:72:freechips.rocketchip.system.DefaultRV32Config.fir@6129.4]
  wire [4:0] _T_13_0_a_bits_source; // @[Xbar.scala 225:18:freechips.rocketchip.system.DefaultRV32Config.fir@4994.4 BundleMap.scala 248:19:freechips.rocketchip.system.DefaultRV32Config.fir@5006.4 Xbar.scala 231:29:freechips.rocketchip.system.DefaultRV32Config.fir@5014.4]
  wire [90:0] _T_525; // @[Mux.scala 27:72:freechips.rocketchip.system.DefaultRV32Config.fir@6137.4]
  wire [90:0] _T_526; // @[Mux.scala 27:72:freechips.rocketchip.system.DefaultRV32Config.fir@6138.4]
  wire [40:0] _T_532; // @[Mux.scala 27:72:freechips.rocketchip.system.DefaultRV32Config.fir@6144.4]
  wire [90:0] _T_540; // @[Mux.scala 27:72:freechips.rocketchip.system.DefaultRV32Config.fir@6152.4]
  wire [90:0] _T_541; // @[Mux.scala 27:72:freechips.rocketchip.system.DefaultRV32Config.fir@6153.4]
  wire [90:0] _T_542; // @[Mux.scala 27:72:freechips.rocketchip.system.DefaultRV32Config.fir@6154.4]
  wire  _T_570; // @[Arbiter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@6253.4]
  wire  _T_595; // @[Arbiter.scala 26:27:freechips.rocketchip.system.DefaultRV32Config.fir@6282.4]
  wire  _T_596; // @[Arbiter.scala 26:18:freechips.rocketchip.system.DefaultRV32Config.fir@6283.4]
  wire [1:0] _T_597; // @[Arbiter.scala 27:29:freechips.rocketchip.system.DefaultRV32Config.fir@6285.6]
  wire [2:0] _T_598; // @[package.scala 217:48:freechips.rocketchip.system.DefaultRV32Config.fir@6286.6]
  wire [1:0] _T_600; // @[package.scala 217:43:freechips.rocketchip.system.DefaultRV32Config.fir@6288.6]
  wire  _T_606; // @[Arbiter.scala 88:79:freechips.rocketchip.system.DefaultRV32Config.fir@6298.4]
  wire  _T_607; // @[Arbiter.scala 88:79:freechips.rocketchip.system.DefaultRV32Config.fir@6299.4]
  wire  _T_613; // @[Arbiter.scala 95:53:freechips.rocketchip.system.DefaultRV32Config.fir@6309.4]
  wire  _T_615; // @[Arbiter.scala 96:67:freechips.rocketchip.system.DefaultRV32Config.fir@6311.4]
  wire  _T_618; // @[Arbiter.scala 96:67:freechips.rocketchip.system.DefaultRV32Config.fir@6314.4]
  wire  _T_619; // @[Arbiter.scala 96:64:freechips.rocketchip.system.DefaultRV32Config.fir@6315.4]
  wire  _T_622; // @[Arbiter.scala 96:13:freechips.rocketchip.system.DefaultRV32Config.fir@6318.4]
  wire  _T_623; // @[Arbiter.scala 96:13:freechips.rocketchip.system.DefaultRV32Config.fir@6319.4]
  wire  _T_624; // @[Arbiter.scala 98:36:freechips.rocketchip.system.DefaultRV32Config.fir@6324.4]
  wire  _T_625; // @[Arbiter.scala 98:15:freechips.rocketchip.system.DefaultRV32Config.fir@6325.4]
  wire  _T_627; // @[Arbiter.scala 98:41:freechips.rocketchip.system.DefaultRV32Config.fir@6327.4]
  wire  _T_629; // @[Arbiter.scala 98:14:freechips.rocketchip.system.DefaultRV32Config.fir@6329.4]
  wire  _T_630; // @[Arbiter.scala 98:14:freechips.rocketchip.system.DefaultRV32Config.fir@6330.4]
  wire  _T_634; // @[Arbiter.scala 99:41:freechips.rocketchip.system.DefaultRV32Config.fir@6338.4]
  wire  _T_636; // @[Arbiter.scala 99:14:freechips.rocketchip.system.DefaultRV32Config.fir@6340.4]
  wire  _T_637; // @[Arbiter.scala 99:14:freechips.rocketchip.system.DefaultRV32Config.fir@6341.4]
  wire [9:0] _T_638; // @[Arbiter.scala 102:73:freechips.rocketchip.system.DefaultRV32Config.fir@6346.4]
  wire [9:0] _T_639; // @[Arbiter.scala 102:73:freechips.rocketchip.system.DefaultRV32Config.fir@6347.4]
  wire [9:0] _T_640; // @[Arbiter.scala 103:44:freechips.rocketchip.system.DefaultRV32Config.fir@6348.4]
  wire  _T_649_0; // @[Arbiter.scala 108:30:freechips.rocketchip.system.DefaultRV32Config.fir@6360.4]
  wire  _T_649_1; // @[Arbiter.scala 108:30:freechips.rocketchip.system.DefaultRV32Config.fir@6360.4]
  wire  _T_655; // @[Mux.scala 27:72:freechips.rocketchip.system.DefaultRV32Config.fir@6370.4]
  wire  _T_656; // @[Mux.scala 27:72:freechips.rocketchip.system.DefaultRV32Config.fir@6371.4]
  wire  _T_657; // @[Mux.scala 27:72:freechips.rocketchip.system.DefaultRV32Config.fir@6372.4]
  wire  _T_659; // @[Arbiter.scala 116:29:freechips.rocketchip.system.DefaultRV32Config.fir@6375.4]
  wire  _T_643; // @[ReadyValidCancel.scala 52:33:freechips.rocketchip.system.DefaultRV32Config.fir@6351.4]
  wire [9:0] _GEN_20; // @[Arbiter.scala 104:52:freechips.rocketchip.system.DefaultRV32Config.fir@6352.4]
  wire [9:0] _T_645; // @[Arbiter.scala 104:52:freechips.rocketchip.system.DefaultRV32Config.fir@6353.4]
  wire [90:0] _T_678; // @[Mux.scala 27:72:freechips.rocketchip.system.DefaultRV32Config.fir@6397.4]
  wire [90:0] _T_693; // @[Mux.scala 27:72:freechips.rocketchip.system.DefaultRV32Config.fir@6412.4]
  wire [90:0] _T_694; // @[Mux.scala 27:72:freechips.rocketchip.system.DefaultRV32Config.fir@6413.4]
  wire  _T_724; // @[Arbiter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@6528.4]
  wire  _T_749; // @[Arbiter.scala 26:27:freechips.rocketchip.system.DefaultRV32Config.fir@6557.4]
  wire  _T_750; // @[Arbiter.scala 26:18:freechips.rocketchip.system.DefaultRV32Config.fir@6558.4]
  wire [1:0] _T_751; // @[Arbiter.scala 27:29:freechips.rocketchip.system.DefaultRV32Config.fir@6560.6]
  wire [2:0] _T_752; // @[package.scala 217:48:freechips.rocketchip.system.DefaultRV32Config.fir@6561.6]
  wire [1:0] _T_754; // @[package.scala 217:43:freechips.rocketchip.system.DefaultRV32Config.fir@6563.6]
  wire  _T_760; // @[Arbiter.scala 88:79:freechips.rocketchip.system.DefaultRV32Config.fir@6573.4]
  wire  _T_761; // @[Arbiter.scala 88:79:freechips.rocketchip.system.DefaultRV32Config.fir@6574.4]
  wire  _T_767; // @[Arbiter.scala 95:53:freechips.rocketchip.system.DefaultRV32Config.fir@6584.4]
  wire  _T_769; // @[Arbiter.scala 96:67:freechips.rocketchip.system.DefaultRV32Config.fir@6586.4]
  wire  _T_772; // @[Arbiter.scala 96:67:freechips.rocketchip.system.DefaultRV32Config.fir@6589.4]
  wire  _T_773; // @[Arbiter.scala 96:64:freechips.rocketchip.system.DefaultRV32Config.fir@6590.4]
  wire  _T_776; // @[Arbiter.scala 96:13:freechips.rocketchip.system.DefaultRV32Config.fir@6593.4]
  wire  _T_777; // @[Arbiter.scala 96:13:freechips.rocketchip.system.DefaultRV32Config.fir@6594.4]
  wire  _T_778; // @[Arbiter.scala 98:36:freechips.rocketchip.system.DefaultRV32Config.fir@6599.4]
  wire  _T_779; // @[Arbiter.scala 98:15:freechips.rocketchip.system.DefaultRV32Config.fir@6600.4]
  wire  _T_781; // @[Arbiter.scala 98:41:freechips.rocketchip.system.DefaultRV32Config.fir@6602.4]
  wire  _T_783; // @[Arbiter.scala 98:14:freechips.rocketchip.system.DefaultRV32Config.fir@6604.4]
  wire  _T_784; // @[Arbiter.scala 98:14:freechips.rocketchip.system.DefaultRV32Config.fir@6605.4]
  wire  _T_788; // @[Arbiter.scala 99:41:freechips.rocketchip.system.DefaultRV32Config.fir@6613.4]
  wire  _T_790; // @[Arbiter.scala 99:14:freechips.rocketchip.system.DefaultRV32Config.fir@6615.4]
  wire  _T_791; // @[Arbiter.scala 99:14:freechips.rocketchip.system.DefaultRV32Config.fir@6616.4]
  wire [9:0] _T_792; // @[Arbiter.scala 102:73:freechips.rocketchip.system.DefaultRV32Config.fir@6621.4]
  wire [9:0] _T_793; // @[Arbiter.scala 102:73:freechips.rocketchip.system.DefaultRV32Config.fir@6622.4]
  wire [9:0] _T_794; // @[Arbiter.scala 103:44:freechips.rocketchip.system.DefaultRV32Config.fir@6623.4]
  wire  _T_803_0; // @[Arbiter.scala 108:30:freechips.rocketchip.system.DefaultRV32Config.fir@6635.4]
  wire  _T_803_1; // @[Arbiter.scala 108:30:freechips.rocketchip.system.DefaultRV32Config.fir@6635.4]
  wire  _T_809; // @[Mux.scala 27:72:freechips.rocketchip.system.DefaultRV32Config.fir@6645.4]
  wire  _T_810; // @[Mux.scala 27:72:freechips.rocketchip.system.DefaultRV32Config.fir@6646.4]
  wire  _T_811; // @[Mux.scala 27:72:freechips.rocketchip.system.DefaultRV32Config.fir@6647.4]
  wire  _T_813; // @[Arbiter.scala 116:29:freechips.rocketchip.system.DefaultRV32Config.fir@6650.4]
  wire  _T_797; // @[ReadyValidCancel.scala 52:33:freechips.rocketchip.system.DefaultRV32Config.fir@6626.4]
  wire [9:0] _GEN_21; // @[Arbiter.scala 104:52:freechips.rocketchip.system.DefaultRV32Config.fir@6627.4]
  wire [9:0] _T_799; // @[Arbiter.scala 104:52:freechips.rocketchip.system.DefaultRV32Config.fir@6628.4]
  wire [90:0] _T_832; // @[Mux.scala 27:72:freechips.rocketchip.system.DefaultRV32Config.fir@6672.4]
  wire [90:0] _T_847; // @[Mux.scala 27:72:freechips.rocketchip.system.DefaultRV32Config.fir@6687.4]
  wire [90:0] _T_848; // @[Mux.scala 27:72:freechips.rocketchip.system.DefaultRV32Config.fir@6688.4]
  wire  _T_884; // @[Arbiter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@6858.4]
  wire  _T_914; // @[Arbiter.scala 26:27:freechips.rocketchip.system.DefaultRV32Config.fir@6892.4]
  wire  _T_915; // @[Arbiter.scala 26:18:freechips.rocketchip.system.DefaultRV32Config.fir@6893.4]
  wire [2:0] _T_916; // @[Arbiter.scala 27:29:freechips.rocketchip.system.DefaultRV32Config.fir@6895.6]
  wire [3:0] _T_917; // @[package.scala 217:48:freechips.rocketchip.system.DefaultRV32Config.fir@6896.6]
  wire [2:0] _T_919; // @[package.scala 217:43:freechips.rocketchip.system.DefaultRV32Config.fir@6898.6]
  wire [4:0] _T_920; // @[package.scala 217:48:freechips.rocketchip.system.DefaultRV32Config.fir@6899.6]
  wire [2:0] _T_922; // @[package.scala 217:43:freechips.rocketchip.system.DefaultRV32Config.fir@6901.6]
  wire  _T_938; // @[Arbiter.scala 95:53:freechips.rocketchip.system.DefaultRV32Config.fir@6928.4]
  wire  _T_939; // @[Arbiter.scala 95:53:freechips.rocketchip.system.DefaultRV32Config.fir@6929.4]
  wire  _T_941; // @[Arbiter.scala 96:67:freechips.rocketchip.system.DefaultRV32Config.fir@6931.4]
  wire  _T_944; // @[Arbiter.scala 96:67:freechips.rocketchip.system.DefaultRV32Config.fir@6934.4]
  wire  _T_945; // @[Arbiter.scala 96:64:freechips.rocketchip.system.DefaultRV32Config.fir@6935.4]
  wire  _T_946; // @[Arbiter.scala 96:61:freechips.rocketchip.system.DefaultRV32Config.fir@6936.4]
  wire  _T_947; // @[Arbiter.scala 96:67:freechips.rocketchip.system.DefaultRV32Config.fir@6937.4]
  wire  _T_948; // @[Arbiter.scala 96:64:freechips.rocketchip.system.DefaultRV32Config.fir@6938.4]
  wire  _T_950; // @[Arbiter.scala 96:82:freechips.rocketchip.system.DefaultRV32Config.fir@6940.4]
  wire  _T_952; // @[Arbiter.scala 96:13:freechips.rocketchip.system.DefaultRV32Config.fir@6942.4]
  wire  _T_953; // @[Arbiter.scala 96:13:freechips.rocketchip.system.DefaultRV32Config.fir@6943.4]
  wire  _T_954; // @[Arbiter.scala 98:36:freechips.rocketchip.system.DefaultRV32Config.fir@6948.4]
  wire  _T_955; // @[Arbiter.scala 98:36:freechips.rocketchip.system.DefaultRV32Config.fir@6949.4]
  wire  _T_956; // @[Arbiter.scala 98:15:freechips.rocketchip.system.DefaultRV32Config.fir@6950.4]
  wire  _T_959; // @[Arbiter.scala 98:41:freechips.rocketchip.system.DefaultRV32Config.fir@6953.4]
  wire  _T_961; // @[Arbiter.scala 98:14:freechips.rocketchip.system.DefaultRV32Config.fir@6955.4]
  wire  _T_962; // @[Arbiter.scala 98:14:freechips.rocketchip.system.DefaultRV32Config.fir@6956.4]
  wire  _T_968; // @[Arbiter.scala 99:41:freechips.rocketchip.system.DefaultRV32Config.fir@6966.4]
  wire  _T_970; // @[Arbiter.scala 99:14:freechips.rocketchip.system.DefaultRV32Config.fir@6968.4]
  wire  _T_971; // @[Arbiter.scala 99:14:freechips.rocketchip.system.DefaultRV32Config.fir@6969.4]
  wire [9:0] _T_972; // @[Arbiter.scala 102:73:freechips.rocketchip.system.DefaultRV32Config.fir@6974.4]
  wire [3:0] _T_973; // @[Arbiter.scala 102:73:freechips.rocketchip.system.DefaultRV32Config.fir@6975.4]
  wire [5:0] _T_974; // @[Arbiter.scala 102:73:freechips.rocketchip.system.DefaultRV32Config.fir@6976.4]
  wire [9:0] _GEN_22; // @[Arbiter.scala 103:44:freechips.rocketchip.system.DefaultRV32Config.fir@6977.4]
  wire [9:0] _T_975; // @[Arbiter.scala 103:44:freechips.rocketchip.system.DefaultRV32Config.fir@6977.4]
  wire [9:0] _GEN_23; // @[Arbiter.scala 103:44:freechips.rocketchip.system.DefaultRV32Config.fir@6978.4]
  wire [9:0] _T_976; // @[Arbiter.scala 103:44:freechips.rocketchip.system.DefaultRV32Config.fir@6978.4]
  wire  _T_993; // @[Mux.scala 27:72:freechips.rocketchip.system.DefaultRV32Config.fir@7005.4]
  wire  _T_994; // @[Mux.scala 27:72:freechips.rocketchip.system.DefaultRV32Config.fir@7006.4]
  wire  _T_996; // @[Mux.scala 27:72:freechips.rocketchip.system.DefaultRV32Config.fir@7008.4]
  wire  _T_995; // @[Mux.scala 27:72:freechips.rocketchip.system.DefaultRV32Config.fir@7007.4]
  wire  _T_997; // @[Mux.scala 27:72:freechips.rocketchip.system.DefaultRV32Config.fir@7009.4]
  wire  _T_999; // @[Arbiter.scala 116:29:freechips.rocketchip.system.DefaultRV32Config.fir@7012.4]
  wire  _T_979; // @[ReadyValidCancel.scala 52:33:freechips.rocketchip.system.DefaultRV32Config.fir@6981.4]
  wire [9:0] _GEN_24; // @[Arbiter.scala 104:52:freechips.rocketchip.system.DefaultRV32Config.fir@6982.4]
  wire [9:0] _T_981; // @[Arbiter.scala 104:52:freechips.rocketchip.system.DefaultRV32Config.fir@6983.4]
  wire  _T_1056; // @[Arbiter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@7187.4]
  wire  _T_1086; // @[Arbiter.scala 26:27:freechips.rocketchip.system.DefaultRV32Config.fir@7221.4]
  wire  _T_1087; // @[Arbiter.scala 26:18:freechips.rocketchip.system.DefaultRV32Config.fir@7222.4]
  wire [2:0] _T_1088; // @[Arbiter.scala 27:29:freechips.rocketchip.system.DefaultRV32Config.fir@7224.6]
  wire [3:0] _T_1089; // @[package.scala 217:48:freechips.rocketchip.system.DefaultRV32Config.fir@7225.6]
  wire [2:0] _T_1091; // @[package.scala 217:43:freechips.rocketchip.system.DefaultRV32Config.fir@7227.6]
  wire [4:0] _T_1092; // @[package.scala 217:48:freechips.rocketchip.system.DefaultRV32Config.fir@7228.6]
  wire [2:0] _T_1094; // @[package.scala 217:43:freechips.rocketchip.system.DefaultRV32Config.fir@7230.6]
  wire  _T_1110; // @[Arbiter.scala 95:53:freechips.rocketchip.system.DefaultRV32Config.fir@7257.4]
  wire  _T_1111; // @[Arbiter.scala 95:53:freechips.rocketchip.system.DefaultRV32Config.fir@7258.4]
  wire  _T_1113; // @[Arbiter.scala 96:67:freechips.rocketchip.system.DefaultRV32Config.fir@7260.4]
  wire  _T_1116; // @[Arbiter.scala 96:67:freechips.rocketchip.system.DefaultRV32Config.fir@7263.4]
  wire  _T_1117; // @[Arbiter.scala 96:64:freechips.rocketchip.system.DefaultRV32Config.fir@7264.4]
  wire  _T_1118; // @[Arbiter.scala 96:61:freechips.rocketchip.system.DefaultRV32Config.fir@7265.4]
  wire  _T_1119; // @[Arbiter.scala 96:67:freechips.rocketchip.system.DefaultRV32Config.fir@7266.4]
  wire  _T_1120; // @[Arbiter.scala 96:64:freechips.rocketchip.system.DefaultRV32Config.fir@7267.4]
  wire  _T_1122; // @[Arbiter.scala 96:82:freechips.rocketchip.system.DefaultRV32Config.fir@7269.4]
  wire  _T_1124; // @[Arbiter.scala 96:13:freechips.rocketchip.system.DefaultRV32Config.fir@7271.4]
  wire  _T_1125; // @[Arbiter.scala 96:13:freechips.rocketchip.system.DefaultRV32Config.fir@7272.4]
  wire  _T_1126; // @[Arbiter.scala 98:36:freechips.rocketchip.system.DefaultRV32Config.fir@7277.4]
  wire  _T_1127; // @[Arbiter.scala 98:36:freechips.rocketchip.system.DefaultRV32Config.fir@7278.4]
  wire  _T_1128; // @[Arbiter.scala 98:15:freechips.rocketchip.system.DefaultRV32Config.fir@7279.4]
  wire  _T_1131; // @[Arbiter.scala 98:41:freechips.rocketchip.system.DefaultRV32Config.fir@7282.4]
  wire  _T_1133; // @[Arbiter.scala 98:14:freechips.rocketchip.system.DefaultRV32Config.fir@7284.4]
  wire  _T_1134; // @[Arbiter.scala 98:14:freechips.rocketchip.system.DefaultRV32Config.fir@7285.4]
  wire  _T_1140; // @[Arbiter.scala 99:41:freechips.rocketchip.system.DefaultRV32Config.fir@7295.4]
  wire  _T_1142; // @[Arbiter.scala 99:14:freechips.rocketchip.system.DefaultRV32Config.fir@7297.4]
  wire  _T_1143; // @[Arbiter.scala 99:14:freechips.rocketchip.system.DefaultRV32Config.fir@7298.4]
  wire [9:0] _T_1144; // @[Arbiter.scala 102:73:freechips.rocketchip.system.DefaultRV32Config.fir@7303.4]
  wire [3:0] _T_1145; // @[Arbiter.scala 102:73:freechips.rocketchip.system.DefaultRV32Config.fir@7304.4]
  wire [5:0] _T_1146; // @[Arbiter.scala 102:73:freechips.rocketchip.system.DefaultRV32Config.fir@7305.4]
  wire [9:0] _GEN_25; // @[Arbiter.scala 103:44:freechips.rocketchip.system.DefaultRV32Config.fir@7306.4]
  wire [9:0] _T_1147; // @[Arbiter.scala 103:44:freechips.rocketchip.system.DefaultRV32Config.fir@7306.4]
  wire [9:0] _GEN_26; // @[Arbiter.scala 103:44:freechips.rocketchip.system.DefaultRV32Config.fir@7307.4]
  wire [9:0] _T_1148; // @[Arbiter.scala 103:44:freechips.rocketchip.system.DefaultRV32Config.fir@7307.4]
  wire  _T_1165; // @[Mux.scala 27:72:freechips.rocketchip.system.DefaultRV32Config.fir@7334.4]
  wire  _T_1166; // @[Mux.scala 27:72:freechips.rocketchip.system.DefaultRV32Config.fir@7335.4]
  wire  _T_1168; // @[Mux.scala 27:72:freechips.rocketchip.system.DefaultRV32Config.fir@7337.4]
  wire  _T_1167; // @[Mux.scala 27:72:freechips.rocketchip.system.DefaultRV32Config.fir@7336.4]
  wire  _T_1169; // @[Mux.scala 27:72:freechips.rocketchip.system.DefaultRV32Config.fir@7338.4]
  wire  _T_1171; // @[Arbiter.scala 116:29:freechips.rocketchip.system.DefaultRV32Config.fir@7341.4]
  wire  _T_1151; // @[ReadyValidCancel.scala 52:33:freechips.rocketchip.system.DefaultRV32Config.fir@7310.4]
  wire [9:0] _GEN_27; // @[Arbiter.scala 104:52:freechips.rocketchip.system.DefaultRV32Config.fir@7311.4]
  wire [9:0] _T_1153; // @[Arbiter.scala 104:52:freechips.rocketchip.system.DefaultRV32Config.fir@7312.4]
  TLMonitor TLMonitor ( // @[Nodes.scala 25:25:freechips.rocketchip.system.DefaultRV32Config.fir@4804.4]
    .clock(TLMonitor_clock),
    .reset(TLMonitor_reset),
    .io_in_a_ready(TLMonitor_io_in_a_ready),
    .io_in_a_valid(TLMonitor_io_in_a_valid),
    .io_in_a_bits_opcode(TLMonitor_io_in_a_bits_opcode),
    .io_in_a_bits_param(TLMonitor_io_in_a_bits_param),
    .io_in_a_bits_size(TLMonitor_io_in_a_bits_size),
    .io_in_a_bits_source(TLMonitor_io_in_a_bits_source),
    .io_in_a_bits_address(TLMonitor_io_in_a_bits_address),
    .io_in_a_bits_mask(TLMonitor_io_in_a_bits_mask),
    .io_in_a_bits_corrupt(TLMonitor_io_in_a_bits_corrupt),
    .io_in_d_ready(TLMonitor_io_in_d_ready),
    .io_in_d_valid(TLMonitor_io_in_d_valid),
    .io_in_d_bits_opcode(TLMonitor_io_in_d_bits_opcode),
    .io_in_d_bits_param(TLMonitor_io_in_d_bits_param),
    .io_in_d_bits_size(TLMonitor_io_in_d_bits_size),
    .io_in_d_bits_source(TLMonitor_io_in_d_bits_source),
    .io_in_d_bits_sink(TLMonitor_io_in_d_bits_sink),
    .io_in_d_bits_denied(TLMonitor_io_in_d_bits_denied),
    .io_in_d_bits_corrupt(TLMonitor_io_in_d_bits_corrupt)
  );
  TLMonitor_1 TLMonitor_1 ( // @[Nodes.scala 25:25:freechips.rocketchip.system.DefaultRV32Config.fir@4834.4]
    .clock(TLMonitor_1_clock),
    .reset(TLMonitor_1_reset),
    .io_in_a_ready(TLMonitor_1_io_in_a_ready),
    .io_in_a_valid(TLMonitor_1_io_in_a_valid),
    .io_in_a_bits_opcode(TLMonitor_1_io_in_a_bits_opcode),
    .io_in_a_bits_param(TLMonitor_1_io_in_a_bits_param),
    .io_in_a_bits_size(TLMonitor_1_io_in_a_bits_size),
    .io_in_a_bits_source(TLMonitor_1_io_in_a_bits_source),
    .io_in_a_bits_address(TLMonitor_1_io_in_a_bits_address),
    .io_in_a_bits_mask(TLMonitor_1_io_in_a_bits_mask),
    .io_in_a_bits_corrupt(TLMonitor_1_io_in_a_bits_corrupt),
    .io_in_b_ready(TLMonitor_1_io_in_b_ready),
    .io_in_b_valid(TLMonitor_1_io_in_b_valid),
    .io_in_b_bits_param(TLMonitor_1_io_in_b_bits_param),
    .io_in_b_bits_address(TLMonitor_1_io_in_b_bits_address),
    .io_in_c_ready(TLMonitor_1_io_in_c_ready),
    .io_in_c_valid(TLMonitor_1_io_in_c_valid),
    .io_in_c_bits_opcode(TLMonitor_1_io_in_c_bits_opcode),
    .io_in_c_bits_param(TLMonitor_1_io_in_c_bits_param),
    .io_in_c_bits_size(TLMonitor_1_io_in_c_bits_size),
    .io_in_c_bits_source(TLMonitor_1_io_in_c_bits_source),
    .io_in_c_bits_address(TLMonitor_1_io_in_c_bits_address),
    .io_in_c_bits_corrupt(TLMonitor_1_io_in_c_bits_corrupt),
    .io_in_d_ready(TLMonitor_1_io_in_d_ready),
    .io_in_d_valid(TLMonitor_1_io_in_d_valid),
    .io_in_d_bits_opcode(TLMonitor_1_io_in_d_bits_opcode),
    .io_in_d_bits_param(TLMonitor_1_io_in_d_bits_param),
    .io_in_d_bits_size(TLMonitor_1_io_in_d_bits_size),
    .io_in_d_bits_source(TLMonitor_1_io_in_d_bits_source),
    .io_in_d_bits_sink(TLMonitor_1_io_in_d_bits_sink),
    .io_in_d_bits_denied(TLMonitor_1_io_in_d_bits_denied),
    .io_in_d_bits_corrupt(TLMonitor_1_io_in_d_bits_corrupt),
    .io_in_e_valid(TLMonitor_1_io_in_e_valid),
    .io_in_e_bits_sink(TLMonitor_1_io_in_e_bits_sink)
  );
  assign _T_883 = _T_882 == 10'h0; // @[Arbiter.scala 79:28:freechips.rocketchip.system.DefaultRV32Config.fir@6857.4]
  assign _T_180 = ~auto_out_2_d_bits_source[4]; // @[Parameters.scala 55:32:freechips.rocketchip.system.DefaultRV32Config.fir@5462.4]
  assign _T_383 = auto_out_2_d_valid & _T_180; // @[Xbar.scala 173:40:freechips.rocketchip.system.DefaultRV32Config.fir@5931.4]
  assign _T_164 = ~auto_out_1_d_bits_source[4]; // @[Parameters.scala 55:32:freechips.rocketchip.system.DefaultRV32Config.fir@5446.4]
  assign _T_374 = auto_out_1_d_valid & _T_164; // @[Xbar.scala 173:40:freechips.rocketchip.system.DefaultRV32Config.fir@5902.4]
  assign _T_148 = ~auto_out_0_d_bits_source[4]; // @[Parameters.scala 55:32:freechips.rocketchip.system.DefaultRV32Config.fir@5430.4]
  assign _T_365 = auto_out_0_d_valid & _T_148; // @[Xbar.scala 173:40:freechips.rocketchip.system.DefaultRV32Config.fir@5873.4]
  assign _T_892 = {_T_383,_T_374,_T_365}; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@6866.4]
  assign _T_899 = ~_T_898; // @[Arbiter.scala 23:30:freechips.rocketchip.system.DefaultRV32Config.fir@6877.4]
  assign _T_900 = _T_892 & _T_899; // @[Arbiter.scala 23:28:freechips.rocketchip.system.DefaultRV32Config.fir@6878.4]
  assign _T_901 = {_T_900,_T_383,_T_374,_T_365}; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@6879.4]
  assign _GEN_5 = {{1'd0}, _T_901[5:1]}; // @[package.scala 226:43:freechips.rocketchip.system.DefaultRV32Config.fir@6881.4]
  assign _T_903 = _T_901 | _GEN_5; // @[package.scala 226:43:freechips.rocketchip.system.DefaultRV32Config.fir@6881.4]
  assign _GEN_6 = {{2'd0}, _T_903[5:2]}; // @[package.scala 226:43:freechips.rocketchip.system.DefaultRV32Config.fir@6883.4]
  assign _T_905 = _T_903 | _GEN_6; // @[package.scala 226:43:freechips.rocketchip.system.DefaultRV32Config.fir@6883.4]
  assign _T_908 = {_T_898, 3'h0}; // @[Arbiter.scala 24:66:freechips.rocketchip.system.DefaultRV32Config.fir@6886.4]
  assign _GEN_7 = {{1'd0}, _T_905[5:1]}; // @[Arbiter.scala 24:58:freechips.rocketchip.system.DefaultRV32Config.fir@6887.4]
  assign _T_909 = _GEN_7 | _T_908; // @[Arbiter.scala 24:58:freechips.rocketchip.system.DefaultRV32Config.fir@6887.4]
  assign _T_912 = _T_909[5:3] & _T_909[2:0]; // @[Arbiter.scala 25:39:freechips.rocketchip.system.DefaultRV32Config.fir@6890.4]
  assign _T_913 = ~_T_912; // @[Arbiter.scala 25:18:freechips.rocketchip.system.DefaultRV32Config.fir@6891.4]
  assign _T_929 = _T_913[0] & _T_365; // @[Arbiter.scala 88:79:freechips.rocketchip.system.DefaultRV32Config.fir@6913.4]
  assign _T_985_0 = _T_883 ? _T_929 : _T_984_0; // @[Arbiter.scala 108:30:freechips.rocketchip.system.DefaultRV32Config.fir@6991.4]
  assign _T_20_0_d_bits_sink = {{1'd0}, auto_out_0_d_bits_sink}; // @[Xbar.scala 282:19:freechips.rocketchip.system.DefaultRV32Config.fir@5123.4 BundleMap.scala 248:19:freechips.rocketchip.system.DefaultRV32Config.fir@5172.4 Xbar.scala 317:28:freechips.rocketchip.system.DefaultRV32Config.fir@5180.4]
  assign _T_1012 = {auto_out_0_d_bits_opcode,auto_out_0_d_bits_param,auto_out_0_d_bits_size,auto_out_0_d_bits_source,_T_20_0_d_bits_sink,auto_out_0_d_bits_denied,auto_out_0_d_bits_data,auto_out_0_d_bits_corrupt}; // @[Mux.scala 27:72:freechips.rocketchip.system.DefaultRV32Config.fir@7028.4]
  assign _T_1013 = _T_985_0 ? _T_1012 : 50'h0; // @[Mux.scala 27:72:freechips.rocketchip.system.DefaultRV32Config.fir@7029.4]
  assign _T_930 = _T_913[1] & _T_374; // @[Arbiter.scala 88:79:freechips.rocketchip.system.DefaultRV32Config.fir@6914.4]
  assign _T_985_1 = _T_883 ? _T_930 : _T_984_1; // @[Arbiter.scala 108:30:freechips.rocketchip.system.DefaultRV32Config.fir@6991.4]
  assign _T_20_1_d_bits_size = {{1'd0}, auto_out_1_d_bits_size}; // @[Xbar.scala 282:19:freechips.rocketchip.system.DefaultRV32Config.fir@5123.4 BundleMap.scala 248:19:freechips.rocketchip.system.DefaultRV32Config.fir@5227.4]
  assign _T_1020 = {auto_out_1_d_bits_opcode,auto_out_1_d_bits_param,_T_20_1_d_bits_size,auto_out_1_d_bits_source,auto_out_1_d_bits_sink,auto_out_1_d_bits_denied,auto_out_1_d_bits_data,auto_out_1_d_bits_corrupt}; // @[Mux.scala 27:72:freechips.rocketchip.system.DefaultRV32Config.fir@7036.4]
  assign _T_1021 = _T_985_1 ? _T_1020 : 50'h0; // @[Mux.scala 27:72:freechips.rocketchip.system.DefaultRV32Config.fir@7037.4]
  assign _T_1030 = _T_1013 | _T_1021; // @[Mux.scala 27:72:freechips.rocketchip.system.DefaultRV32Config.fir@7046.4]
  assign _T_931 = _T_913[2] & _T_383; // @[Arbiter.scala 88:79:freechips.rocketchip.system.DefaultRV32Config.fir@6915.4]
  assign _T_985_2 = _T_883 ? _T_931 : _T_984_2; // @[Arbiter.scala 108:30:freechips.rocketchip.system.DefaultRV32Config.fir@6991.4]
  assign _T_1028 = {auto_out_2_d_bits_opcode,2'h0,auto_out_2_d_bits_size,auto_out_2_d_bits_source,2'h0,auto_out_2_d_bits_denied,auto_out_2_d_bits_data,auto_out_2_d_bits_corrupt}; // @[Mux.scala 27:72:freechips.rocketchip.system.DefaultRV32Config.fir@7044.4]
  assign _T_1029 = _T_985_2 ? _T_1028 : 50'h0; // @[Mux.scala 27:72:freechips.rocketchip.system.DefaultRV32Config.fir@7045.4]
  assign _T_1031 = _T_1030 | _T_1029; // @[Mux.scala 27:72:freechips.rocketchip.system.DefaultRV32Config.fir@7047.4]
  assign _GEN_8 = {{3'd0}, auto_in_1_a_bits_source}; // @[Xbar.scala 231:55:freechips.rocketchip.system.DefaultRV32Config.fir@5083.4]
  assign _T_16 = _GEN_8 | 5'h10; // @[Xbar.scala 231:55:freechips.rocketchip.system.DefaultRV32Config.fir@5083.4]
  assign _GEN_9 = {{3'd0}, auto_in_1_c_bits_source}; // @[Xbar.scala 253:55:freechips.rocketchip.system.DefaultRV32Config.fir@5106.4]
  assign _T_1055 = _T_1054 == 10'h0; // @[Arbiter.scala 79:28:freechips.rocketchip.system.DefaultRV32Config.fir@7186.4]
  assign _T_188 = auto_out_2_d_bits_source[4:2] == 3'h4; // @[Parameters.scala 55:32:freechips.rocketchip.system.DefaultRV32Config.fir@5470.4]
  assign _T_385 = auto_out_2_d_valid & _T_188; // @[Xbar.scala 173:40:freechips.rocketchip.system.DefaultRV32Config.fir@5942.4]
  assign _T_172 = auto_out_1_d_bits_source[4:2] == 3'h4; // @[Parameters.scala 55:32:freechips.rocketchip.system.DefaultRV32Config.fir@5454.4]
  assign _T_376 = auto_out_1_d_valid & _T_172; // @[Xbar.scala 173:40:freechips.rocketchip.system.DefaultRV32Config.fir@5913.4]
  assign _T_156 = auto_out_0_d_bits_source[4:2] == 3'h4; // @[Parameters.scala 55:32:freechips.rocketchip.system.DefaultRV32Config.fir@5438.4]
  assign _T_367 = auto_out_0_d_valid & _T_156; // @[Xbar.scala 173:40:freechips.rocketchip.system.DefaultRV32Config.fir@5884.4]
  assign _T_1064 = {_T_385,_T_376,_T_367}; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@7195.4]
  assign _T_1071 = ~_T_1070; // @[Arbiter.scala 23:30:freechips.rocketchip.system.DefaultRV32Config.fir@7206.4]
  assign _T_1072 = _T_1064 & _T_1071; // @[Arbiter.scala 23:28:freechips.rocketchip.system.DefaultRV32Config.fir@7207.4]
  assign _T_1073 = {_T_1072,_T_385,_T_376,_T_367}; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@7208.4]
  assign _GEN_10 = {{1'd0}, _T_1073[5:1]}; // @[package.scala 226:43:freechips.rocketchip.system.DefaultRV32Config.fir@7210.4]
  assign _T_1075 = _T_1073 | _GEN_10; // @[package.scala 226:43:freechips.rocketchip.system.DefaultRV32Config.fir@7210.4]
  assign _GEN_11 = {{2'd0}, _T_1075[5:2]}; // @[package.scala 226:43:freechips.rocketchip.system.DefaultRV32Config.fir@7212.4]
  assign _T_1077 = _T_1075 | _GEN_11; // @[package.scala 226:43:freechips.rocketchip.system.DefaultRV32Config.fir@7212.4]
  assign _T_1080 = {_T_1070, 3'h0}; // @[Arbiter.scala 24:66:freechips.rocketchip.system.DefaultRV32Config.fir@7215.4]
  assign _GEN_12 = {{1'd0}, _T_1077[5:1]}; // @[Arbiter.scala 24:58:freechips.rocketchip.system.DefaultRV32Config.fir@7216.4]
  assign _T_1081 = _GEN_12 | _T_1080; // @[Arbiter.scala 24:58:freechips.rocketchip.system.DefaultRV32Config.fir@7216.4]
  assign _T_1084 = _T_1081[5:3] & _T_1081[2:0]; // @[Arbiter.scala 25:39:freechips.rocketchip.system.DefaultRV32Config.fir@7219.4]
  assign _T_1085 = ~_T_1084; // @[Arbiter.scala 25:18:freechips.rocketchip.system.DefaultRV32Config.fir@7220.4]
  assign _T_1101 = _T_1085[0] & _T_367; // @[Arbiter.scala 88:79:freechips.rocketchip.system.DefaultRV32Config.fir@7242.4]
  assign _T_1157_0 = _T_1055 ? _T_1101 : _T_1156_0; // @[Arbiter.scala 108:30:freechips.rocketchip.system.DefaultRV32Config.fir@7320.4]
  assign _T_1185 = _T_1157_0 ? _T_1012 : 50'h0; // @[Mux.scala 27:72:freechips.rocketchip.system.DefaultRV32Config.fir@7358.4]
  assign _T_1102 = _T_1085[1] & _T_376; // @[Arbiter.scala 88:79:freechips.rocketchip.system.DefaultRV32Config.fir@7243.4]
  assign _T_1157_1 = _T_1055 ? _T_1102 : _T_1156_1; // @[Arbiter.scala 108:30:freechips.rocketchip.system.DefaultRV32Config.fir@7320.4]
  assign _T_1193 = _T_1157_1 ? _T_1020 : 50'h0; // @[Mux.scala 27:72:freechips.rocketchip.system.DefaultRV32Config.fir@7366.4]
  assign _T_1202 = _T_1185 | _T_1193; // @[Mux.scala 27:72:freechips.rocketchip.system.DefaultRV32Config.fir@7375.4]
  assign _T_1103 = _T_1085[2] & _T_385; // @[Arbiter.scala 88:79:freechips.rocketchip.system.DefaultRV32Config.fir@7244.4]
  assign _T_1157_2 = _T_1055 ? _T_1103 : _T_1156_2; // @[Arbiter.scala 108:30:freechips.rocketchip.system.DefaultRV32Config.fir@7320.4]
  assign _T_1201 = _T_1157_2 ? _T_1028 : 50'h0; // @[Mux.scala 27:72:freechips.rocketchip.system.DefaultRV32Config.fir@7374.4]
  assign _T_1203 = _T_1202 | _T_1201; // @[Mux.scala 27:72:freechips.rocketchip.system.DefaultRV32Config.fir@7376.4]
  assign _T_26 = {1'b0,$signed(auto_in_0_a_bits_address)}; // @[Parameters.scala 137:49:freechips.rocketchip.system.DefaultRV32Config.fir@5308.4]
  assign _T_28 = $signed(_T_26) & 33'shc0000000; // @[Parameters.scala 137:52:freechips.rocketchip.system.DefaultRV32Config.fir@5310.4]
  assign _T_29 = $signed(_T_28) == 33'sh0; // @[Parameters.scala 137:67:freechips.rocketchip.system.DefaultRV32Config.fir@5311.4]
  assign _T_31 = auto_in_0_a_bits_address ^ 32'h80000000; // @[Parameters.scala 137:31:freechips.rocketchip.system.DefaultRV32Config.fir@5313.4]
  assign _T_32 = {1'b0,$signed(_T_31)}; // @[Parameters.scala 137:49:freechips.rocketchip.system.DefaultRV32Config.fir@5314.4]
  assign _T_34 = $signed(_T_32) & 33'shc0000000; // @[Parameters.scala 137:52:freechips.rocketchip.system.DefaultRV32Config.fir@5316.4]
  assign _T_35 = $signed(_T_34) == 33'sh0; // @[Parameters.scala 137:67:freechips.rocketchip.system.DefaultRV32Config.fir@5317.4]
  assign _T_37 = auto_in_0_a_bits_address ^ 32'h40000000; // @[Parameters.scala 137:31:freechips.rocketchip.system.DefaultRV32Config.fir@5319.4]
  assign _T_38 = {1'b0,$signed(_T_37)}; // @[Parameters.scala 137:49:freechips.rocketchip.system.DefaultRV32Config.fir@5320.4]
  assign _T_40 = $signed(_T_38) & 33'shc0000000; // @[Parameters.scala 137:52:freechips.rocketchip.system.DefaultRV32Config.fir@5322.4]
  assign _T_41 = $signed(_T_40) == 33'sh0; // @[Parameters.scala 137:67:freechips.rocketchip.system.DefaultRV32Config.fir@5323.4]
  assign _T_44 = {1'b0,$signed(auto_in_1_a_bits_address)}; // @[Parameters.scala 137:49:freechips.rocketchip.system.DefaultRV32Config.fir@5326.4]
  assign _T_46 = $signed(_T_44) & 33'shc0000000; // @[Parameters.scala 137:52:freechips.rocketchip.system.DefaultRV32Config.fir@5328.4]
  assign _T_47 = $signed(_T_46) == 33'sh0; // @[Parameters.scala 137:67:freechips.rocketchip.system.DefaultRV32Config.fir@5329.4]
  assign _T_49 = auto_in_1_a_bits_address ^ 32'h80000000; // @[Parameters.scala 137:31:freechips.rocketchip.system.DefaultRV32Config.fir@5331.4]
  assign _T_50 = {1'b0,$signed(_T_49)}; // @[Parameters.scala 137:49:freechips.rocketchip.system.DefaultRV32Config.fir@5332.4]
  assign _T_52 = $signed(_T_50) & 33'shc0000000; // @[Parameters.scala 137:52:freechips.rocketchip.system.DefaultRV32Config.fir@5334.4]
  assign _T_53 = $signed(_T_52) == 33'sh0; // @[Parameters.scala 137:67:freechips.rocketchip.system.DefaultRV32Config.fir@5335.4]
  assign _T_55 = auto_in_1_a_bits_address ^ 32'h40000000; // @[Parameters.scala 137:31:freechips.rocketchip.system.DefaultRV32Config.fir@5337.4]
  assign _T_56 = {1'b0,$signed(_T_55)}; // @[Parameters.scala 137:49:freechips.rocketchip.system.DefaultRV32Config.fir@5338.4]
  assign _T_58 = $signed(_T_56) & 33'shc0000000; // @[Parameters.scala 137:52:freechips.rocketchip.system.DefaultRV32Config.fir@5340.4]
  assign _T_59 = $signed(_T_58) == 33'sh0; // @[Parameters.scala 137:67:freechips.rocketchip.system.DefaultRV32Config.fir@5341.4]
  assign _T_210 = 27'hfff << auto_in_0_a_bits_size; // @[package.scala 207:77:freechips.rocketchip.system.DefaultRV32Config.fir@5492.4]
  assign _T_212 = ~_T_210[11:0]; // @[package.scala 207:46:freechips.rocketchip.system.DefaultRV32Config.fir@5494.4]
  assign _T_215 = ~auto_in_0_a_bits_opcode[2]; // @[Edges.scala 93:28:freechips.rocketchip.system.DefaultRV32Config.fir@5497.4]
  assign _T_216 = _T_215 ? _T_212[11:2] : 10'h0; // @[Edges.scala 222:14:freechips.rocketchip.system.DefaultRV32Config.fir@5498.4]
  assign _T_218 = 27'hfff << auto_in_1_a_bits_size; // @[package.scala 207:77:freechips.rocketchip.system.DefaultRV32Config.fir@5500.4]
  assign _T_220 = ~_T_218[11:0]; // @[package.scala 207:46:freechips.rocketchip.system.DefaultRV32Config.fir@5502.4]
  assign _T_223 = ~auto_in_1_a_bits_opcode[2]; // @[Edges.scala 93:28:freechips.rocketchip.system.DefaultRV32Config.fir@5505.4]
  assign _T_224 = _T_223 ? _T_220[11:2] : 10'h0; // @[Edges.scala 222:14:freechips.rocketchip.system.DefaultRV32Config.fir@5506.4]
  assign _T_264 = 27'hfff << auto_out_0_d_bits_size; // @[package.scala 207:77:freechips.rocketchip.system.DefaultRV32Config.fir@5546.4]
  assign _T_266 = ~_T_264[11:0]; // @[package.scala 207:46:freechips.rocketchip.system.DefaultRV32Config.fir@5548.4]
  assign _T_269 = auto_out_0_d_bits_opcode[0] ? _T_266[11:2] : 10'h0; // @[Edges.scala 222:14:freechips.rocketchip.system.DefaultRV32Config.fir@5551.4]
  assign _T_271 = 21'h3f << _T_20_1_d_bits_size; // @[package.scala 207:77:freechips.rocketchip.system.DefaultRV32Config.fir@5553.4]
  assign _T_273 = ~_T_271[5:0]; // @[package.scala 207:46:freechips.rocketchip.system.DefaultRV32Config.fir@5555.4]
  assign _T_276 = auto_out_1_d_bits_opcode[0] ? _T_273[5:2] : 4'h0; // @[Edges.scala 222:14:freechips.rocketchip.system.DefaultRV32Config.fir@5558.4]
  assign _T_278 = 23'hff << auto_out_2_d_bits_size; // @[package.scala 207:77:freechips.rocketchip.system.DefaultRV32Config.fir@5560.4]
  assign _T_280 = ~_T_278[7:0]; // @[package.scala 207:46:freechips.rocketchip.system.DefaultRV32Config.fir@5562.4]
  assign _T_283 = auto_out_2_d_bits_opcode[0] ? _T_280[7:2] : 6'h0; // @[Edges.scala 222:14:freechips.rocketchip.system.DefaultRV32Config.fir@5565.4]
  assign _T_286 = auto_in_0_a_valid & _T_29; // @[Xbar.scala 422:50:freechips.rocketchip.system.DefaultRV32Config.fir@5584.4]
  assign _T_288 = auto_in_0_a_valid & _T_35; // @[Xbar.scala 422:50:freechips.rocketchip.system.DefaultRV32Config.fir@5603.4]
  assign _T_290 = auto_in_0_a_valid & _T_41; // @[Xbar.scala 422:50:freechips.rocketchip.system.DefaultRV32Config.fir@5622.4]
  assign _T_417 = _T_416 == 10'h0; // @[Arbiter.scala 79:28:freechips.rocketchip.system.DefaultRV32Config.fir@5993.4]
  assign _T_299 = auto_in_1_a_valid & _T_47; // @[Xbar.scala 422:50:freechips.rocketchip.system.DefaultRV32Config.fir@5650.4]
  assign _T_423 = {_T_299,_T_286}; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@5999.4]
  assign _T_430 = ~_T_429; // @[Arbiter.scala 23:30:freechips.rocketchip.system.DefaultRV32Config.fir@6010.4]
  assign _T_431 = _T_423 & _T_430; // @[Arbiter.scala 23:28:freechips.rocketchip.system.DefaultRV32Config.fir@6011.4]
  assign _T_432 = {_T_431,_T_299,_T_286}; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@6012.4]
  assign _GEN_13 = {{1'd0}, _T_432[3:1]}; // @[package.scala 226:43:freechips.rocketchip.system.DefaultRV32Config.fir@6014.4]
  assign _T_434 = _T_432 | _GEN_13; // @[package.scala 226:43:freechips.rocketchip.system.DefaultRV32Config.fir@6014.4]
  assign _T_437 = {_T_429, 2'h0}; // @[Arbiter.scala 24:66:freechips.rocketchip.system.DefaultRV32Config.fir@6017.4]
  assign _GEN_14 = {{1'd0}, _T_434[3:1]}; // @[Arbiter.scala 24:58:freechips.rocketchip.system.DefaultRV32Config.fir@6018.4]
  assign _T_438 = _GEN_14 | _T_437; // @[Arbiter.scala 24:58:freechips.rocketchip.system.DefaultRV32Config.fir@6018.4]
  assign _T_441 = _T_438[3:2] & _T_438[1:0]; // @[Arbiter.scala 25:39:freechips.rocketchip.system.DefaultRV32Config.fir@6021.4]
  assign _T_442 = ~_T_441; // @[Arbiter.scala 25:18:freechips.rocketchip.system.DefaultRV32Config.fir@6022.4]
  assign _T_499_0 = _T_417 ? _T_442[0] : _T_496_0; // @[Arbiter.scala 112:24:freechips.rocketchip.system.DefaultRV32Config.fir@6105.4]
  assign _T_500 = auto_out_0_a_ready & _T_499_0; // @[Arbiter.scala 114:31:freechips.rocketchip.system.DefaultRV32Config.fir@6106.4]
  assign _T_291 = _T_29 & _T_500; // @[Mux.scala 27:72:freechips.rocketchip.system.DefaultRV32Config.fir@5624.4]
  assign _T_569 = _T_568 == 10'h0; // @[Arbiter.scala 79:28:freechips.rocketchip.system.DefaultRV32Config.fir@6252.4]
  assign _T_301 = auto_in_1_a_valid & _T_53; // @[Xbar.scala 422:50:freechips.rocketchip.system.DefaultRV32Config.fir@5669.4]
  assign _T_575 = {_T_301,_T_288}; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@6258.4]
  assign _T_582 = ~_T_581; // @[Arbiter.scala 23:30:freechips.rocketchip.system.DefaultRV32Config.fir@6269.4]
  assign _T_583 = _T_575 & _T_582; // @[Arbiter.scala 23:28:freechips.rocketchip.system.DefaultRV32Config.fir@6270.4]
  assign _T_584 = {_T_583,_T_301,_T_288}; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@6271.4]
  assign _GEN_15 = {{1'd0}, _T_584[3:1]}; // @[package.scala 226:43:freechips.rocketchip.system.DefaultRV32Config.fir@6273.4]
  assign _T_586 = _T_584 | _GEN_15; // @[package.scala 226:43:freechips.rocketchip.system.DefaultRV32Config.fir@6273.4]
  assign _T_589 = {_T_581, 2'h0}; // @[Arbiter.scala 24:66:freechips.rocketchip.system.DefaultRV32Config.fir@6276.4]
  assign _GEN_16 = {{1'd0}, _T_586[3:1]}; // @[Arbiter.scala 24:58:freechips.rocketchip.system.DefaultRV32Config.fir@6277.4]
  assign _T_590 = _GEN_16 | _T_589; // @[Arbiter.scala 24:58:freechips.rocketchip.system.DefaultRV32Config.fir@6277.4]
  assign _T_593 = _T_590[3:2] & _T_590[1:0]; // @[Arbiter.scala 25:39:freechips.rocketchip.system.DefaultRV32Config.fir@6280.4]
  assign _T_594 = ~_T_593; // @[Arbiter.scala 25:18:freechips.rocketchip.system.DefaultRV32Config.fir@6281.4]
  assign _T_651_0 = _T_569 ? _T_594[0] : _T_648_0; // @[Arbiter.scala 112:24:freechips.rocketchip.system.DefaultRV32Config.fir@6364.4]
  assign _T_652 = auto_out_1_a_ready & _T_651_0; // @[Arbiter.scala 114:31:freechips.rocketchip.system.DefaultRV32Config.fir@6365.4]
  assign _T_292 = _T_35 & _T_652; // @[Mux.scala 27:72:freechips.rocketchip.system.DefaultRV32Config.fir@5625.4]
  assign _T_723 = _T_722 == 10'h0; // @[Arbiter.scala 79:28:freechips.rocketchip.system.DefaultRV32Config.fir@6527.4]
  assign _T_303 = auto_in_1_a_valid & _T_59; // @[Xbar.scala 422:50:freechips.rocketchip.system.DefaultRV32Config.fir@5688.4]
  assign _T_729 = {_T_303,_T_290}; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@6533.4]
  assign _T_736 = ~_T_735; // @[Arbiter.scala 23:30:freechips.rocketchip.system.DefaultRV32Config.fir@6544.4]
  assign _T_737 = _T_729 & _T_736; // @[Arbiter.scala 23:28:freechips.rocketchip.system.DefaultRV32Config.fir@6545.4]
  assign _T_738 = {_T_737,_T_303,_T_290}; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@6546.4]
  assign _GEN_17 = {{1'd0}, _T_738[3:1]}; // @[package.scala 226:43:freechips.rocketchip.system.DefaultRV32Config.fir@6548.4]
  assign _T_740 = _T_738 | _GEN_17; // @[package.scala 226:43:freechips.rocketchip.system.DefaultRV32Config.fir@6548.4]
  assign _T_743 = {_T_735, 2'h0}; // @[Arbiter.scala 24:66:freechips.rocketchip.system.DefaultRV32Config.fir@6551.4]
  assign _GEN_18 = {{1'd0}, _T_740[3:1]}; // @[Arbiter.scala 24:58:freechips.rocketchip.system.DefaultRV32Config.fir@6552.4]
  assign _T_744 = _GEN_18 | _T_743; // @[Arbiter.scala 24:58:freechips.rocketchip.system.DefaultRV32Config.fir@6552.4]
  assign _T_747 = _T_744[3:2] & _T_744[1:0]; // @[Arbiter.scala 25:39:freechips.rocketchip.system.DefaultRV32Config.fir@6555.4]
  assign _T_748 = ~_T_747; // @[Arbiter.scala 25:18:freechips.rocketchip.system.DefaultRV32Config.fir@6556.4]
  assign _T_805_0 = _T_723 ? _T_748[0] : _T_802_0; // @[Arbiter.scala 112:24:freechips.rocketchip.system.DefaultRV32Config.fir@6639.4]
  assign _T_806 = auto_out_2_a_ready & _T_805_0; // @[Arbiter.scala 114:31:freechips.rocketchip.system.DefaultRV32Config.fir@6640.4]
  assign _T_293 = _T_41 & _T_806; // @[Mux.scala 27:72:freechips.rocketchip.system.DefaultRV32Config.fir@5626.4]
  assign _T_294 = _T_291 | _T_292; // @[Mux.scala 27:72:freechips.rocketchip.system.DefaultRV32Config.fir@5627.4]
  assign _T_499_1 = _T_417 ? _T_442[1] : _T_496_1; // @[Arbiter.scala 112:24:freechips.rocketchip.system.DefaultRV32Config.fir@6105.4]
  assign _T_501 = auto_out_0_a_ready & _T_499_1; // @[Arbiter.scala 114:31:freechips.rocketchip.system.DefaultRV32Config.fir@6108.4]
  assign _T_304 = _T_47 & _T_501; // @[Mux.scala 27:72:freechips.rocketchip.system.DefaultRV32Config.fir@5690.4]
  assign _T_651_1 = _T_569 ? _T_594[1] : _T_648_1; // @[Arbiter.scala 112:24:freechips.rocketchip.system.DefaultRV32Config.fir@6364.4]
  assign _T_653 = auto_out_1_a_ready & _T_651_1; // @[Arbiter.scala 114:31:freechips.rocketchip.system.DefaultRV32Config.fir@6367.4]
  assign _T_305 = _T_53 & _T_653; // @[Mux.scala 27:72:freechips.rocketchip.system.DefaultRV32Config.fir@5691.4]
  assign _T_805_1 = _T_723 ? _T_748[1] : _T_802_1; // @[Arbiter.scala 112:24:freechips.rocketchip.system.DefaultRV32Config.fir@6639.4]
  assign _T_807 = auto_out_2_a_ready & _T_805_1; // @[Arbiter.scala 114:31:freechips.rocketchip.system.DefaultRV32Config.fir@6642.4]
  assign _T_306 = _T_59 & _T_807; // @[Mux.scala 27:72:freechips.rocketchip.system.DefaultRV32Config.fir@5692.4]
  assign _T_307 = _T_304 | _T_305; // @[Mux.scala 27:72:freechips.rocketchip.system.DefaultRV32Config.fir@5693.4]
  assign _T_987_0 = _T_883 ? _T_913[0] : _T_984_0; // @[Arbiter.scala 112:24:freechips.rocketchip.system.DefaultRV32Config.fir@6996.4]
  assign _T_988 = auto_in_0_d_ready & _T_987_0; // @[Arbiter.scala 114:31:freechips.rocketchip.system.DefaultRV32Config.fir@6997.4]
  assign _T_368 = _T_148 & _T_988; // @[Mux.scala 27:72:freechips.rocketchip.system.DefaultRV32Config.fir@5886.4]
  assign _T_1159_0 = _T_1055 ? _T_1085[0] : _T_1156_0; // @[Arbiter.scala 112:24:freechips.rocketchip.system.DefaultRV32Config.fir@7325.4]
  assign _T_1160 = auto_in_1_d_ready & _T_1159_0; // @[Arbiter.scala 114:31:freechips.rocketchip.system.DefaultRV32Config.fir@7326.4]
  assign _T_369 = _T_156 & _T_1160; // @[Mux.scala 27:72:freechips.rocketchip.system.DefaultRV32Config.fir@5887.4]
  assign _T_987_1 = _T_883 ? _T_913[1] : _T_984_1; // @[Arbiter.scala 112:24:freechips.rocketchip.system.DefaultRV32Config.fir@6996.4]
  assign _T_989 = auto_in_0_d_ready & _T_987_1; // @[Arbiter.scala 114:31:freechips.rocketchip.system.DefaultRV32Config.fir@6999.4]
  assign _T_377 = _T_164 & _T_989; // @[Mux.scala 27:72:freechips.rocketchip.system.DefaultRV32Config.fir@5915.4]
  assign _T_1159_1 = _T_1055 ? _T_1085[1] : _T_1156_1; // @[Arbiter.scala 112:24:freechips.rocketchip.system.DefaultRV32Config.fir@7325.4]
  assign _T_1161 = auto_in_1_d_ready & _T_1159_1; // @[Arbiter.scala 114:31:freechips.rocketchip.system.DefaultRV32Config.fir@7328.4]
  assign _T_378 = _T_172 & _T_1161; // @[Mux.scala 27:72:freechips.rocketchip.system.DefaultRV32Config.fir@5916.4]
  assign _T_987_2 = _T_883 ? _T_913[2] : _T_984_2; // @[Arbiter.scala 112:24:freechips.rocketchip.system.DefaultRV32Config.fir@6996.4]
  assign _T_990 = auto_in_0_d_ready & _T_987_2; // @[Arbiter.scala 114:31:freechips.rocketchip.system.DefaultRV32Config.fir@7001.4]
  assign _T_386 = _T_180 & _T_990; // @[Mux.scala 27:72:freechips.rocketchip.system.DefaultRV32Config.fir@5944.4]
  assign _T_1159_2 = _T_1055 ? _T_1085[2] : _T_1156_2; // @[Arbiter.scala 112:24:freechips.rocketchip.system.DefaultRV32Config.fir@7325.4]
  assign _T_1162 = auto_in_1_d_ready & _T_1159_2; // @[Arbiter.scala 114:31:freechips.rocketchip.system.DefaultRV32Config.fir@7330.4]
  assign _T_387 = _T_188 & _T_1162; // @[Mux.scala 27:72:freechips.rocketchip.system.DefaultRV32Config.fir@5945.4]
  assign _T_418 = _T_417 & auto_out_0_a_ready; // @[Arbiter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@5994.4]
  assign _T_443 = |_T_423; // @[Arbiter.scala 26:27:freechips.rocketchip.system.DefaultRV32Config.fir@6023.4]
  assign _T_444 = _T_418 & _T_443; // @[Arbiter.scala 26:18:freechips.rocketchip.system.DefaultRV32Config.fir@6024.4]
  assign _T_445 = _T_442 & _T_423; // @[Arbiter.scala 27:29:freechips.rocketchip.system.DefaultRV32Config.fir@6026.6]
  assign _T_446 = {_T_445, 1'h0}; // @[package.scala 217:48:freechips.rocketchip.system.DefaultRV32Config.fir@6027.6]
  assign _T_448 = _T_445 | _T_446[1:0]; // @[package.scala 217:43:freechips.rocketchip.system.DefaultRV32Config.fir@6029.6]
  assign _T_454 = _T_442[0] & _T_286; // @[Arbiter.scala 88:79:freechips.rocketchip.system.DefaultRV32Config.fir@6039.4]
  assign _T_455 = _T_442[1] & _T_299; // @[Arbiter.scala 88:79:freechips.rocketchip.system.DefaultRV32Config.fir@6040.4]
  assign _T_461 = _T_454 | _T_455; // @[Arbiter.scala 95:53:freechips.rocketchip.system.DefaultRV32Config.fir@6050.4]
  assign _T_463 = ~_T_454; // @[Arbiter.scala 96:67:freechips.rocketchip.system.DefaultRV32Config.fir@6052.4]
  assign _T_466 = ~_T_455; // @[Arbiter.scala 96:67:freechips.rocketchip.system.DefaultRV32Config.fir@6055.4]
  assign _T_467 = _T_463 | _T_466; // @[Arbiter.scala 96:64:freechips.rocketchip.system.DefaultRV32Config.fir@6056.4]
  assign _T_470 = _T_467 | reset; // @[Arbiter.scala 96:13:freechips.rocketchip.system.DefaultRV32Config.fir@6059.4]
  assign _T_471 = ~_T_470; // @[Arbiter.scala 96:13:freechips.rocketchip.system.DefaultRV32Config.fir@6060.4]
  assign _T_472 = _T_286 | _T_299; // @[Arbiter.scala 98:36:freechips.rocketchip.system.DefaultRV32Config.fir@6065.4]
  assign _T_473 = ~_T_472; // @[Arbiter.scala 98:15:freechips.rocketchip.system.DefaultRV32Config.fir@6066.4]
  assign _T_475 = _T_473 | _T_461; // @[Arbiter.scala 98:41:freechips.rocketchip.system.DefaultRV32Config.fir@6068.4]
  assign _T_477 = _T_475 | reset; // @[Arbiter.scala 98:14:freechips.rocketchip.system.DefaultRV32Config.fir@6070.4]
  assign _T_478 = ~_T_477; // @[Arbiter.scala 98:14:freechips.rocketchip.system.DefaultRV32Config.fir@6071.4]
  assign _T_482 = _T_473 | _T_472; // @[Arbiter.scala 99:41:freechips.rocketchip.system.DefaultRV32Config.fir@6079.4]
  assign _T_484 = _T_482 | reset; // @[Arbiter.scala 99:14:freechips.rocketchip.system.DefaultRV32Config.fir@6081.4]
  assign _T_485 = ~_T_484; // @[Arbiter.scala 99:14:freechips.rocketchip.system.DefaultRV32Config.fir@6082.4]
  assign _T_486 = _T_454 ? _T_216 : 10'h0; // @[Arbiter.scala 102:73:freechips.rocketchip.system.DefaultRV32Config.fir@6087.4]
  assign _T_487 = _T_455 ? _T_224 : 10'h0; // @[Arbiter.scala 102:73:freechips.rocketchip.system.DefaultRV32Config.fir@6088.4]
  assign _T_488 = _T_486 | _T_487; // @[Arbiter.scala 103:44:freechips.rocketchip.system.DefaultRV32Config.fir@6089.4]
  assign _T_497_0 = _T_417 ? _T_454 : _T_496_0; // @[Arbiter.scala 108:30:freechips.rocketchip.system.DefaultRV32Config.fir@6101.4]
  assign _T_497_1 = _T_417 ? _T_455 : _T_496_1; // @[Arbiter.scala 108:30:freechips.rocketchip.system.DefaultRV32Config.fir@6101.4]
  assign _T_503 = _T_496_0 & _T_286; // @[Mux.scala 27:72:freechips.rocketchip.system.DefaultRV32Config.fir@6111.4]
  assign _T_504 = _T_496_1 & _T_299; // @[Mux.scala 27:72:freechips.rocketchip.system.DefaultRV32Config.fir@6112.4]
  assign _T_505 = _T_503 | _T_504; // @[Mux.scala 27:72:freechips.rocketchip.system.DefaultRV32Config.fir@6113.4]
  assign _T_507 = _T_417 ? _T_472 : _T_505; // @[Arbiter.scala 116:29:freechips.rocketchip.system.DefaultRV32Config.fir@6116.4]
  assign _T_491 = auto_out_0_a_ready & _T_507; // @[ReadyValidCancel.scala 52:33:freechips.rocketchip.system.DefaultRV32Config.fir@6092.4]
  assign _GEN_19 = {{9'd0}, _T_491}; // @[Arbiter.scala 104:52:freechips.rocketchip.system.DefaultRV32Config.fir@6093.4]
  assign _T_493 = _T_416 - _GEN_19; // @[Arbiter.scala 104:52:freechips.rocketchip.system.DefaultRV32Config.fir@6094.4]
  assign _T_517 = {auto_in_0_a_bits_user_amba_prot_writealloc,auto_in_0_a_bits_user_amba_prot_privileged,auto_in_0_a_bits_user_amba_prot_secure,auto_in_0_a_bits_user_amba_prot_fetch,auto_in_0_a_bits_mask,auto_in_0_a_bits_data,auto_in_0_a_bits_corrupt}; // @[Mux.scala 27:72:freechips.rocketchip.system.DefaultRV32Config.fir@6129.4]
  assign _T_13_0_a_bits_source = {{1'd0}, auto_in_0_a_bits_source}; // @[Xbar.scala 225:18:freechips.rocketchip.system.DefaultRV32Config.fir@4994.4 BundleMap.scala 248:19:freechips.rocketchip.system.DefaultRV32Config.fir@5006.4 Xbar.scala 231:29:freechips.rocketchip.system.DefaultRV32Config.fir@5014.4]
  assign _T_525 = {auto_in_0_a_bits_opcode,auto_in_0_a_bits_param,auto_in_0_a_bits_size,_T_13_0_a_bits_source,auto_in_0_a_bits_address,auto_in_0_a_bits_user_amba_prot_bufferable,auto_in_0_a_bits_user_amba_prot_modifiable,auto_in_0_a_bits_user_amba_prot_readalloc,_T_517}; // @[Mux.scala 27:72:freechips.rocketchip.system.DefaultRV32Config.fir@6137.4]
  assign _T_526 = _T_497_0 ? _T_525 : 91'h0; // @[Mux.scala 27:72:freechips.rocketchip.system.DefaultRV32Config.fir@6138.4]
  assign _T_532 = {4'h6,auto_in_1_a_bits_mask,auto_in_1_a_bits_data,auto_in_1_a_bits_corrupt}; // @[Mux.scala 27:72:freechips.rocketchip.system.DefaultRV32Config.fir@6144.4]
  assign _T_540 = {auto_in_1_a_bits_opcode,auto_in_1_a_bits_param,auto_in_1_a_bits_size,_T_16,auto_in_1_a_bits_address,1'h0,2'h0,_T_532}; // @[Mux.scala 27:72:freechips.rocketchip.system.DefaultRV32Config.fir@6152.4]
  assign _T_541 = _T_497_1 ? _T_540 : 91'h0; // @[Mux.scala 27:72:freechips.rocketchip.system.DefaultRV32Config.fir@6153.4]
  assign _T_542 = _T_526 | _T_541; // @[Mux.scala 27:72:freechips.rocketchip.system.DefaultRV32Config.fir@6154.4]
  assign _T_570 = _T_569 & auto_out_1_a_ready; // @[Arbiter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@6253.4]
  assign _T_595 = |_T_575; // @[Arbiter.scala 26:27:freechips.rocketchip.system.DefaultRV32Config.fir@6282.4]
  assign _T_596 = _T_570 & _T_595; // @[Arbiter.scala 26:18:freechips.rocketchip.system.DefaultRV32Config.fir@6283.4]
  assign _T_597 = _T_594 & _T_575; // @[Arbiter.scala 27:29:freechips.rocketchip.system.DefaultRV32Config.fir@6285.6]
  assign _T_598 = {_T_597, 1'h0}; // @[package.scala 217:48:freechips.rocketchip.system.DefaultRV32Config.fir@6286.6]
  assign _T_600 = _T_597 | _T_598[1:0]; // @[package.scala 217:43:freechips.rocketchip.system.DefaultRV32Config.fir@6288.6]
  assign _T_606 = _T_594[0] & _T_288; // @[Arbiter.scala 88:79:freechips.rocketchip.system.DefaultRV32Config.fir@6298.4]
  assign _T_607 = _T_594[1] & _T_301; // @[Arbiter.scala 88:79:freechips.rocketchip.system.DefaultRV32Config.fir@6299.4]
  assign _T_613 = _T_606 | _T_607; // @[Arbiter.scala 95:53:freechips.rocketchip.system.DefaultRV32Config.fir@6309.4]
  assign _T_615 = ~_T_606; // @[Arbiter.scala 96:67:freechips.rocketchip.system.DefaultRV32Config.fir@6311.4]
  assign _T_618 = ~_T_607; // @[Arbiter.scala 96:67:freechips.rocketchip.system.DefaultRV32Config.fir@6314.4]
  assign _T_619 = _T_615 | _T_618; // @[Arbiter.scala 96:64:freechips.rocketchip.system.DefaultRV32Config.fir@6315.4]
  assign _T_622 = _T_619 | reset; // @[Arbiter.scala 96:13:freechips.rocketchip.system.DefaultRV32Config.fir@6318.4]
  assign _T_623 = ~_T_622; // @[Arbiter.scala 96:13:freechips.rocketchip.system.DefaultRV32Config.fir@6319.4]
  assign _T_624 = _T_288 | _T_301; // @[Arbiter.scala 98:36:freechips.rocketchip.system.DefaultRV32Config.fir@6324.4]
  assign _T_625 = ~_T_624; // @[Arbiter.scala 98:15:freechips.rocketchip.system.DefaultRV32Config.fir@6325.4]
  assign _T_627 = _T_625 | _T_613; // @[Arbiter.scala 98:41:freechips.rocketchip.system.DefaultRV32Config.fir@6327.4]
  assign _T_629 = _T_627 | reset; // @[Arbiter.scala 98:14:freechips.rocketchip.system.DefaultRV32Config.fir@6329.4]
  assign _T_630 = ~_T_629; // @[Arbiter.scala 98:14:freechips.rocketchip.system.DefaultRV32Config.fir@6330.4]
  assign _T_634 = _T_625 | _T_624; // @[Arbiter.scala 99:41:freechips.rocketchip.system.DefaultRV32Config.fir@6338.4]
  assign _T_636 = _T_634 | reset; // @[Arbiter.scala 99:14:freechips.rocketchip.system.DefaultRV32Config.fir@6340.4]
  assign _T_637 = ~_T_636; // @[Arbiter.scala 99:14:freechips.rocketchip.system.DefaultRV32Config.fir@6341.4]
  assign _T_638 = _T_606 ? _T_216 : 10'h0; // @[Arbiter.scala 102:73:freechips.rocketchip.system.DefaultRV32Config.fir@6346.4]
  assign _T_639 = _T_607 ? _T_224 : 10'h0; // @[Arbiter.scala 102:73:freechips.rocketchip.system.DefaultRV32Config.fir@6347.4]
  assign _T_640 = _T_638 | _T_639; // @[Arbiter.scala 103:44:freechips.rocketchip.system.DefaultRV32Config.fir@6348.4]
  assign _T_649_0 = _T_569 ? _T_606 : _T_648_0; // @[Arbiter.scala 108:30:freechips.rocketchip.system.DefaultRV32Config.fir@6360.4]
  assign _T_649_1 = _T_569 ? _T_607 : _T_648_1; // @[Arbiter.scala 108:30:freechips.rocketchip.system.DefaultRV32Config.fir@6360.4]
  assign _T_655 = _T_648_0 & _T_288; // @[Mux.scala 27:72:freechips.rocketchip.system.DefaultRV32Config.fir@6370.4]
  assign _T_656 = _T_648_1 & _T_301; // @[Mux.scala 27:72:freechips.rocketchip.system.DefaultRV32Config.fir@6371.4]
  assign _T_657 = _T_655 | _T_656; // @[Mux.scala 27:72:freechips.rocketchip.system.DefaultRV32Config.fir@6372.4]
  assign _T_659 = _T_569 ? _T_624 : _T_657; // @[Arbiter.scala 116:29:freechips.rocketchip.system.DefaultRV32Config.fir@6375.4]
  assign _T_643 = auto_out_1_a_ready & _T_659; // @[ReadyValidCancel.scala 52:33:freechips.rocketchip.system.DefaultRV32Config.fir@6351.4]
  assign _GEN_20 = {{9'd0}, _T_643}; // @[Arbiter.scala 104:52:freechips.rocketchip.system.DefaultRV32Config.fir@6352.4]
  assign _T_645 = _T_568 - _GEN_20; // @[Arbiter.scala 104:52:freechips.rocketchip.system.DefaultRV32Config.fir@6353.4]
  assign _T_678 = _T_649_0 ? _T_525 : 91'h0; // @[Mux.scala 27:72:freechips.rocketchip.system.DefaultRV32Config.fir@6397.4]
  assign _T_693 = _T_649_1 ? _T_540 : 91'h0; // @[Mux.scala 27:72:freechips.rocketchip.system.DefaultRV32Config.fir@6412.4]
  assign _T_694 = _T_678 | _T_693; // @[Mux.scala 27:72:freechips.rocketchip.system.DefaultRV32Config.fir@6413.4]
  assign _T_724 = _T_723 & auto_out_2_a_ready; // @[Arbiter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@6528.4]
  assign _T_749 = |_T_729; // @[Arbiter.scala 26:27:freechips.rocketchip.system.DefaultRV32Config.fir@6557.4]
  assign _T_750 = _T_724 & _T_749; // @[Arbiter.scala 26:18:freechips.rocketchip.system.DefaultRV32Config.fir@6558.4]
  assign _T_751 = _T_748 & _T_729; // @[Arbiter.scala 27:29:freechips.rocketchip.system.DefaultRV32Config.fir@6560.6]
  assign _T_752 = {_T_751, 1'h0}; // @[package.scala 217:48:freechips.rocketchip.system.DefaultRV32Config.fir@6561.6]
  assign _T_754 = _T_751 | _T_752[1:0]; // @[package.scala 217:43:freechips.rocketchip.system.DefaultRV32Config.fir@6563.6]
  assign _T_760 = _T_748[0] & _T_290; // @[Arbiter.scala 88:79:freechips.rocketchip.system.DefaultRV32Config.fir@6573.4]
  assign _T_761 = _T_748[1] & _T_303; // @[Arbiter.scala 88:79:freechips.rocketchip.system.DefaultRV32Config.fir@6574.4]
  assign _T_767 = _T_760 | _T_761; // @[Arbiter.scala 95:53:freechips.rocketchip.system.DefaultRV32Config.fir@6584.4]
  assign _T_769 = ~_T_760; // @[Arbiter.scala 96:67:freechips.rocketchip.system.DefaultRV32Config.fir@6586.4]
  assign _T_772 = ~_T_761; // @[Arbiter.scala 96:67:freechips.rocketchip.system.DefaultRV32Config.fir@6589.4]
  assign _T_773 = _T_769 | _T_772; // @[Arbiter.scala 96:64:freechips.rocketchip.system.DefaultRV32Config.fir@6590.4]
  assign _T_776 = _T_773 | reset; // @[Arbiter.scala 96:13:freechips.rocketchip.system.DefaultRV32Config.fir@6593.4]
  assign _T_777 = ~_T_776; // @[Arbiter.scala 96:13:freechips.rocketchip.system.DefaultRV32Config.fir@6594.4]
  assign _T_778 = _T_290 | _T_303; // @[Arbiter.scala 98:36:freechips.rocketchip.system.DefaultRV32Config.fir@6599.4]
  assign _T_779 = ~_T_778; // @[Arbiter.scala 98:15:freechips.rocketchip.system.DefaultRV32Config.fir@6600.4]
  assign _T_781 = _T_779 | _T_767; // @[Arbiter.scala 98:41:freechips.rocketchip.system.DefaultRV32Config.fir@6602.4]
  assign _T_783 = _T_781 | reset; // @[Arbiter.scala 98:14:freechips.rocketchip.system.DefaultRV32Config.fir@6604.4]
  assign _T_784 = ~_T_783; // @[Arbiter.scala 98:14:freechips.rocketchip.system.DefaultRV32Config.fir@6605.4]
  assign _T_788 = _T_779 | _T_778; // @[Arbiter.scala 99:41:freechips.rocketchip.system.DefaultRV32Config.fir@6613.4]
  assign _T_790 = _T_788 | reset; // @[Arbiter.scala 99:14:freechips.rocketchip.system.DefaultRV32Config.fir@6615.4]
  assign _T_791 = ~_T_790; // @[Arbiter.scala 99:14:freechips.rocketchip.system.DefaultRV32Config.fir@6616.4]
  assign _T_792 = _T_760 ? _T_216 : 10'h0; // @[Arbiter.scala 102:73:freechips.rocketchip.system.DefaultRV32Config.fir@6621.4]
  assign _T_793 = _T_761 ? _T_224 : 10'h0; // @[Arbiter.scala 102:73:freechips.rocketchip.system.DefaultRV32Config.fir@6622.4]
  assign _T_794 = _T_792 | _T_793; // @[Arbiter.scala 103:44:freechips.rocketchip.system.DefaultRV32Config.fir@6623.4]
  assign _T_803_0 = _T_723 ? _T_760 : _T_802_0; // @[Arbiter.scala 108:30:freechips.rocketchip.system.DefaultRV32Config.fir@6635.4]
  assign _T_803_1 = _T_723 ? _T_761 : _T_802_1; // @[Arbiter.scala 108:30:freechips.rocketchip.system.DefaultRV32Config.fir@6635.4]
  assign _T_809 = _T_802_0 & _T_290; // @[Mux.scala 27:72:freechips.rocketchip.system.DefaultRV32Config.fir@6645.4]
  assign _T_810 = _T_802_1 & _T_303; // @[Mux.scala 27:72:freechips.rocketchip.system.DefaultRV32Config.fir@6646.4]
  assign _T_811 = _T_809 | _T_810; // @[Mux.scala 27:72:freechips.rocketchip.system.DefaultRV32Config.fir@6647.4]
  assign _T_813 = _T_723 ? _T_778 : _T_811; // @[Arbiter.scala 116:29:freechips.rocketchip.system.DefaultRV32Config.fir@6650.4]
  assign _T_797 = auto_out_2_a_ready & _T_813; // @[ReadyValidCancel.scala 52:33:freechips.rocketchip.system.DefaultRV32Config.fir@6626.4]
  assign _GEN_21 = {{9'd0}, _T_797}; // @[Arbiter.scala 104:52:freechips.rocketchip.system.DefaultRV32Config.fir@6627.4]
  assign _T_799 = _T_722 - _GEN_21; // @[Arbiter.scala 104:52:freechips.rocketchip.system.DefaultRV32Config.fir@6628.4]
  assign _T_832 = _T_803_0 ? _T_525 : 91'h0; // @[Mux.scala 27:72:freechips.rocketchip.system.DefaultRV32Config.fir@6672.4]
  assign _T_847 = _T_803_1 ? _T_540 : 91'h0; // @[Mux.scala 27:72:freechips.rocketchip.system.DefaultRV32Config.fir@6687.4]
  assign _T_848 = _T_832 | _T_847; // @[Mux.scala 27:72:freechips.rocketchip.system.DefaultRV32Config.fir@6688.4]
  assign _T_884 = _T_883 & auto_in_0_d_ready; // @[Arbiter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@6858.4]
  assign _T_914 = |_T_892; // @[Arbiter.scala 26:27:freechips.rocketchip.system.DefaultRV32Config.fir@6892.4]
  assign _T_915 = _T_884 & _T_914; // @[Arbiter.scala 26:18:freechips.rocketchip.system.DefaultRV32Config.fir@6893.4]
  assign _T_916 = _T_913 & _T_892; // @[Arbiter.scala 27:29:freechips.rocketchip.system.DefaultRV32Config.fir@6895.6]
  assign _T_917 = {_T_916, 1'h0}; // @[package.scala 217:48:freechips.rocketchip.system.DefaultRV32Config.fir@6896.6]
  assign _T_919 = _T_916 | _T_917[2:0]; // @[package.scala 217:43:freechips.rocketchip.system.DefaultRV32Config.fir@6898.6]
  assign _T_920 = {_T_919, 2'h0}; // @[package.scala 217:48:freechips.rocketchip.system.DefaultRV32Config.fir@6899.6]
  assign _T_922 = _T_919 | _T_920[2:0]; // @[package.scala 217:43:freechips.rocketchip.system.DefaultRV32Config.fir@6901.6]
  assign _T_938 = _T_929 | _T_930; // @[Arbiter.scala 95:53:freechips.rocketchip.system.DefaultRV32Config.fir@6928.4]
  assign _T_939 = _T_938 | _T_931; // @[Arbiter.scala 95:53:freechips.rocketchip.system.DefaultRV32Config.fir@6929.4]
  assign _T_941 = ~_T_929; // @[Arbiter.scala 96:67:freechips.rocketchip.system.DefaultRV32Config.fir@6931.4]
  assign _T_944 = ~_T_930; // @[Arbiter.scala 96:67:freechips.rocketchip.system.DefaultRV32Config.fir@6934.4]
  assign _T_945 = _T_941 | _T_944; // @[Arbiter.scala 96:64:freechips.rocketchip.system.DefaultRV32Config.fir@6935.4]
  assign _T_946 = ~_T_938; // @[Arbiter.scala 96:61:freechips.rocketchip.system.DefaultRV32Config.fir@6936.4]
  assign _T_947 = ~_T_931; // @[Arbiter.scala 96:67:freechips.rocketchip.system.DefaultRV32Config.fir@6937.4]
  assign _T_948 = _T_946 | _T_947; // @[Arbiter.scala 96:64:freechips.rocketchip.system.DefaultRV32Config.fir@6938.4]
  assign _T_950 = _T_945 & _T_948; // @[Arbiter.scala 96:82:freechips.rocketchip.system.DefaultRV32Config.fir@6940.4]
  assign _T_952 = _T_950 | reset; // @[Arbiter.scala 96:13:freechips.rocketchip.system.DefaultRV32Config.fir@6942.4]
  assign _T_953 = ~_T_952; // @[Arbiter.scala 96:13:freechips.rocketchip.system.DefaultRV32Config.fir@6943.4]
  assign _T_954 = _T_365 | _T_374; // @[Arbiter.scala 98:36:freechips.rocketchip.system.DefaultRV32Config.fir@6948.4]
  assign _T_955 = _T_954 | _T_383; // @[Arbiter.scala 98:36:freechips.rocketchip.system.DefaultRV32Config.fir@6949.4]
  assign _T_956 = ~_T_955; // @[Arbiter.scala 98:15:freechips.rocketchip.system.DefaultRV32Config.fir@6950.4]
  assign _T_959 = _T_956 | _T_939; // @[Arbiter.scala 98:41:freechips.rocketchip.system.DefaultRV32Config.fir@6953.4]
  assign _T_961 = _T_959 | reset; // @[Arbiter.scala 98:14:freechips.rocketchip.system.DefaultRV32Config.fir@6955.4]
  assign _T_962 = ~_T_961; // @[Arbiter.scala 98:14:freechips.rocketchip.system.DefaultRV32Config.fir@6956.4]
  assign _T_968 = _T_956 | _T_955; // @[Arbiter.scala 99:41:freechips.rocketchip.system.DefaultRV32Config.fir@6966.4]
  assign _T_970 = _T_968 | reset; // @[Arbiter.scala 99:14:freechips.rocketchip.system.DefaultRV32Config.fir@6968.4]
  assign _T_971 = ~_T_970; // @[Arbiter.scala 99:14:freechips.rocketchip.system.DefaultRV32Config.fir@6969.4]
  assign _T_972 = _T_929 ? _T_269 : 10'h0; // @[Arbiter.scala 102:73:freechips.rocketchip.system.DefaultRV32Config.fir@6974.4]
  assign _T_973 = _T_930 ? _T_276 : 4'h0; // @[Arbiter.scala 102:73:freechips.rocketchip.system.DefaultRV32Config.fir@6975.4]
  assign _T_974 = _T_931 ? _T_283 : 6'h0; // @[Arbiter.scala 102:73:freechips.rocketchip.system.DefaultRV32Config.fir@6976.4]
  assign _GEN_22 = {{6'd0}, _T_973}; // @[Arbiter.scala 103:44:freechips.rocketchip.system.DefaultRV32Config.fir@6977.4]
  assign _T_975 = _T_972 | _GEN_22; // @[Arbiter.scala 103:44:freechips.rocketchip.system.DefaultRV32Config.fir@6977.4]
  assign _GEN_23 = {{4'd0}, _T_974}; // @[Arbiter.scala 103:44:freechips.rocketchip.system.DefaultRV32Config.fir@6978.4]
  assign _T_976 = _T_975 | _GEN_23; // @[Arbiter.scala 103:44:freechips.rocketchip.system.DefaultRV32Config.fir@6978.4]
  assign _T_993 = _T_984_0 & _T_365; // @[Mux.scala 27:72:freechips.rocketchip.system.DefaultRV32Config.fir@7005.4]
  assign _T_994 = _T_984_1 & _T_374; // @[Mux.scala 27:72:freechips.rocketchip.system.DefaultRV32Config.fir@7006.4]
  assign _T_996 = _T_993 | _T_994; // @[Mux.scala 27:72:freechips.rocketchip.system.DefaultRV32Config.fir@7008.4]
  assign _T_995 = _T_984_2 & _T_383; // @[Mux.scala 27:72:freechips.rocketchip.system.DefaultRV32Config.fir@7007.4]
  assign _T_997 = _T_996 | _T_995; // @[Mux.scala 27:72:freechips.rocketchip.system.DefaultRV32Config.fir@7009.4]
  assign _T_999 = _T_883 ? _T_955 : _T_997; // @[Arbiter.scala 116:29:freechips.rocketchip.system.DefaultRV32Config.fir@7012.4]
  assign _T_979 = auto_in_0_d_ready & _T_999; // @[ReadyValidCancel.scala 52:33:freechips.rocketchip.system.DefaultRV32Config.fir@6981.4]
  assign _GEN_24 = {{9'd0}, _T_979}; // @[Arbiter.scala 104:52:freechips.rocketchip.system.DefaultRV32Config.fir@6982.4]
  assign _T_981 = _T_882 - _GEN_24; // @[Arbiter.scala 104:52:freechips.rocketchip.system.DefaultRV32Config.fir@6983.4]
  assign _T_1056 = _T_1055 & auto_in_1_d_ready; // @[Arbiter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@7187.4]
  assign _T_1086 = |_T_1064; // @[Arbiter.scala 26:27:freechips.rocketchip.system.DefaultRV32Config.fir@7221.4]
  assign _T_1087 = _T_1056 & _T_1086; // @[Arbiter.scala 26:18:freechips.rocketchip.system.DefaultRV32Config.fir@7222.4]
  assign _T_1088 = _T_1085 & _T_1064; // @[Arbiter.scala 27:29:freechips.rocketchip.system.DefaultRV32Config.fir@7224.6]
  assign _T_1089 = {_T_1088, 1'h0}; // @[package.scala 217:48:freechips.rocketchip.system.DefaultRV32Config.fir@7225.6]
  assign _T_1091 = _T_1088 | _T_1089[2:0]; // @[package.scala 217:43:freechips.rocketchip.system.DefaultRV32Config.fir@7227.6]
  assign _T_1092 = {_T_1091, 2'h0}; // @[package.scala 217:48:freechips.rocketchip.system.DefaultRV32Config.fir@7228.6]
  assign _T_1094 = _T_1091 | _T_1092[2:0]; // @[package.scala 217:43:freechips.rocketchip.system.DefaultRV32Config.fir@7230.6]
  assign _T_1110 = _T_1101 | _T_1102; // @[Arbiter.scala 95:53:freechips.rocketchip.system.DefaultRV32Config.fir@7257.4]
  assign _T_1111 = _T_1110 | _T_1103; // @[Arbiter.scala 95:53:freechips.rocketchip.system.DefaultRV32Config.fir@7258.4]
  assign _T_1113 = ~_T_1101; // @[Arbiter.scala 96:67:freechips.rocketchip.system.DefaultRV32Config.fir@7260.4]
  assign _T_1116 = ~_T_1102; // @[Arbiter.scala 96:67:freechips.rocketchip.system.DefaultRV32Config.fir@7263.4]
  assign _T_1117 = _T_1113 | _T_1116; // @[Arbiter.scala 96:64:freechips.rocketchip.system.DefaultRV32Config.fir@7264.4]
  assign _T_1118 = ~_T_1110; // @[Arbiter.scala 96:61:freechips.rocketchip.system.DefaultRV32Config.fir@7265.4]
  assign _T_1119 = ~_T_1103; // @[Arbiter.scala 96:67:freechips.rocketchip.system.DefaultRV32Config.fir@7266.4]
  assign _T_1120 = _T_1118 | _T_1119; // @[Arbiter.scala 96:64:freechips.rocketchip.system.DefaultRV32Config.fir@7267.4]
  assign _T_1122 = _T_1117 & _T_1120; // @[Arbiter.scala 96:82:freechips.rocketchip.system.DefaultRV32Config.fir@7269.4]
  assign _T_1124 = _T_1122 | reset; // @[Arbiter.scala 96:13:freechips.rocketchip.system.DefaultRV32Config.fir@7271.4]
  assign _T_1125 = ~_T_1124; // @[Arbiter.scala 96:13:freechips.rocketchip.system.DefaultRV32Config.fir@7272.4]
  assign _T_1126 = _T_367 | _T_376; // @[Arbiter.scala 98:36:freechips.rocketchip.system.DefaultRV32Config.fir@7277.4]
  assign _T_1127 = _T_1126 | _T_385; // @[Arbiter.scala 98:36:freechips.rocketchip.system.DefaultRV32Config.fir@7278.4]
  assign _T_1128 = ~_T_1127; // @[Arbiter.scala 98:15:freechips.rocketchip.system.DefaultRV32Config.fir@7279.4]
  assign _T_1131 = _T_1128 | _T_1111; // @[Arbiter.scala 98:41:freechips.rocketchip.system.DefaultRV32Config.fir@7282.4]
  assign _T_1133 = _T_1131 | reset; // @[Arbiter.scala 98:14:freechips.rocketchip.system.DefaultRV32Config.fir@7284.4]
  assign _T_1134 = ~_T_1133; // @[Arbiter.scala 98:14:freechips.rocketchip.system.DefaultRV32Config.fir@7285.4]
  assign _T_1140 = _T_1128 | _T_1127; // @[Arbiter.scala 99:41:freechips.rocketchip.system.DefaultRV32Config.fir@7295.4]
  assign _T_1142 = _T_1140 | reset; // @[Arbiter.scala 99:14:freechips.rocketchip.system.DefaultRV32Config.fir@7297.4]
  assign _T_1143 = ~_T_1142; // @[Arbiter.scala 99:14:freechips.rocketchip.system.DefaultRV32Config.fir@7298.4]
  assign _T_1144 = _T_1101 ? _T_269 : 10'h0; // @[Arbiter.scala 102:73:freechips.rocketchip.system.DefaultRV32Config.fir@7303.4]
  assign _T_1145 = _T_1102 ? _T_276 : 4'h0; // @[Arbiter.scala 102:73:freechips.rocketchip.system.DefaultRV32Config.fir@7304.4]
  assign _T_1146 = _T_1103 ? _T_283 : 6'h0; // @[Arbiter.scala 102:73:freechips.rocketchip.system.DefaultRV32Config.fir@7305.4]
  assign _GEN_25 = {{6'd0}, _T_1145}; // @[Arbiter.scala 103:44:freechips.rocketchip.system.DefaultRV32Config.fir@7306.4]
  assign _T_1147 = _T_1144 | _GEN_25; // @[Arbiter.scala 103:44:freechips.rocketchip.system.DefaultRV32Config.fir@7306.4]
  assign _GEN_26 = {{4'd0}, _T_1146}; // @[Arbiter.scala 103:44:freechips.rocketchip.system.DefaultRV32Config.fir@7307.4]
  assign _T_1148 = _T_1147 | _GEN_26; // @[Arbiter.scala 103:44:freechips.rocketchip.system.DefaultRV32Config.fir@7307.4]
  assign _T_1165 = _T_1156_0 & _T_367; // @[Mux.scala 27:72:freechips.rocketchip.system.DefaultRV32Config.fir@7334.4]
  assign _T_1166 = _T_1156_1 & _T_376; // @[Mux.scala 27:72:freechips.rocketchip.system.DefaultRV32Config.fir@7335.4]
  assign _T_1168 = _T_1165 | _T_1166; // @[Mux.scala 27:72:freechips.rocketchip.system.DefaultRV32Config.fir@7337.4]
  assign _T_1167 = _T_1156_2 & _T_385; // @[Mux.scala 27:72:freechips.rocketchip.system.DefaultRV32Config.fir@7336.4]
  assign _T_1169 = _T_1168 | _T_1167; // @[Mux.scala 27:72:freechips.rocketchip.system.DefaultRV32Config.fir@7338.4]
  assign _T_1171 = _T_1055 ? _T_1127 : _T_1169; // @[Arbiter.scala 116:29:freechips.rocketchip.system.DefaultRV32Config.fir@7341.4]
  assign _T_1151 = auto_in_1_d_ready & _T_1171; // @[ReadyValidCancel.scala 52:33:freechips.rocketchip.system.DefaultRV32Config.fir@7310.4]
  assign _GEN_27 = {{9'd0}, _T_1151}; // @[Arbiter.scala 104:52:freechips.rocketchip.system.DefaultRV32Config.fir@7311.4]
  assign _T_1153 = _T_1054 - _GEN_27; // @[Arbiter.scala 104:52:freechips.rocketchip.system.DefaultRV32Config.fir@7312.4]
  assign auto_in_1_a_ready = _T_307 | _T_306; // @[LazyModule.scala 303:16:freechips.rocketchip.system.DefaultRV32Config.fir@4889.4]
  assign auto_in_1_b_valid = auto_out_1_b_valid; // @[LazyModule.scala 303:16:freechips.rocketchip.system.DefaultRV32Config.fir@4889.4]
  assign auto_in_1_b_bits_param = auto_out_1_b_bits_param; // @[LazyModule.scala 303:16:freechips.rocketchip.system.DefaultRV32Config.fir@4889.4]
  assign auto_in_1_b_bits_address = auto_out_1_b_bits_address; // @[LazyModule.scala 303:16:freechips.rocketchip.system.DefaultRV32Config.fir@4889.4]
  assign auto_in_1_c_ready = auto_out_1_c_ready; // @[LazyModule.scala 303:16:freechips.rocketchip.system.DefaultRV32Config.fir@4889.4]
  assign auto_in_1_d_valid = _T_1055 ? _T_1127 : _T_1169; // @[LazyModule.scala 303:16:freechips.rocketchip.system.DefaultRV32Config.fir@4889.4]
  assign auto_in_1_d_bits_opcode = _T_1203[49:47]; // @[LazyModule.scala 303:16:freechips.rocketchip.system.DefaultRV32Config.fir@4889.4]
  assign auto_in_1_d_bits_param = _T_1203[46:45]; // @[LazyModule.scala 303:16:freechips.rocketchip.system.DefaultRV32Config.fir@4889.4]
  assign auto_in_1_d_bits_size = _T_1203[44:41]; // @[LazyModule.scala 303:16:freechips.rocketchip.system.DefaultRV32Config.fir@4889.4]
  assign auto_in_1_d_bits_source = _T_1203[37:36]; // @[LazyModule.scala 303:16:freechips.rocketchip.system.DefaultRV32Config.fir@4889.4]
  assign auto_in_1_d_bits_sink = _T_1203[35:34]; // @[LazyModule.scala 303:16:freechips.rocketchip.system.DefaultRV32Config.fir@4889.4]
  assign auto_in_1_d_bits_denied = _T_1203[33]; // @[LazyModule.scala 303:16:freechips.rocketchip.system.DefaultRV32Config.fir@4889.4]
  assign auto_in_1_d_bits_data = _T_1203[32:1]; // @[LazyModule.scala 303:16:freechips.rocketchip.system.DefaultRV32Config.fir@4889.4]
  assign auto_in_1_d_bits_corrupt = _T_1203[0]; // @[LazyModule.scala 303:16:freechips.rocketchip.system.DefaultRV32Config.fir@4889.4]
  assign auto_in_0_a_ready = _T_294 | _T_293; // @[LazyModule.scala 303:16:freechips.rocketchip.system.DefaultRV32Config.fir@4888.4]
  assign auto_in_0_d_valid = _T_883 ? _T_955 : _T_997; // @[LazyModule.scala 303:16:freechips.rocketchip.system.DefaultRV32Config.fir@4888.4]
  assign auto_in_0_d_bits_opcode = _T_1031[49:47]; // @[LazyModule.scala 303:16:freechips.rocketchip.system.DefaultRV32Config.fir@4888.4]
  assign auto_in_0_d_bits_param = _T_1031[46:45]; // @[LazyModule.scala 303:16:freechips.rocketchip.system.DefaultRV32Config.fir@4888.4]
  assign auto_in_0_d_bits_size = _T_1031[44:41]; // @[LazyModule.scala 303:16:freechips.rocketchip.system.DefaultRV32Config.fir@4888.4]
  assign auto_in_0_d_bits_source = _T_1031[39:36]; // @[LazyModule.scala 303:16:freechips.rocketchip.system.DefaultRV32Config.fir@4888.4]
  assign auto_in_0_d_bits_sink = _T_1031[35:34]; // @[LazyModule.scala 303:16:freechips.rocketchip.system.DefaultRV32Config.fir@4888.4]
  assign auto_in_0_d_bits_denied = _T_1031[33]; // @[LazyModule.scala 303:16:freechips.rocketchip.system.DefaultRV32Config.fir@4888.4]
  assign auto_in_0_d_bits_data = _T_1031[32:1]; // @[LazyModule.scala 303:16:freechips.rocketchip.system.DefaultRV32Config.fir@4888.4]
  assign auto_in_0_d_bits_corrupt = _T_1031[0]; // @[LazyModule.scala 303:16:freechips.rocketchip.system.DefaultRV32Config.fir@4888.4]
  assign auto_out_2_a_valid = _T_723 ? _T_778 : _T_811; // @[LazyModule.scala 305:12:freechips.rocketchip.system.DefaultRV32Config.fir@4887.4]
  assign auto_out_2_a_bits_opcode = _T_848[90:88]; // @[LazyModule.scala 305:12:freechips.rocketchip.system.DefaultRV32Config.fir@4887.4]
  assign auto_out_2_a_bits_param = _T_848[87:85]; // @[LazyModule.scala 305:12:freechips.rocketchip.system.DefaultRV32Config.fir@4887.4]
  assign auto_out_2_a_bits_size = _T_848[84:81]; // @[LazyModule.scala 305:12:freechips.rocketchip.system.DefaultRV32Config.fir@4887.4]
  assign auto_out_2_a_bits_source = _T_848[80:76]; // @[LazyModule.scala 305:12:freechips.rocketchip.system.DefaultRV32Config.fir@4887.4]
  assign auto_out_2_a_bits_address = _T_848[74:44]; // @[LazyModule.scala 305:12:freechips.rocketchip.system.DefaultRV32Config.fir@4887.4]
  assign auto_out_2_a_bits_user_amba_prot_bufferable = _T_848[43]; // @[LazyModule.scala 305:12:freechips.rocketchip.system.DefaultRV32Config.fir@4887.4]
  assign auto_out_2_a_bits_user_amba_prot_modifiable = _T_848[42]; // @[LazyModule.scala 305:12:freechips.rocketchip.system.DefaultRV32Config.fir@4887.4]
  assign auto_out_2_a_bits_user_amba_prot_readalloc = _T_848[41]; // @[LazyModule.scala 305:12:freechips.rocketchip.system.DefaultRV32Config.fir@4887.4]
  assign auto_out_2_a_bits_user_amba_prot_writealloc = _T_848[40]; // @[LazyModule.scala 305:12:freechips.rocketchip.system.DefaultRV32Config.fir@4887.4]
  assign auto_out_2_a_bits_user_amba_prot_privileged = _T_848[39]; // @[LazyModule.scala 305:12:freechips.rocketchip.system.DefaultRV32Config.fir@4887.4]
  assign auto_out_2_a_bits_user_amba_prot_secure = _T_848[38]; // @[LazyModule.scala 305:12:freechips.rocketchip.system.DefaultRV32Config.fir@4887.4]
  assign auto_out_2_a_bits_user_amba_prot_fetch = _T_848[37]; // @[LazyModule.scala 305:12:freechips.rocketchip.system.DefaultRV32Config.fir@4887.4]
  assign auto_out_2_a_bits_mask = _T_848[36:33]; // @[LazyModule.scala 305:12:freechips.rocketchip.system.DefaultRV32Config.fir@4887.4]
  assign auto_out_2_a_bits_data = _T_848[32:1]; // @[LazyModule.scala 305:12:freechips.rocketchip.system.DefaultRV32Config.fir@4887.4]
  assign auto_out_2_a_bits_corrupt = _T_848[0]; // @[LazyModule.scala 305:12:freechips.rocketchip.system.DefaultRV32Config.fir@4887.4]
  assign auto_out_2_d_ready = _T_386 | _T_387; // @[LazyModule.scala 305:12:freechips.rocketchip.system.DefaultRV32Config.fir@4887.4]
  assign auto_out_1_a_valid = _T_569 ? _T_624 : _T_657; // @[LazyModule.scala 305:12:freechips.rocketchip.system.DefaultRV32Config.fir@4886.4]
  assign auto_out_1_a_bits_opcode = _T_694[90:88]; // @[LazyModule.scala 305:12:freechips.rocketchip.system.DefaultRV32Config.fir@4886.4]
  assign auto_out_1_a_bits_param = _T_694[87:85]; // @[LazyModule.scala 305:12:freechips.rocketchip.system.DefaultRV32Config.fir@4886.4]
  assign auto_out_1_a_bits_size = _T_694[83:81]; // @[LazyModule.scala 305:12:freechips.rocketchip.system.DefaultRV32Config.fir@4886.4]
  assign auto_out_1_a_bits_source = _T_694[80:76]; // @[LazyModule.scala 305:12:freechips.rocketchip.system.DefaultRV32Config.fir@4886.4]
  assign auto_out_1_a_bits_address = _T_694[75:44]; // @[LazyModule.scala 305:12:freechips.rocketchip.system.DefaultRV32Config.fir@4886.4]
  assign auto_out_1_a_bits_user_amba_prot_bufferable = _T_694[43]; // @[LazyModule.scala 305:12:freechips.rocketchip.system.DefaultRV32Config.fir@4886.4]
  assign auto_out_1_a_bits_user_amba_prot_modifiable = _T_694[42]; // @[LazyModule.scala 305:12:freechips.rocketchip.system.DefaultRV32Config.fir@4886.4]
  assign auto_out_1_a_bits_user_amba_prot_readalloc = _T_694[41]; // @[LazyModule.scala 305:12:freechips.rocketchip.system.DefaultRV32Config.fir@4886.4]
  assign auto_out_1_a_bits_user_amba_prot_writealloc = _T_694[40]; // @[LazyModule.scala 305:12:freechips.rocketchip.system.DefaultRV32Config.fir@4886.4]
  assign auto_out_1_a_bits_user_amba_prot_privileged = _T_694[39]; // @[LazyModule.scala 305:12:freechips.rocketchip.system.DefaultRV32Config.fir@4886.4]
  assign auto_out_1_a_bits_user_amba_prot_secure = _T_694[38]; // @[LazyModule.scala 305:12:freechips.rocketchip.system.DefaultRV32Config.fir@4886.4]
  assign auto_out_1_a_bits_user_amba_prot_fetch = _T_694[37]; // @[LazyModule.scala 305:12:freechips.rocketchip.system.DefaultRV32Config.fir@4886.4]
  assign auto_out_1_a_bits_mask = _T_694[36:33]; // @[LazyModule.scala 305:12:freechips.rocketchip.system.DefaultRV32Config.fir@4886.4]
  assign auto_out_1_a_bits_data = _T_694[32:1]; // @[LazyModule.scala 305:12:freechips.rocketchip.system.DefaultRV32Config.fir@4886.4]
  assign auto_out_1_a_bits_corrupt = _T_694[0]; // @[LazyModule.scala 305:12:freechips.rocketchip.system.DefaultRV32Config.fir@4886.4]
  assign auto_out_1_b_ready = auto_in_1_b_ready; // @[LazyModule.scala 305:12:freechips.rocketchip.system.DefaultRV32Config.fir@4886.4]
  assign auto_out_1_c_valid = auto_in_1_c_valid; // @[LazyModule.scala 305:12:freechips.rocketchip.system.DefaultRV32Config.fir@4886.4]
  assign auto_out_1_c_bits_opcode = auto_in_1_c_bits_opcode; // @[LazyModule.scala 305:12:freechips.rocketchip.system.DefaultRV32Config.fir@4886.4]
  assign auto_out_1_c_bits_param = auto_in_1_c_bits_param; // @[LazyModule.scala 305:12:freechips.rocketchip.system.DefaultRV32Config.fir@4886.4]
  assign auto_out_1_c_bits_size = auto_in_1_c_bits_size[2:0]; // @[LazyModule.scala 305:12:freechips.rocketchip.system.DefaultRV32Config.fir@4886.4]
  assign auto_out_1_c_bits_source = _GEN_9 | 5'h10; // @[LazyModule.scala 305:12:freechips.rocketchip.system.DefaultRV32Config.fir@4886.4]
  assign auto_out_1_c_bits_address = auto_in_1_c_bits_address; // @[LazyModule.scala 305:12:freechips.rocketchip.system.DefaultRV32Config.fir@4886.4]
  assign auto_out_1_c_bits_data = auto_in_1_c_bits_data; // @[LazyModule.scala 305:12:freechips.rocketchip.system.DefaultRV32Config.fir@4886.4]
  assign auto_out_1_c_bits_corrupt = auto_in_1_c_bits_corrupt; // @[LazyModule.scala 305:12:freechips.rocketchip.system.DefaultRV32Config.fir@4886.4]
  assign auto_out_1_d_ready = _T_377 | _T_378; // @[LazyModule.scala 305:12:freechips.rocketchip.system.DefaultRV32Config.fir@4886.4]
  assign auto_out_1_e_valid = auto_in_1_e_valid; // @[LazyModule.scala 305:12:freechips.rocketchip.system.DefaultRV32Config.fir@4886.4]
  assign auto_out_1_e_bits_sink = auto_in_1_e_bits_sink; // @[LazyModule.scala 305:12:freechips.rocketchip.system.DefaultRV32Config.fir@4886.4]
  assign auto_out_0_a_valid = _T_417 ? _T_472 : _T_505; // @[LazyModule.scala 305:12:freechips.rocketchip.system.DefaultRV32Config.fir@4885.4]
  assign auto_out_0_a_bits_opcode = _T_542[90:88]; // @[LazyModule.scala 305:12:freechips.rocketchip.system.DefaultRV32Config.fir@4885.4]
  assign auto_out_0_a_bits_param = _T_542[87:85]; // @[LazyModule.scala 305:12:freechips.rocketchip.system.DefaultRV32Config.fir@4885.4]
  assign auto_out_0_a_bits_size = _T_542[84:81]; // @[LazyModule.scala 305:12:freechips.rocketchip.system.DefaultRV32Config.fir@4885.4]
  assign auto_out_0_a_bits_source = _T_542[80:76]; // @[LazyModule.scala 305:12:freechips.rocketchip.system.DefaultRV32Config.fir@4885.4]
  assign auto_out_0_a_bits_address = _T_542[71:44]; // @[LazyModule.scala 305:12:freechips.rocketchip.system.DefaultRV32Config.fir@4885.4]
  assign auto_out_0_a_bits_mask = _T_542[36:33]; // @[LazyModule.scala 305:12:freechips.rocketchip.system.DefaultRV32Config.fir@4885.4]
  assign auto_out_0_a_bits_data = _T_542[32:1]; // @[LazyModule.scala 305:12:freechips.rocketchip.system.DefaultRV32Config.fir@4885.4]
  assign auto_out_0_a_bits_corrupt = _T_542[0]; // @[LazyModule.scala 305:12:freechips.rocketchip.system.DefaultRV32Config.fir@4885.4]
  assign auto_out_0_d_ready = _T_368 | _T_369; // @[LazyModule.scala 305:12:freechips.rocketchip.system.DefaultRV32Config.fir@4885.4]
  assign TLMonitor_clock = clock; // @[:freechips.rocketchip.system.DefaultRV32Config.fir@4805.4]
  assign TLMonitor_reset = reset; // @[:freechips.rocketchip.system.DefaultRV32Config.fir@4806.4]
  assign TLMonitor_io_in_a_ready = _T_294 | _T_293; // @[Nodes.scala 26:19:freechips.rocketchip.system.DefaultRV32Config.fir@4833.4]
  assign TLMonitor_io_in_a_valid = auto_in_0_a_valid; // @[Nodes.scala 26:19:freechips.rocketchip.system.DefaultRV32Config.fir@4832.4]
  assign TLMonitor_io_in_a_bits_opcode = auto_in_0_a_bits_opcode; // @[Nodes.scala 26:19:freechips.rocketchip.system.DefaultRV32Config.fir@4831.4]
  assign TLMonitor_io_in_a_bits_param = auto_in_0_a_bits_param; // @[Nodes.scala 26:19:freechips.rocketchip.system.DefaultRV32Config.fir@4830.4]
  assign TLMonitor_io_in_a_bits_size = auto_in_0_a_bits_size; // @[Nodes.scala 26:19:freechips.rocketchip.system.DefaultRV32Config.fir@4829.4]
  assign TLMonitor_io_in_a_bits_source = auto_in_0_a_bits_source; // @[Nodes.scala 26:19:freechips.rocketchip.system.DefaultRV32Config.fir@4828.4]
  assign TLMonitor_io_in_a_bits_address = auto_in_0_a_bits_address; // @[Nodes.scala 26:19:freechips.rocketchip.system.DefaultRV32Config.fir@4827.4]
  assign TLMonitor_io_in_a_bits_mask = auto_in_0_a_bits_mask; // @[Nodes.scala 26:19:freechips.rocketchip.system.DefaultRV32Config.fir@4819.4]
  assign TLMonitor_io_in_a_bits_corrupt = auto_in_0_a_bits_corrupt; // @[Nodes.scala 26:19:freechips.rocketchip.system.DefaultRV32Config.fir@4817.4]
  assign TLMonitor_io_in_d_ready = auto_in_0_d_ready; // @[Nodes.scala 26:19:freechips.rocketchip.system.DefaultRV32Config.fir@4816.4]
  assign TLMonitor_io_in_d_valid = _T_883 ? _T_955 : _T_997; // @[Nodes.scala 26:19:freechips.rocketchip.system.DefaultRV32Config.fir@4815.4]
  assign TLMonitor_io_in_d_bits_opcode = _T_1031[49:47]; // @[Nodes.scala 26:19:freechips.rocketchip.system.DefaultRV32Config.fir@4814.4]
  assign TLMonitor_io_in_d_bits_param = _T_1031[46:45]; // @[Nodes.scala 26:19:freechips.rocketchip.system.DefaultRV32Config.fir@4813.4]
  assign TLMonitor_io_in_d_bits_size = _T_1031[44:41]; // @[Nodes.scala 26:19:freechips.rocketchip.system.DefaultRV32Config.fir@4812.4]
  assign TLMonitor_io_in_d_bits_source = _T_1031[39:36]; // @[Nodes.scala 26:19:freechips.rocketchip.system.DefaultRV32Config.fir@4811.4]
  assign TLMonitor_io_in_d_bits_sink = _T_1031[35:34]; // @[Nodes.scala 26:19:freechips.rocketchip.system.DefaultRV32Config.fir@4810.4]
  assign TLMonitor_io_in_d_bits_denied = _T_1031[33]; // @[Nodes.scala 26:19:freechips.rocketchip.system.DefaultRV32Config.fir@4809.4]
  assign TLMonitor_io_in_d_bits_corrupt = _T_1031[0]; // @[Nodes.scala 26:19:freechips.rocketchip.system.DefaultRV32Config.fir@4807.4]
  assign TLMonitor_1_clock = clock; // @[:freechips.rocketchip.system.DefaultRV32Config.fir@4835.4]
  assign TLMonitor_1_reset = reset; // @[:freechips.rocketchip.system.DefaultRV32Config.fir@4836.4]
  assign TLMonitor_1_io_in_a_ready = _T_307 | _T_306; // @[Nodes.scala 26:19:freechips.rocketchip.system.DefaultRV32Config.fir@4878.4]
  assign TLMonitor_1_io_in_a_valid = auto_in_1_a_valid; // @[Nodes.scala 26:19:freechips.rocketchip.system.DefaultRV32Config.fir@4877.4]
  assign TLMonitor_1_io_in_a_bits_opcode = auto_in_1_a_bits_opcode; // @[Nodes.scala 26:19:freechips.rocketchip.system.DefaultRV32Config.fir@4876.4]
  assign TLMonitor_1_io_in_a_bits_param = auto_in_1_a_bits_param; // @[Nodes.scala 26:19:freechips.rocketchip.system.DefaultRV32Config.fir@4875.4]
  assign TLMonitor_1_io_in_a_bits_size = auto_in_1_a_bits_size; // @[Nodes.scala 26:19:freechips.rocketchip.system.DefaultRV32Config.fir@4874.4]
  assign TLMonitor_1_io_in_a_bits_source = auto_in_1_a_bits_source; // @[Nodes.scala 26:19:freechips.rocketchip.system.DefaultRV32Config.fir@4873.4]
  assign TLMonitor_1_io_in_a_bits_address = auto_in_1_a_bits_address; // @[Nodes.scala 26:19:freechips.rocketchip.system.DefaultRV32Config.fir@4872.4]
  assign TLMonitor_1_io_in_a_bits_mask = auto_in_1_a_bits_mask; // @[Nodes.scala 26:19:freechips.rocketchip.system.DefaultRV32Config.fir@4871.4]
  assign TLMonitor_1_io_in_a_bits_corrupt = auto_in_1_a_bits_corrupt; // @[Nodes.scala 26:19:freechips.rocketchip.system.DefaultRV32Config.fir@4869.4]
  assign TLMonitor_1_io_in_b_ready = auto_in_1_b_ready; // @[Nodes.scala 26:19:freechips.rocketchip.system.DefaultRV32Config.fir@4868.4]
  assign TLMonitor_1_io_in_b_valid = auto_out_1_b_valid; // @[Nodes.scala 26:19:freechips.rocketchip.system.DefaultRV32Config.fir@4867.4]
  assign TLMonitor_1_io_in_b_bits_param = auto_out_1_b_bits_param; // @[Nodes.scala 26:19:freechips.rocketchip.system.DefaultRV32Config.fir@4865.4]
  assign TLMonitor_1_io_in_b_bits_address = auto_out_1_b_bits_address; // @[Nodes.scala 26:19:freechips.rocketchip.system.DefaultRV32Config.fir@4862.4]
  assign TLMonitor_1_io_in_c_ready = auto_out_1_c_ready; // @[Nodes.scala 26:19:freechips.rocketchip.system.DefaultRV32Config.fir@4858.4]
  assign TLMonitor_1_io_in_c_valid = auto_in_1_c_valid; // @[Nodes.scala 26:19:freechips.rocketchip.system.DefaultRV32Config.fir@4857.4]
  assign TLMonitor_1_io_in_c_bits_opcode = auto_in_1_c_bits_opcode; // @[Nodes.scala 26:19:freechips.rocketchip.system.DefaultRV32Config.fir@4856.4]
  assign TLMonitor_1_io_in_c_bits_param = auto_in_1_c_bits_param; // @[Nodes.scala 26:19:freechips.rocketchip.system.DefaultRV32Config.fir@4855.4]
  assign TLMonitor_1_io_in_c_bits_size = auto_in_1_c_bits_size; // @[Nodes.scala 26:19:freechips.rocketchip.system.DefaultRV32Config.fir@4854.4]
  assign TLMonitor_1_io_in_c_bits_source = auto_in_1_c_bits_source; // @[Nodes.scala 26:19:freechips.rocketchip.system.DefaultRV32Config.fir@4853.4]
  assign TLMonitor_1_io_in_c_bits_address = auto_in_1_c_bits_address; // @[Nodes.scala 26:19:freechips.rocketchip.system.DefaultRV32Config.fir@4852.4]
  assign TLMonitor_1_io_in_c_bits_corrupt = auto_in_1_c_bits_corrupt; // @[Nodes.scala 26:19:freechips.rocketchip.system.DefaultRV32Config.fir@4850.4]
  assign TLMonitor_1_io_in_d_ready = auto_in_1_d_ready; // @[Nodes.scala 26:19:freechips.rocketchip.system.DefaultRV32Config.fir@4849.4]
  assign TLMonitor_1_io_in_d_valid = _T_1055 ? _T_1127 : _T_1169; // @[Nodes.scala 26:19:freechips.rocketchip.system.DefaultRV32Config.fir@4848.4]
  assign TLMonitor_1_io_in_d_bits_opcode = _T_1203[49:47]; // @[Nodes.scala 26:19:freechips.rocketchip.system.DefaultRV32Config.fir@4847.4]
  assign TLMonitor_1_io_in_d_bits_param = _T_1203[46:45]; // @[Nodes.scala 26:19:freechips.rocketchip.system.DefaultRV32Config.fir@4846.4]
  assign TLMonitor_1_io_in_d_bits_size = _T_1203[44:41]; // @[Nodes.scala 26:19:freechips.rocketchip.system.DefaultRV32Config.fir@4845.4]
  assign TLMonitor_1_io_in_d_bits_source = _T_1203[37:36]; // @[Nodes.scala 26:19:freechips.rocketchip.system.DefaultRV32Config.fir@4844.4]
  assign TLMonitor_1_io_in_d_bits_sink = _T_1203[35:34]; // @[Nodes.scala 26:19:freechips.rocketchip.system.DefaultRV32Config.fir@4843.4]
  assign TLMonitor_1_io_in_d_bits_denied = _T_1203[33]; // @[Nodes.scala 26:19:freechips.rocketchip.system.DefaultRV32Config.fir@4842.4]
  assign TLMonitor_1_io_in_d_bits_corrupt = _T_1203[0]; // @[Nodes.scala 26:19:freechips.rocketchip.system.DefaultRV32Config.fir@4840.4]
  assign TLMonitor_1_io_in_e_valid = auto_in_1_e_valid; // @[Nodes.scala 26:19:freechips.rocketchip.system.DefaultRV32Config.fir@4838.4]
  assign TLMonitor_1_io_in_e_bits_sink = auto_in_1_e_bits_sink; // @[Nodes.scala 26:19:freechips.rocketchip.system.DefaultRV32Config.fir@4837.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_882 = _RAND_0[9:0];
  _RAND_1 = {1{`RANDOM}};
  _T_898 = _RAND_1[2:0];
  _RAND_2 = {1{`RANDOM}};
  _T_984_0 = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  _T_984_1 = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  _T_984_2 = _RAND_4[0:0];
  _RAND_5 = {1{`RANDOM}};
  _T_1054 = _RAND_5[9:0];
  _RAND_6 = {1{`RANDOM}};
  _T_1070 = _RAND_6[2:0];
  _RAND_7 = {1{`RANDOM}};
  _T_1156_0 = _RAND_7[0:0];
  _RAND_8 = {1{`RANDOM}};
  _T_1156_1 = _RAND_8[0:0];
  _RAND_9 = {1{`RANDOM}};
  _T_1156_2 = _RAND_9[0:0];
  _RAND_10 = {1{`RANDOM}};
  _T_416 = _RAND_10[9:0];
  _RAND_11 = {1{`RANDOM}};
  _T_429 = _RAND_11[1:0];
  _RAND_12 = {1{`RANDOM}};
  _T_496_0 = _RAND_12[0:0];
  _RAND_13 = {1{`RANDOM}};
  _T_568 = _RAND_13[9:0];
  _RAND_14 = {1{`RANDOM}};
  _T_581 = _RAND_14[1:0];
  _RAND_15 = {1{`RANDOM}};
  _T_648_0 = _RAND_15[0:0];
  _RAND_16 = {1{`RANDOM}};
  _T_722 = _RAND_16[9:0];
  _RAND_17 = {1{`RANDOM}};
  _T_735 = _RAND_17[1:0];
  _RAND_18 = {1{`RANDOM}};
  _T_802_0 = _RAND_18[0:0];
  _RAND_19 = {1{`RANDOM}};
  _T_496_1 = _RAND_19[0:0];
  _RAND_20 = {1{`RANDOM}};
  _T_648_1 = _RAND_20[0:0];
  _RAND_21 = {1{`RANDOM}};
  _T_802_1 = _RAND_21[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      _T_882 <= 10'h0;
    end else if (_T_884) begin
      _T_882 <= _T_976;
    end else begin
      _T_882 <= _T_981;
    end
    if (reset) begin
      _T_898 <= 3'h7;
    end else if (_T_915) begin
      _T_898 <= _T_922;
    end
    if (reset) begin
      _T_984_0 <= 1'h0;
    end else if (_T_883) begin
      _T_984_0 <= _T_929;
    end
    if (reset) begin
      _T_984_1 <= 1'h0;
    end else if (_T_883) begin
      _T_984_1 <= _T_930;
    end
    if (reset) begin
      _T_984_2 <= 1'h0;
    end else if (_T_883) begin
      _T_984_2 <= _T_931;
    end
    if (reset) begin
      _T_1054 <= 10'h0;
    end else if (_T_1056) begin
      _T_1054 <= _T_1148;
    end else begin
      _T_1054 <= _T_1153;
    end
    if (reset) begin
      _T_1070 <= 3'h7;
    end else if (_T_1087) begin
      _T_1070 <= _T_1094;
    end
    if (reset) begin
      _T_1156_0 <= 1'h0;
    end else if (_T_1055) begin
      _T_1156_0 <= _T_1101;
    end
    if (reset) begin
      _T_1156_1 <= 1'h0;
    end else if (_T_1055) begin
      _T_1156_1 <= _T_1102;
    end
    if (reset) begin
      _T_1156_2 <= 1'h0;
    end else if (_T_1055) begin
      _T_1156_2 <= _T_1103;
    end
    if (reset) begin
      _T_416 <= 10'h0;
    end else if (_T_418) begin
      _T_416 <= _T_488;
    end else begin
      _T_416 <= _T_493;
    end
    if (reset) begin
      _T_429 <= 2'h3;
    end else if (_T_444) begin
      _T_429 <= _T_448;
    end
    if (reset) begin
      _T_496_0 <= 1'h0;
    end else if (_T_417) begin
      _T_496_0 <= _T_454;
    end
    if (reset) begin
      _T_568 <= 10'h0;
    end else if (_T_570) begin
      _T_568 <= _T_640;
    end else begin
      _T_568 <= _T_645;
    end
    if (reset) begin
      _T_581 <= 2'h3;
    end else if (_T_596) begin
      _T_581 <= _T_600;
    end
    if (reset) begin
      _T_648_0 <= 1'h0;
    end else if (_T_569) begin
      _T_648_0 <= _T_606;
    end
    if (reset) begin
      _T_722 <= 10'h0;
    end else if (_T_724) begin
      _T_722 <= _T_794;
    end else begin
      _T_722 <= _T_799;
    end
    if (reset) begin
      _T_735 <= 2'h3;
    end else if (_T_750) begin
      _T_735 <= _T_754;
    end
    if (reset) begin
      _T_802_0 <= 1'h0;
    end else if (_T_723) begin
      _T_802_0 <= _T_760;
    end
    if (reset) begin
      _T_496_1 <= 1'h0;
    end else if (_T_417) begin
      _T_496_1 <= _T_455;
    end
    if (reset) begin
      _T_648_1 <= 1'h0;
    end else if (_T_569) begin
      _T_648_1 <= _T_607;
    end
    if (reset) begin
      _T_802_1 <= 1'h0;
    end else if (_T_723) begin
      _T_802_1 <= _T_761;
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_471) begin
          $fwrite(32'h80000002,"Assertion failed\n    at Arbiter.scala:96 assert((prefixOR zip earlyWinner) map { case (p,w) => !p || !w } reduce {_ && _})\n"); // @[Arbiter.scala 96:13:freechips.rocketchip.system.DefaultRV32Config.fir@6062.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_471) begin
          $fatal; // @[Arbiter.scala 96:13:freechips.rocketchip.system.DefaultRV32Config.fir@6063.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_478) begin
          $fwrite(32'h80000002,"Assertion failed\n    at Arbiter.scala:98 assert (!earlyValids.reduce(_||_) || earlyWinner.reduce(_||_))\n"); // @[Arbiter.scala 98:14:freechips.rocketchip.system.DefaultRV32Config.fir@6073.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_478) begin
          $fatal; // @[Arbiter.scala 98:14:freechips.rocketchip.system.DefaultRV32Config.fir@6074.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_485) begin
          $fwrite(32'h80000002,"Assertion failed\n    at Arbiter.scala:99 assert (!validQuals .reduce(_||_) || validQuals .reduce(_||_))\n"); // @[Arbiter.scala 99:14:freechips.rocketchip.system.DefaultRV32Config.fir@6084.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_485) begin
          $fatal; // @[Arbiter.scala 99:14:freechips.rocketchip.system.DefaultRV32Config.fir@6085.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_623) begin
          $fwrite(32'h80000002,"Assertion failed\n    at Arbiter.scala:96 assert((prefixOR zip earlyWinner) map { case (p,w) => !p || !w } reduce {_ && _})\n"); // @[Arbiter.scala 96:13:freechips.rocketchip.system.DefaultRV32Config.fir@6321.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_623) begin
          $fatal; // @[Arbiter.scala 96:13:freechips.rocketchip.system.DefaultRV32Config.fir@6322.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_630) begin
          $fwrite(32'h80000002,"Assertion failed\n    at Arbiter.scala:98 assert (!earlyValids.reduce(_||_) || earlyWinner.reduce(_||_))\n"); // @[Arbiter.scala 98:14:freechips.rocketchip.system.DefaultRV32Config.fir@6332.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_630) begin
          $fatal; // @[Arbiter.scala 98:14:freechips.rocketchip.system.DefaultRV32Config.fir@6333.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_637) begin
          $fwrite(32'h80000002,"Assertion failed\n    at Arbiter.scala:99 assert (!validQuals .reduce(_||_) || validQuals .reduce(_||_))\n"); // @[Arbiter.scala 99:14:freechips.rocketchip.system.DefaultRV32Config.fir@6343.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_637) begin
          $fatal; // @[Arbiter.scala 99:14:freechips.rocketchip.system.DefaultRV32Config.fir@6344.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_777) begin
          $fwrite(32'h80000002,"Assertion failed\n    at Arbiter.scala:96 assert((prefixOR zip earlyWinner) map { case (p,w) => !p || !w } reduce {_ && _})\n"); // @[Arbiter.scala 96:13:freechips.rocketchip.system.DefaultRV32Config.fir@6596.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_777) begin
          $fatal; // @[Arbiter.scala 96:13:freechips.rocketchip.system.DefaultRV32Config.fir@6597.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_784) begin
          $fwrite(32'h80000002,"Assertion failed\n    at Arbiter.scala:98 assert (!earlyValids.reduce(_||_) || earlyWinner.reduce(_||_))\n"); // @[Arbiter.scala 98:14:freechips.rocketchip.system.DefaultRV32Config.fir@6607.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_784) begin
          $fatal; // @[Arbiter.scala 98:14:freechips.rocketchip.system.DefaultRV32Config.fir@6608.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_791) begin
          $fwrite(32'h80000002,"Assertion failed\n    at Arbiter.scala:99 assert (!validQuals .reduce(_||_) || validQuals .reduce(_||_))\n"); // @[Arbiter.scala 99:14:freechips.rocketchip.system.DefaultRV32Config.fir@6618.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_791) begin
          $fatal; // @[Arbiter.scala 99:14:freechips.rocketchip.system.DefaultRV32Config.fir@6619.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_953) begin
          $fwrite(32'h80000002,"Assertion failed\n    at Arbiter.scala:96 assert((prefixOR zip earlyWinner) map { case (p,w) => !p || !w } reduce {_ && _})\n"); // @[Arbiter.scala 96:13:freechips.rocketchip.system.DefaultRV32Config.fir@6945.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_953) begin
          $fatal; // @[Arbiter.scala 96:13:freechips.rocketchip.system.DefaultRV32Config.fir@6946.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_962) begin
          $fwrite(32'h80000002,"Assertion failed\n    at Arbiter.scala:98 assert (!earlyValids.reduce(_||_) || earlyWinner.reduce(_||_))\n"); // @[Arbiter.scala 98:14:freechips.rocketchip.system.DefaultRV32Config.fir@6958.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_962) begin
          $fatal; // @[Arbiter.scala 98:14:freechips.rocketchip.system.DefaultRV32Config.fir@6959.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_971) begin
          $fwrite(32'h80000002,"Assertion failed\n    at Arbiter.scala:99 assert (!validQuals .reduce(_||_) || validQuals .reduce(_||_))\n"); // @[Arbiter.scala 99:14:freechips.rocketchip.system.DefaultRV32Config.fir@6971.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_971) begin
          $fatal; // @[Arbiter.scala 99:14:freechips.rocketchip.system.DefaultRV32Config.fir@6972.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1125) begin
          $fwrite(32'h80000002,"Assertion failed\n    at Arbiter.scala:96 assert((prefixOR zip earlyWinner) map { case (p,w) => !p || !w } reduce {_ && _})\n"); // @[Arbiter.scala 96:13:freechips.rocketchip.system.DefaultRV32Config.fir@7274.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_1125) begin
          $fatal; // @[Arbiter.scala 96:13:freechips.rocketchip.system.DefaultRV32Config.fir@7275.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1134) begin
          $fwrite(32'h80000002,"Assertion failed\n    at Arbiter.scala:98 assert (!earlyValids.reduce(_||_) || earlyWinner.reduce(_||_))\n"); // @[Arbiter.scala 98:14:freechips.rocketchip.system.DefaultRV32Config.fir@7287.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_1134) begin
          $fatal; // @[Arbiter.scala 98:14:freechips.rocketchip.system.DefaultRV32Config.fir@7288.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1143) begin
          $fwrite(32'h80000002,"Assertion failed\n    at Arbiter.scala:99 assert (!validQuals .reduce(_||_) || validQuals .reduce(_||_))\n"); // @[Arbiter.scala 99:14:freechips.rocketchip.system.DefaultRV32Config.fir@7300.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_1143) begin
          $fatal; // @[Arbiter.scala 99:14:freechips.rocketchip.system.DefaultRV32Config.fir@7301.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
  end
endmodule
