module AXI4UserYanker( // @[:freechips.rocketchip.system.DefaultRV32Config.fir@23249.2]
  input         clock, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@23250.4]
  input         reset, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@23251.4]
  output        auto_in_aw_ready, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@23252.4]
  input         auto_in_aw_valid, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@23252.4]
  input  [3:0]  auto_in_aw_bits_id, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@23252.4]
  input  [30:0] auto_in_aw_bits_addr, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@23252.4]
  input  [7:0]  auto_in_aw_bits_len, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@23252.4]
  input  [2:0]  auto_in_aw_bits_size, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@23252.4]
  input  [1:0]  auto_in_aw_bits_burst, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@23252.4]
  input         auto_in_aw_bits_lock, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@23252.4]
  input  [3:0]  auto_in_aw_bits_cache, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@23252.4]
  input  [2:0]  auto_in_aw_bits_prot, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@23252.4]
  input  [3:0]  auto_in_aw_bits_qos, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@23252.4]
  input  [3:0]  auto_in_aw_bits_echo_tl_state_size, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@23252.4]
  input  [4:0]  auto_in_aw_bits_echo_tl_state_source, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@23252.4]
  output        auto_in_w_ready, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@23252.4]
  input         auto_in_w_valid, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@23252.4]
  input  [31:0] auto_in_w_bits_data, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@23252.4]
  input  [3:0]  auto_in_w_bits_strb, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@23252.4]
  input         auto_in_w_bits_last, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@23252.4]
  input         auto_in_b_ready, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@23252.4]
  output        auto_in_b_valid, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@23252.4]
  output [3:0]  auto_in_b_bits_id, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@23252.4]
  output [1:0]  auto_in_b_bits_resp, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@23252.4]
  output [3:0]  auto_in_b_bits_echo_tl_state_size, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@23252.4]
  output [4:0]  auto_in_b_bits_echo_tl_state_source, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@23252.4]
  output        auto_in_ar_ready, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@23252.4]
  input         auto_in_ar_valid, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@23252.4]
  input  [3:0]  auto_in_ar_bits_id, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@23252.4]
  input  [30:0] auto_in_ar_bits_addr, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@23252.4]
  input  [7:0]  auto_in_ar_bits_len, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@23252.4]
  input  [2:0]  auto_in_ar_bits_size, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@23252.4]
  input  [1:0]  auto_in_ar_bits_burst, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@23252.4]
  input         auto_in_ar_bits_lock, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@23252.4]
  input  [3:0]  auto_in_ar_bits_cache, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@23252.4]
  input  [2:0]  auto_in_ar_bits_prot, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@23252.4]
  input  [3:0]  auto_in_ar_bits_qos, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@23252.4]
  input  [3:0]  auto_in_ar_bits_echo_tl_state_size, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@23252.4]
  input  [4:0]  auto_in_ar_bits_echo_tl_state_source, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@23252.4]
  input         auto_in_r_ready, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@23252.4]
  output        auto_in_r_valid, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@23252.4]
  output [3:0]  auto_in_r_bits_id, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@23252.4]
  output [31:0] auto_in_r_bits_data, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@23252.4]
  output [1:0]  auto_in_r_bits_resp, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@23252.4]
  output [3:0]  auto_in_r_bits_echo_tl_state_size, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@23252.4]
  output [4:0]  auto_in_r_bits_echo_tl_state_source, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@23252.4]
  output        auto_in_r_bits_last, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@23252.4]
  input         auto_out_aw_ready, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@23252.4]
  output        auto_out_aw_valid, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@23252.4]
  output [3:0]  auto_out_aw_bits_id, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@23252.4]
  output [30:0] auto_out_aw_bits_addr, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@23252.4]
  output [7:0]  auto_out_aw_bits_len, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@23252.4]
  output [2:0]  auto_out_aw_bits_size, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@23252.4]
  output [1:0]  auto_out_aw_bits_burst, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@23252.4]
  output        auto_out_aw_bits_lock, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@23252.4]
  output [3:0]  auto_out_aw_bits_cache, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@23252.4]
  output [2:0]  auto_out_aw_bits_prot, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@23252.4]
  output [3:0]  auto_out_aw_bits_qos, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@23252.4]
  input         auto_out_w_ready, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@23252.4]
  output        auto_out_w_valid, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@23252.4]
  output [31:0] auto_out_w_bits_data, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@23252.4]
  output [3:0]  auto_out_w_bits_strb, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@23252.4]
  output        auto_out_w_bits_last, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@23252.4]
  output        auto_out_b_ready, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@23252.4]
  input         auto_out_b_valid, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@23252.4]
  input  [3:0]  auto_out_b_bits_id, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@23252.4]
  input  [1:0]  auto_out_b_bits_resp, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@23252.4]
  input         auto_out_ar_ready, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@23252.4]
  output        auto_out_ar_valid, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@23252.4]
  output [3:0]  auto_out_ar_bits_id, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@23252.4]
  output [30:0] auto_out_ar_bits_addr, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@23252.4]
  output [7:0]  auto_out_ar_bits_len, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@23252.4]
  output [2:0]  auto_out_ar_bits_size, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@23252.4]
  output [1:0]  auto_out_ar_bits_burst, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@23252.4]
  output        auto_out_ar_bits_lock, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@23252.4]
  output [3:0]  auto_out_ar_bits_cache, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@23252.4]
  output [2:0]  auto_out_ar_bits_prot, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@23252.4]
  output [3:0]  auto_out_ar_bits_qos, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@23252.4]
  output        auto_out_r_ready, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@23252.4]
  input         auto_out_r_valid, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@23252.4]
  input  [3:0]  auto_out_r_bits_id, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@23252.4]
  input  [31:0] auto_out_r_bits_data, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@23252.4]
  input  [1:0]  auto_out_r_bits_resp, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@23252.4]
  input         auto_out_r_bits_last // @[:freechips.rocketchip.system.DefaultRV32Config.fir@23252.4]
);
  wire  QueueCompatibility_clock; // @[UserYanker.scala 39:17:freechips.rocketchip.system.DefaultRV32Config.fir@23263.4]
  wire  QueueCompatibility_reset; // @[UserYanker.scala 39:17:freechips.rocketchip.system.DefaultRV32Config.fir@23263.4]
  wire  QueueCompatibility_io_enq_ready; // @[UserYanker.scala 39:17:freechips.rocketchip.system.DefaultRV32Config.fir@23263.4]
  wire  QueueCompatibility_io_enq_valid; // @[UserYanker.scala 39:17:freechips.rocketchip.system.DefaultRV32Config.fir@23263.4]
  wire [3:0] QueueCompatibility_io_enq_bits_tl_state_size; // @[UserYanker.scala 39:17:freechips.rocketchip.system.DefaultRV32Config.fir@23263.4]
  wire [4:0] QueueCompatibility_io_enq_bits_tl_state_source; // @[UserYanker.scala 39:17:freechips.rocketchip.system.DefaultRV32Config.fir@23263.4]
  wire  QueueCompatibility_io_deq_ready; // @[UserYanker.scala 39:17:freechips.rocketchip.system.DefaultRV32Config.fir@23263.4]
  wire  QueueCompatibility_io_deq_valid; // @[UserYanker.scala 39:17:freechips.rocketchip.system.DefaultRV32Config.fir@23263.4]
  wire [3:0] QueueCompatibility_io_deq_bits_tl_state_size; // @[UserYanker.scala 39:17:freechips.rocketchip.system.DefaultRV32Config.fir@23263.4]
  wire [4:0] QueueCompatibility_io_deq_bits_tl_state_source; // @[UserYanker.scala 39:17:freechips.rocketchip.system.DefaultRV32Config.fir@23263.4]
  wire  QueueCompatibility_1_clock; // @[UserYanker.scala 39:17:freechips.rocketchip.system.DefaultRV32Config.fir@23267.4]
  wire  QueueCompatibility_1_reset; // @[UserYanker.scala 39:17:freechips.rocketchip.system.DefaultRV32Config.fir@23267.4]
  wire  QueueCompatibility_1_io_enq_ready; // @[UserYanker.scala 39:17:freechips.rocketchip.system.DefaultRV32Config.fir@23267.4]
  wire  QueueCompatibility_1_io_enq_valid; // @[UserYanker.scala 39:17:freechips.rocketchip.system.DefaultRV32Config.fir@23267.4]
  wire [3:0] QueueCompatibility_1_io_enq_bits_tl_state_size; // @[UserYanker.scala 39:17:freechips.rocketchip.system.DefaultRV32Config.fir@23267.4]
  wire [4:0] QueueCompatibility_1_io_enq_bits_tl_state_source; // @[UserYanker.scala 39:17:freechips.rocketchip.system.DefaultRV32Config.fir@23267.4]
  wire  QueueCompatibility_1_io_deq_ready; // @[UserYanker.scala 39:17:freechips.rocketchip.system.DefaultRV32Config.fir@23267.4]
  wire  QueueCompatibility_1_io_deq_valid; // @[UserYanker.scala 39:17:freechips.rocketchip.system.DefaultRV32Config.fir@23267.4]
  wire [3:0] QueueCompatibility_1_io_deq_bits_tl_state_size; // @[UserYanker.scala 39:17:freechips.rocketchip.system.DefaultRV32Config.fir@23267.4]
  wire [4:0] QueueCompatibility_1_io_deq_bits_tl_state_source; // @[UserYanker.scala 39:17:freechips.rocketchip.system.DefaultRV32Config.fir@23267.4]
  wire  QueueCompatibility_2_clock; // @[UserYanker.scala 39:17:freechips.rocketchip.system.DefaultRV32Config.fir@23271.4]
  wire  QueueCompatibility_2_reset; // @[UserYanker.scala 39:17:freechips.rocketchip.system.DefaultRV32Config.fir@23271.4]
  wire  QueueCompatibility_2_io_enq_ready; // @[UserYanker.scala 39:17:freechips.rocketchip.system.DefaultRV32Config.fir@23271.4]
  wire  QueueCompatibility_2_io_enq_valid; // @[UserYanker.scala 39:17:freechips.rocketchip.system.DefaultRV32Config.fir@23271.4]
  wire [3:0] QueueCompatibility_2_io_enq_bits_tl_state_size; // @[UserYanker.scala 39:17:freechips.rocketchip.system.DefaultRV32Config.fir@23271.4]
  wire [4:0] QueueCompatibility_2_io_enq_bits_tl_state_source; // @[UserYanker.scala 39:17:freechips.rocketchip.system.DefaultRV32Config.fir@23271.4]
  wire  QueueCompatibility_2_io_deq_ready; // @[UserYanker.scala 39:17:freechips.rocketchip.system.DefaultRV32Config.fir@23271.4]
  wire  QueueCompatibility_2_io_deq_valid; // @[UserYanker.scala 39:17:freechips.rocketchip.system.DefaultRV32Config.fir@23271.4]
  wire [3:0] QueueCompatibility_2_io_deq_bits_tl_state_size; // @[UserYanker.scala 39:17:freechips.rocketchip.system.DefaultRV32Config.fir@23271.4]
  wire [4:0] QueueCompatibility_2_io_deq_bits_tl_state_source; // @[UserYanker.scala 39:17:freechips.rocketchip.system.DefaultRV32Config.fir@23271.4]
  wire  QueueCompatibility_3_clock; // @[UserYanker.scala 39:17:freechips.rocketchip.system.DefaultRV32Config.fir@23275.4]
  wire  QueueCompatibility_3_reset; // @[UserYanker.scala 39:17:freechips.rocketchip.system.DefaultRV32Config.fir@23275.4]
  wire  QueueCompatibility_3_io_enq_ready; // @[UserYanker.scala 39:17:freechips.rocketchip.system.DefaultRV32Config.fir@23275.4]
  wire  QueueCompatibility_3_io_enq_valid; // @[UserYanker.scala 39:17:freechips.rocketchip.system.DefaultRV32Config.fir@23275.4]
  wire [3:0] QueueCompatibility_3_io_enq_bits_tl_state_size; // @[UserYanker.scala 39:17:freechips.rocketchip.system.DefaultRV32Config.fir@23275.4]
  wire [4:0] QueueCompatibility_3_io_enq_bits_tl_state_source; // @[UserYanker.scala 39:17:freechips.rocketchip.system.DefaultRV32Config.fir@23275.4]
  wire  QueueCompatibility_3_io_deq_ready; // @[UserYanker.scala 39:17:freechips.rocketchip.system.DefaultRV32Config.fir@23275.4]
  wire  QueueCompatibility_3_io_deq_valid; // @[UserYanker.scala 39:17:freechips.rocketchip.system.DefaultRV32Config.fir@23275.4]
  wire [3:0] QueueCompatibility_3_io_deq_bits_tl_state_size; // @[UserYanker.scala 39:17:freechips.rocketchip.system.DefaultRV32Config.fir@23275.4]
  wire [4:0] QueueCompatibility_3_io_deq_bits_tl_state_source; // @[UserYanker.scala 39:17:freechips.rocketchip.system.DefaultRV32Config.fir@23275.4]
  wire  QueueCompatibility_4_clock; // @[UserYanker.scala 39:17:freechips.rocketchip.system.DefaultRV32Config.fir@23279.4]
  wire  QueueCompatibility_4_reset; // @[UserYanker.scala 39:17:freechips.rocketchip.system.DefaultRV32Config.fir@23279.4]
  wire  QueueCompatibility_4_io_enq_ready; // @[UserYanker.scala 39:17:freechips.rocketchip.system.DefaultRV32Config.fir@23279.4]
  wire  QueueCompatibility_4_io_enq_valid; // @[UserYanker.scala 39:17:freechips.rocketchip.system.DefaultRV32Config.fir@23279.4]
  wire [3:0] QueueCompatibility_4_io_enq_bits_tl_state_size; // @[UserYanker.scala 39:17:freechips.rocketchip.system.DefaultRV32Config.fir@23279.4]
  wire [4:0] QueueCompatibility_4_io_enq_bits_tl_state_source; // @[UserYanker.scala 39:17:freechips.rocketchip.system.DefaultRV32Config.fir@23279.4]
  wire  QueueCompatibility_4_io_deq_ready; // @[UserYanker.scala 39:17:freechips.rocketchip.system.DefaultRV32Config.fir@23279.4]
  wire  QueueCompatibility_4_io_deq_valid; // @[UserYanker.scala 39:17:freechips.rocketchip.system.DefaultRV32Config.fir@23279.4]
  wire [3:0] QueueCompatibility_4_io_deq_bits_tl_state_size; // @[UserYanker.scala 39:17:freechips.rocketchip.system.DefaultRV32Config.fir@23279.4]
  wire [4:0] QueueCompatibility_4_io_deq_bits_tl_state_source; // @[UserYanker.scala 39:17:freechips.rocketchip.system.DefaultRV32Config.fir@23279.4]
  wire  QueueCompatibility_5_clock; // @[UserYanker.scala 39:17:freechips.rocketchip.system.DefaultRV32Config.fir@23305.4]
  wire  QueueCompatibility_5_reset; // @[UserYanker.scala 39:17:freechips.rocketchip.system.DefaultRV32Config.fir@23305.4]
  wire  QueueCompatibility_5_io_enq_ready; // @[UserYanker.scala 39:17:freechips.rocketchip.system.DefaultRV32Config.fir@23305.4]
  wire  QueueCompatibility_5_io_enq_valid; // @[UserYanker.scala 39:17:freechips.rocketchip.system.DefaultRV32Config.fir@23305.4]
  wire [3:0] QueueCompatibility_5_io_enq_bits_tl_state_size; // @[UserYanker.scala 39:17:freechips.rocketchip.system.DefaultRV32Config.fir@23305.4]
  wire [4:0] QueueCompatibility_5_io_enq_bits_tl_state_source; // @[UserYanker.scala 39:17:freechips.rocketchip.system.DefaultRV32Config.fir@23305.4]
  wire  QueueCompatibility_5_io_deq_ready; // @[UserYanker.scala 39:17:freechips.rocketchip.system.DefaultRV32Config.fir@23305.4]
  wire  QueueCompatibility_5_io_deq_valid; // @[UserYanker.scala 39:17:freechips.rocketchip.system.DefaultRV32Config.fir@23305.4]
  wire [3:0] QueueCompatibility_5_io_deq_bits_tl_state_size; // @[UserYanker.scala 39:17:freechips.rocketchip.system.DefaultRV32Config.fir@23305.4]
  wire [4:0] QueueCompatibility_5_io_deq_bits_tl_state_source; // @[UserYanker.scala 39:17:freechips.rocketchip.system.DefaultRV32Config.fir@23305.4]
  wire  QueueCompatibility_6_clock; // @[UserYanker.scala 39:17:freechips.rocketchip.system.DefaultRV32Config.fir@23309.4]
  wire  QueueCompatibility_6_reset; // @[UserYanker.scala 39:17:freechips.rocketchip.system.DefaultRV32Config.fir@23309.4]
  wire  QueueCompatibility_6_io_enq_ready; // @[UserYanker.scala 39:17:freechips.rocketchip.system.DefaultRV32Config.fir@23309.4]
  wire  QueueCompatibility_6_io_enq_valid; // @[UserYanker.scala 39:17:freechips.rocketchip.system.DefaultRV32Config.fir@23309.4]
  wire [3:0] QueueCompatibility_6_io_enq_bits_tl_state_size; // @[UserYanker.scala 39:17:freechips.rocketchip.system.DefaultRV32Config.fir@23309.4]
  wire [4:0] QueueCompatibility_6_io_enq_bits_tl_state_source; // @[UserYanker.scala 39:17:freechips.rocketchip.system.DefaultRV32Config.fir@23309.4]
  wire  QueueCompatibility_6_io_deq_ready; // @[UserYanker.scala 39:17:freechips.rocketchip.system.DefaultRV32Config.fir@23309.4]
  wire  QueueCompatibility_6_io_deq_valid; // @[UserYanker.scala 39:17:freechips.rocketchip.system.DefaultRV32Config.fir@23309.4]
  wire [3:0] QueueCompatibility_6_io_deq_bits_tl_state_size; // @[UserYanker.scala 39:17:freechips.rocketchip.system.DefaultRV32Config.fir@23309.4]
  wire [4:0] QueueCompatibility_6_io_deq_bits_tl_state_source; // @[UserYanker.scala 39:17:freechips.rocketchip.system.DefaultRV32Config.fir@23309.4]
  wire  QueueCompatibility_7_clock; // @[UserYanker.scala 39:17:freechips.rocketchip.system.DefaultRV32Config.fir@23313.4]
  wire  QueueCompatibility_7_reset; // @[UserYanker.scala 39:17:freechips.rocketchip.system.DefaultRV32Config.fir@23313.4]
  wire  QueueCompatibility_7_io_enq_ready; // @[UserYanker.scala 39:17:freechips.rocketchip.system.DefaultRV32Config.fir@23313.4]
  wire  QueueCompatibility_7_io_enq_valid; // @[UserYanker.scala 39:17:freechips.rocketchip.system.DefaultRV32Config.fir@23313.4]
  wire [3:0] QueueCompatibility_7_io_enq_bits_tl_state_size; // @[UserYanker.scala 39:17:freechips.rocketchip.system.DefaultRV32Config.fir@23313.4]
  wire [4:0] QueueCompatibility_7_io_enq_bits_tl_state_source; // @[UserYanker.scala 39:17:freechips.rocketchip.system.DefaultRV32Config.fir@23313.4]
  wire  QueueCompatibility_7_io_deq_ready; // @[UserYanker.scala 39:17:freechips.rocketchip.system.DefaultRV32Config.fir@23313.4]
  wire  QueueCompatibility_7_io_deq_valid; // @[UserYanker.scala 39:17:freechips.rocketchip.system.DefaultRV32Config.fir@23313.4]
  wire [3:0] QueueCompatibility_7_io_deq_bits_tl_state_size; // @[UserYanker.scala 39:17:freechips.rocketchip.system.DefaultRV32Config.fir@23313.4]
  wire [4:0] QueueCompatibility_7_io_deq_bits_tl_state_source; // @[UserYanker.scala 39:17:freechips.rocketchip.system.DefaultRV32Config.fir@23313.4]
  wire  QueueCompatibility_8_clock; // @[UserYanker.scala 39:17:freechips.rocketchip.system.DefaultRV32Config.fir@23317.4]
  wire  QueueCompatibility_8_reset; // @[UserYanker.scala 39:17:freechips.rocketchip.system.DefaultRV32Config.fir@23317.4]
  wire  QueueCompatibility_8_io_enq_ready; // @[UserYanker.scala 39:17:freechips.rocketchip.system.DefaultRV32Config.fir@23317.4]
  wire  QueueCompatibility_8_io_enq_valid; // @[UserYanker.scala 39:17:freechips.rocketchip.system.DefaultRV32Config.fir@23317.4]
  wire [3:0] QueueCompatibility_8_io_enq_bits_tl_state_size; // @[UserYanker.scala 39:17:freechips.rocketchip.system.DefaultRV32Config.fir@23317.4]
  wire [4:0] QueueCompatibility_8_io_enq_bits_tl_state_source; // @[UserYanker.scala 39:17:freechips.rocketchip.system.DefaultRV32Config.fir@23317.4]
  wire  QueueCompatibility_8_io_deq_ready; // @[UserYanker.scala 39:17:freechips.rocketchip.system.DefaultRV32Config.fir@23317.4]
  wire  QueueCompatibility_8_io_deq_valid; // @[UserYanker.scala 39:17:freechips.rocketchip.system.DefaultRV32Config.fir@23317.4]
  wire [3:0] QueueCompatibility_8_io_deq_bits_tl_state_size; // @[UserYanker.scala 39:17:freechips.rocketchip.system.DefaultRV32Config.fir@23317.4]
  wire [4:0] QueueCompatibility_8_io_deq_bits_tl_state_source; // @[UserYanker.scala 39:17:freechips.rocketchip.system.DefaultRV32Config.fir@23317.4]
  wire  QueueCompatibility_9_clock; // @[UserYanker.scala 39:17:freechips.rocketchip.system.DefaultRV32Config.fir@23321.4]
  wire  QueueCompatibility_9_reset; // @[UserYanker.scala 39:17:freechips.rocketchip.system.DefaultRV32Config.fir@23321.4]
  wire  QueueCompatibility_9_io_enq_ready; // @[UserYanker.scala 39:17:freechips.rocketchip.system.DefaultRV32Config.fir@23321.4]
  wire  QueueCompatibility_9_io_enq_valid; // @[UserYanker.scala 39:17:freechips.rocketchip.system.DefaultRV32Config.fir@23321.4]
  wire [3:0] QueueCompatibility_9_io_enq_bits_tl_state_size; // @[UserYanker.scala 39:17:freechips.rocketchip.system.DefaultRV32Config.fir@23321.4]
  wire [4:0] QueueCompatibility_9_io_enq_bits_tl_state_source; // @[UserYanker.scala 39:17:freechips.rocketchip.system.DefaultRV32Config.fir@23321.4]
  wire  QueueCompatibility_9_io_deq_ready; // @[UserYanker.scala 39:17:freechips.rocketchip.system.DefaultRV32Config.fir@23321.4]
  wire  QueueCompatibility_9_io_deq_valid; // @[UserYanker.scala 39:17:freechips.rocketchip.system.DefaultRV32Config.fir@23321.4]
  wire [3:0] QueueCompatibility_9_io_deq_bits_tl_state_size; // @[UserYanker.scala 39:17:freechips.rocketchip.system.DefaultRV32Config.fir@23321.4]
  wire [4:0] QueueCompatibility_9_io_deq_bits_tl_state_source; // @[UserYanker.scala 39:17:freechips.rocketchip.system.DefaultRV32Config.fir@23321.4]
  wire  _T_24_0; // @[UserYanker.scala 47:25:freechips.rocketchip.system.DefaultRV32Config.fir@23347.4 UserYanker.scala 47:25:freechips.rocketchip.system.DefaultRV32Config.fir@23349.4]
  wire  _T_24_1; // @[UserYanker.scala 47:25:freechips.rocketchip.system.DefaultRV32Config.fir@23347.4 UserYanker.scala 47:25:freechips.rocketchip.system.DefaultRV32Config.fir@23350.4]
  wire  _GEN_1; // @[UserYanker.scala 48:36:freechips.rocketchip.system.DefaultRV32Config.fir@23365.4]
  wire  _T_24_2; // @[UserYanker.scala 47:25:freechips.rocketchip.system.DefaultRV32Config.fir@23347.4 UserYanker.scala 47:25:freechips.rocketchip.system.DefaultRV32Config.fir@23351.4]
  wire  _GEN_2; // @[UserYanker.scala 48:36:freechips.rocketchip.system.DefaultRV32Config.fir@23365.4]
  wire  _T_24_3; // @[UserYanker.scala 47:25:freechips.rocketchip.system.DefaultRV32Config.fir@23347.4 UserYanker.scala 47:25:freechips.rocketchip.system.DefaultRV32Config.fir@23352.4]
  wire  _GEN_3; // @[UserYanker.scala 48:36:freechips.rocketchip.system.DefaultRV32Config.fir@23365.4]
  wire  _T_24_4; // @[UserYanker.scala 47:25:freechips.rocketchip.system.DefaultRV32Config.fir@23347.4 UserYanker.scala 47:25:freechips.rocketchip.system.DefaultRV32Config.fir@23353.4]
  wire  _GEN_4; // @[UserYanker.scala 48:36:freechips.rocketchip.system.DefaultRV32Config.fir@23365.4]
  wire  _GEN_5; // @[UserYanker.scala 48:36:freechips.rocketchip.system.DefaultRV32Config.fir@23365.4]
  wire  _GEN_6; // @[UserYanker.scala 48:36:freechips.rocketchip.system.DefaultRV32Config.fir@23365.4]
  wire  _GEN_7; // @[UserYanker.scala 48:36:freechips.rocketchip.system.DefaultRV32Config.fir@23365.4]
  wire  _GEN_8; // @[UserYanker.scala 48:36:freechips.rocketchip.system.DefaultRV32Config.fir@23365.4]
  wire  _GEN_9; // @[UserYanker.scala 48:36:freechips.rocketchip.system.DefaultRV32Config.fir@23365.4]
  wire  _GEN_10; // @[UserYanker.scala 48:36:freechips.rocketchip.system.DefaultRV32Config.fir@23365.4]
  wire  _GEN_11; // @[UserYanker.scala 48:36:freechips.rocketchip.system.DefaultRV32Config.fir@23365.4]
  wire  _GEN_12; // @[UserYanker.scala 48:36:freechips.rocketchip.system.DefaultRV32Config.fir@23365.4]
  wire  _GEN_13; // @[UserYanker.scala 48:36:freechips.rocketchip.system.DefaultRV32Config.fir@23365.4]
  wire  _GEN_14; // @[UserYanker.scala 48:36:freechips.rocketchip.system.DefaultRV32Config.fir@23365.4]
  wire  _GEN_15; // @[UserYanker.scala 48:36:freechips.rocketchip.system.DefaultRV32Config.fir@23365.4]
  wire  _T_29; // @[UserYanker.scala 55:15:freechips.rocketchip.system.DefaultRV32Config.fir@23414.4]
  wire  _T_27_0; // @[UserYanker.scala 53:24:freechips.rocketchip.system.DefaultRV32Config.fir@23378.4 UserYanker.scala 53:24:freechips.rocketchip.system.DefaultRV32Config.fir@23380.4]
  wire  _T_27_1; // @[UserYanker.scala 53:24:freechips.rocketchip.system.DefaultRV32Config.fir@23378.4 UserYanker.scala 53:24:freechips.rocketchip.system.DefaultRV32Config.fir@23381.4]
  wire  _GEN_17; // @[UserYanker.scala 55:28:freechips.rocketchip.system.DefaultRV32Config.fir@23415.4]
  wire  _T_27_2; // @[UserYanker.scala 53:24:freechips.rocketchip.system.DefaultRV32Config.fir@23378.4 UserYanker.scala 53:24:freechips.rocketchip.system.DefaultRV32Config.fir@23382.4]
  wire  _GEN_18; // @[UserYanker.scala 55:28:freechips.rocketchip.system.DefaultRV32Config.fir@23415.4]
  wire  _T_27_3; // @[UserYanker.scala 53:24:freechips.rocketchip.system.DefaultRV32Config.fir@23378.4 UserYanker.scala 53:24:freechips.rocketchip.system.DefaultRV32Config.fir@23383.4]
  wire  _GEN_19; // @[UserYanker.scala 55:28:freechips.rocketchip.system.DefaultRV32Config.fir@23415.4]
  wire  _T_27_4; // @[UserYanker.scala 53:24:freechips.rocketchip.system.DefaultRV32Config.fir@23378.4 UserYanker.scala 53:24:freechips.rocketchip.system.DefaultRV32Config.fir@23384.4]
  wire  _GEN_20; // @[UserYanker.scala 55:28:freechips.rocketchip.system.DefaultRV32Config.fir@23415.4]
  wire  _GEN_21; // @[UserYanker.scala 55:28:freechips.rocketchip.system.DefaultRV32Config.fir@23415.4]
  wire  _GEN_22; // @[UserYanker.scala 55:28:freechips.rocketchip.system.DefaultRV32Config.fir@23415.4]
  wire  _GEN_23; // @[UserYanker.scala 55:28:freechips.rocketchip.system.DefaultRV32Config.fir@23415.4]
  wire  _GEN_24; // @[UserYanker.scala 55:28:freechips.rocketchip.system.DefaultRV32Config.fir@23415.4]
  wire  _GEN_25; // @[UserYanker.scala 55:28:freechips.rocketchip.system.DefaultRV32Config.fir@23415.4]
  wire  _GEN_26; // @[UserYanker.scala 55:28:freechips.rocketchip.system.DefaultRV32Config.fir@23415.4]
  wire  _GEN_27; // @[UserYanker.scala 55:28:freechips.rocketchip.system.DefaultRV32Config.fir@23415.4]
  wire  _GEN_28; // @[UserYanker.scala 55:28:freechips.rocketchip.system.DefaultRV32Config.fir@23415.4]
  wire  _GEN_29; // @[UserYanker.scala 55:28:freechips.rocketchip.system.DefaultRV32Config.fir@23415.4]
  wire  _GEN_30; // @[UserYanker.scala 55:28:freechips.rocketchip.system.DefaultRV32Config.fir@23415.4]
  wire  _GEN_31; // @[UserYanker.scala 55:28:freechips.rocketchip.system.DefaultRV32Config.fir@23415.4]
  wire  _T_30; // @[UserYanker.scala 55:28:freechips.rocketchip.system.DefaultRV32Config.fir@23415.4]
  wire  _T_32; // @[UserYanker.scala 55:14:freechips.rocketchip.system.DefaultRV32Config.fir@23417.4]
  wire  _T_33; // @[UserYanker.scala 55:14:freechips.rocketchip.system.DefaultRV32Config.fir@23418.4]
  wire [3:0] _T_28_0_tl_state_size; // @[UserYanker.scala 54:23:freechips.rocketchip.system.DefaultRV32Config.fir@23396.4 UserYanker.scala 54:23:freechips.rocketchip.system.DefaultRV32Config.fir@23398.4]
  wire [4:0] _T_28_0_tl_state_source; // @[UserYanker.scala 54:23:freechips.rocketchip.system.DefaultRV32Config.fir@23396.4 UserYanker.scala 54:23:freechips.rocketchip.system.DefaultRV32Config.fir@23398.4]
  wire [3:0] _T_28_1_tl_state_size; // @[UserYanker.scala 54:23:freechips.rocketchip.system.DefaultRV32Config.fir@23396.4 UserYanker.scala 54:23:freechips.rocketchip.system.DefaultRV32Config.fir@23399.4]
  wire [3:0] _GEN_34; // @[BundleMap.scala 248:19:freechips.rocketchip.system.DefaultRV32Config.fir@23431.4]
  wire [4:0] _T_28_1_tl_state_source; // @[UserYanker.scala 54:23:freechips.rocketchip.system.DefaultRV32Config.fir@23396.4 UserYanker.scala 54:23:freechips.rocketchip.system.DefaultRV32Config.fir@23399.4]
  wire [4:0] _GEN_35; // @[BundleMap.scala 248:19:freechips.rocketchip.system.DefaultRV32Config.fir@23431.4]
  wire [3:0] _T_28_2_tl_state_size; // @[UserYanker.scala 54:23:freechips.rocketchip.system.DefaultRV32Config.fir@23396.4 UserYanker.scala 54:23:freechips.rocketchip.system.DefaultRV32Config.fir@23400.4]
  wire [3:0] _GEN_36; // @[BundleMap.scala 248:19:freechips.rocketchip.system.DefaultRV32Config.fir@23431.4]
  wire [4:0] _T_28_2_tl_state_source; // @[UserYanker.scala 54:23:freechips.rocketchip.system.DefaultRV32Config.fir@23396.4 UserYanker.scala 54:23:freechips.rocketchip.system.DefaultRV32Config.fir@23400.4]
  wire [4:0] _GEN_37; // @[BundleMap.scala 248:19:freechips.rocketchip.system.DefaultRV32Config.fir@23431.4]
  wire [3:0] _T_28_3_tl_state_size; // @[UserYanker.scala 54:23:freechips.rocketchip.system.DefaultRV32Config.fir@23396.4 UserYanker.scala 54:23:freechips.rocketchip.system.DefaultRV32Config.fir@23401.4]
  wire [3:0] _GEN_38; // @[BundleMap.scala 248:19:freechips.rocketchip.system.DefaultRV32Config.fir@23431.4]
  wire [4:0] _T_28_3_tl_state_source; // @[UserYanker.scala 54:23:freechips.rocketchip.system.DefaultRV32Config.fir@23396.4 UserYanker.scala 54:23:freechips.rocketchip.system.DefaultRV32Config.fir@23401.4]
  wire [4:0] _GEN_39; // @[BundleMap.scala 248:19:freechips.rocketchip.system.DefaultRV32Config.fir@23431.4]
  wire [3:0] _T_28_4_tl_state_size; // @[UserYanker.scala 54:23:freechips.rocketchip.system.DefaultRV32Config.fir@23396.4 UserYanker.scala 54:23:freechips.rocketchip.system.DefaultRV32Config.fir@23402.4]
  wire [3:0] _GEN_40; // @[BundleMap.scala 248:19:freechips.rocketchip.system.DefaultRV32Config.fir@23431.4]
  wire [4:0] _T_28_4_tl_state_source; // @[UserYanker.scala 54:23:freechips.rocketchip.system.DefaultRV32Config.fir@23396.4 UserYanker.scala 54:23:freechips.rocketchip.system.DefaultRV32Config.fir@23402.4]
  wire [4:0] _GEN_41; // @[BundleMap.scala 248:19:freechips.rocketchip.system.DefaultRV32Config.fir@23431.4]
  wire [3:0] _GEN_42; // @[BundleMap.scala 248:19:freechips.rocketchip.system.DefaultRV32Config.fir@23431.4]
  wire [4:0] _GEN_43; // @[BundleMap.scala 248:19:freechips.rocketchip.system.DefaultRV32Config.fir@23431.4]
  wire [3:0] _GEN_44; // @[BundleMap.scala 248:19:freechips.rocketchip.system.DefaultRV32Config.fir@23431.4]
  wire [4:0] _GEN_45; // @[BundleMap.scala 248:19:freechips.rocketchip.system.DefaultRV32Config.fir@23431.4]
  wire [3:0] _GEN_46; // @[BundleMap.scala 248:19:freechips.rocketchip.system.DefaultRV32Config.fir@23431.4]
  wire [4:0] _GEN_47; // @[BundleMap.scala 248:19:freechips.rocketchip.system.DefaultRV32Config.fir@23431.4]
  wire [3:0] _GEN_48; // @[BundleMap.scala 248:19:freechips.rocketchip.system.DefaultRV32Config.fir@23431.4]
  wire [4:0] _GEN_49; // @[BundleMap.scala 248:19:freechips.rocketchip.system.DefaultRV32Config.fir@23431.4]
  wire [3:0] _GEN_50; // @[BundleMap.scala 248:19:freechips.rocketchip.system.DefaultRV32Config.fir@23431.4]
  wire [4:0] _GEN_51; // @[BundleMap.scala 248:19:freechips.rocketchip.system.DefaultRV32Config.fir@23431.4]
  wire [3:0] _GEN_52; // @[BundleMap.scala 248:19:freechips.rocketchip.system.DefaultRV32Config.fir@23431.4]
  wire [4:0] _GEN_53; // @[BundleMap.scala 248:19:freechips.rocketchip.system.DefaultRV32Config.fir@23431.4]
  wire [3:0] _GEN_54; // @[BundleMap.scala 248:19:freechips.rocketchip.system.DefaultRV32Config.fir@23431.4]
  wire [4:0] _GEN_55; // @[BundleMap.scala 248:19:freechips.rocketchip.system.DefaultRV32Config.fir@23431.4]
  wire [3:0] _GEN_56; // @[BundleMap.scala 248:19:freechips.rocketchip.system.DefaultRV32Config.fir@23431.4]
  wire [4:0] _GEN_57; // @[BundleMap.scala 248:19:freechips.rocketchip.system.DefaultRV32Config.fir@23431.4]
  wire [3:0] _GEN_58; // @[BundleMap.scala 248:19:freechips.rocketchip.system.DefaultRV32Config.fir@23431.4]
  wire [4:0] _GEN_59; // @[BundleMap.scala 248:19:freechips.rocketchip.system.DefaultRV32Config.fir@23431.4]
  wire [3:0] _GEN_60; // @[BundleMap.scala 248:19:freechips.rocketchip.system.DefaultRV32Config.fir@23431.4]
  wire [4:0] _GEN_61; // @[BundleMap.scala 248:19:freechips.rocketchip.system.DefaultRV32Config.fir@23431.4]
  wire [15:0] _T_35; // @[OneHot.scala 65:12:freechips.rocketchip.system.DefaultRV32Config.fir@23434.4]
  wire [15:0] _T_54; // @[OneHot.scala 65:12:freechips.rocketchip.system.DefaultRV32Config.fir@23453.4]
  wire  _T_72; // @[UserYanker.scala 62:37:freechips.rocketchip.system.DefaultRV32Config.fir@23471.4]
  wire  _T_73; // @[UserYanker.scala 62:53:freechips.rocketchip.system.DefaultRV32Config.fir@23472.4]
  wire  _T_75; // @[UserYanker.scala 63:37:freechips.rocketchip.system.DefaultRV32Config.fir@23475.4]
  wire  _T_78; // @[UserYanker.scala 62:53:freechips.rocketchip.system.DefaultRV32Config.fir@23481.4]
  wire  _T_83; // @[UserYanker.scala 62:53:freechips.rocketchip.system.DefaultRV32Config.fir@23490.4]
  wire  _T_88; // @[UserYanker.scala 62:53:freechips.rocketchip.system.DefaultRV32Config.fir@23499.4]
  wire  _T_93; // @[UserYanker.scala 62:53:freechips.rocketchip.system.DefaultRV32Config.fir@23508.4]
  wire  _T_152_0; // @[UserYanker.scala 68:25:freechips.rocketchip.system.DefaultRV32Config.fir@23615.4 UserYanker.scala 68:25:freechips.rocketchip.system.DefaultRV32Config.fir@23617.4]
  wire  _T_152_1; // @[UserYanker.scala 68:25:freechips.rocketchip.system.DefaultRV32Config.fir@23615.4 UserYanker.scala 68:25:freechips.rocketchip.system.DefaultRV32Config.fir@23618.4]
  wire  _GEN_65; // @[UserYanker.scala 69:36:freechips.rocketchip.system.DefaultRV32Config.fir@23633.4]
  wire  _T_152_2; // @[UserYanker.scala 68:25:freechips.rocketchip.system.DefaultRV32Config.fir@23615.4 UserYanker.scala 68:25:freechips.rocketchip.system.DefaultRV32Config.fir@23619.4]
  wire  _GEN_66; // @[UserYanker.scala 69:36:freechips.rocketchip.system.DefaultRV32Config.fir@23633.4]
  wire  _T_152_3; // @[UserYanker.scala 68:25:freechips.rocketchip.system.DefaultRV32Config.fir@23615.4 UserYanker.scala 68:25:freechips.rocketchip.system.DefaultRV32Config.fir@23620.4]
  wire  _GEN_67; // @[UserYanker.scala 69:36:freechips.rocketchip.system.DefaultRV32Config.fir@23633.4]
  wire  _T_152_4; // @[UserYanker.scala 68:25:freechips.rocketchip.system.DefaultRV32Config.fir@23615.4 UserYanker.scala 68:25:freechips.rocketchip.system.DefaultRV32Config.fir@23621.4]
  wire  _GEN_68; // @[UserYanker.scala 69:36:freechips.rocketchip.system.DefaultRV32Config.fir@23633.4]
  wire  _GEN_69; // @[UserYanker.scala 69:36:freechips.rocketchip.system.DefaultRV32Config.fir@23633.4]
  wire  _GEN_70; // @[UserYanker.scala 69:36:freechips.rocketchip.system.DefaultRV32Config.fir@23633.4]
  wire  _GEN_71; // @[UserYanker.scala 69:36:freechips.rocketchip.system.DefaultRV32Config.fir@23633.4]
  wire  _GEN_72; // @[UserYanker.scala 69:36:freechips.rocketchip.system.DefaultRV32Config.fir@23633.4]
  wire  _GEN_73; // @[UserYanker.scala 69:36:freechips.rocketchip.system.DefaultRV32Config.fir@23633.4]
  wire  _GEN_74; // @[UserYanker.scala 69:36:freechips.rocketchip.system.DefaultRV32Config.fir@23633.4]
  wire  _GEN_75; // @[UserYanker.scala 69:36:freechips.rocketchip.system.DefaultRV32Config.fir@23633.4]
  wire  _GEN_76; // @[UserYanker.scala 69:36:freechips.rocketchip.system.DefaultRV32Config.fir@23633.4]
  wire  _GEN_77; // @[UserYanker.scala 69:36:freechips.rocketchip.system.DefaultRV32Config.fir@23633.4]
  wire  _GEN_78; // @[UserYanker.scala 69:36:freechips.rocketchip.system.DefaultRV32Config.fir@23633.4]
  wire  _GEN_79; // @[UserYanker.scala 69:36:freechips.rocketchip.system.DefaultRV32Config.fir@23633.4]
  wire  _T_157; // @[UserYanker.scala 76:15:freechips.rocketchip.system.DefaultRV32Config.fir@23682.4]
  wire  _T_155_0; // @[UserYanker.scala 74:24:freechips.rocketchip.system.DefaultRV32Config.fir@23646.4 UserYanker.scala 74:24:freechips.rocketchip.system.DefaultRV32Config.fir@23648.4]
  wire  _T_155_1; // @[UserYanker.scala 74:24:freechips.rocketchip.system.DefaultRV32Config.fir@23646.4 UserYanker.scala 74:24:freechips.rocketchip.system.DefaultRV32Config.fir@23649.4]
  wire  _GEN_81; // @[UserYanker.scala 76:28:freechips.rocketchip.system.DefaultRV32Config.fir@23683.4]
  wire  _T_155_2; // @[UserYanker.scala 74:24:freechips.rocketchip.system.DefaultRV32Config.fir@23646.4 UserYanker.scala 74:24:freechips.rocketchip.system.DefaultRV32Config.fir@23650.4]
  wire  _GEN_82; // @[UserYanker.scala 76:28:freechips.rocketchip.system.DefaultRV32Config.fir@23683.4]
  wire  _T_155_3; // @[UserYanker.scala 74:24:freechips.rocketchip.system.DefaultRV32Config.fir@23646.4 UserYanker.scala 74:24:freechips.rocketchip.system.DefaultRV32Config.fir@23651.4]
  wire  _GEN_83; // @[UserYanker.scala 76:28:freechips.rocketchip.system.DefaultRV32Config.fir@23683.4]
  wire  _T_155_4; // @[UserYanker.scala 74:24:freechips.rocketchip.system.DefaultRV32Config.fir@23646.4 UserYanker.scala 74:24:freechips.rocketchip.system.DefaultRV32Config.fir@23652.4]
  wire  _GEN_84; // @[UserYanker.scala 76:28:freechips.rocketchip.system.DefaultRV32Config.fir@23683.4]
  wire  _GEN_85; // @[UserYanker.scala 76:28:freechips.rocketchip.system.DefaultRV32Config.fir@23683.4]
  wire  _GEN_86; // @[UserYanker.scala 76:28:freechips.rocketchip.system.DefaultRV32Config.fir@23683.4]
  wire  _GEN_87; // @[UserYanker.scala 76:28:freechips.rocketchip.system.DefaultRV32Config.fir@23683.4]
  wire  _GEN_88; // @[UserYanker.scala 76:28:freechips.rocketchip.system.DefaultRV32Config.fir@23683.4]
  wire  _GEN_89; // @[UserYanker.scala 76:28:freechips.rocketchip.system.DefaultRV32Config.fir@23683.4]
  wire  _GEN_90; // @[UserYanker.scala 76:28:freechips.rocketchip.system.DefaultRV32Config.fir@23683.4]
  wire  _GEN_91; // @[UserYanker.scala 76:28:freechips.rocketchip.system.DefaultRV32Config.fir@23683.4]
  wire  _GEN_92; // @[UserYanker.scala 76:28:freechips.rocketchip.system.DefaultRV32Config.fir@23683.4]
  wire  _GEN_93; // @[UserYanker.scala 76:28:freechips.rocketchip.system.DefaultRV32Config.fir@23683.4]
  wire  _GEN_94; // @[UserYanker.scala 76:28:freechips.rocketchip.system.DefaultRV32Config.fir@23683.4]
  wire  _GEN_95; // @[UserYanker.scala 76:28:freechips.rocketchip.system.DefaultRV32Config.fir@23683.4]
  wire  _T_158; // @[UserYanker.scala 76:28:freechips.rocketchip.system.DefaultRV32Config.fir@23683.4]
  wire  _T_160; // @[UserYanker.scala 76:14:freechips.rocketchip.system.DefaultRV32Config.fir@23685.4]
  wire  _T_161; // @[UserYanker.scala 76:14:freechips.rocketchip.system.DefaultRV32Config.fir@23686.4]
  wire [3:0] _T_156_0_tl_state_size; // @[UserYanker.scala 75:23:freechips.rocketchip.system.DefaultRV32Config.fir@23664.4 UserYanker.scala 75:23:freechips.rocketchip.system.DefaultRV32Config.fir@23666.4]
  wire [4:0] _T_156_0_tl_state_source; // @[UserYanker.scala 75:23:freechips.rocketchip.system.DefaultRV32Config.fir@23664.4 UserYanker.scala 75:23:freechips.rocketchip.system.DefaultRV32Config.fir@23666.4]
  wire [3:0] _T_156_1_tl_state_size; // @[UserYanker.scala 75:23:freechips.rocketchip.system.DefaultRV32Config.fir@23664.4 UserYanker.scala 75:23:freechips.rocketchip.system.DefaultRV32Config.fir@23667.4]
  wire [3:0] _GEN_98; // @[BundleMap.scala 248:19:freechips.rocketchip.system.DefaultRV32Config.fir@23697.4]
  wire [4:0] _T_156_1_tl_state_source; // @[UserYanker.scala 75:23:freechips.rocketchip.system.DefaultRV32Config.fir@23664.4 UserYanker.scala 75:23:freechips.rocketchip.system.DefaultRV32Config.fir@23667.4]
  wire [4:0] _GEN_99; // @[BundleMap.scala 248:19:freechips.rocketchip.system.DefaultRV32Config.fir@23697.4]
  wire [3:0] _T_156_2_tl_state_size; // @[UserYanker.scala 75:23:freechips.rocketchip.system.DefaultRV32Config.fir@23664.4 UserYanker.scala 75:23:freechips.rocketchip.system.DefaultRV32Config.fir@23668.4]
  wire [3:0] _GEN_100; // @[BundleMap.scala 248:19:freechips.rocketchip.system.DefaultRV32Config.fir@23697.4]
  wire [4:0] _T_156_2_tl_state_source; // @[UserYanker.scala 75:23:freechips.rocketchip.system.DefaultRV32Config.fir@23664.4 UserYanker.scala 75:23:freechips.rocketchip.system.DefaultRV32Config.fir@23668.4]
  wire [4:0] _GEN_101; // @[BundleMap.scala 248:19:freechips.rocketchip.system.DefaultRV32Config.fir@23697.4]
  wire [3:0] _T_156_3_tl_state_size; // @[UserYanker.scala 75:23:freechips.rocketchip.system.DefaultRV32Config.fir@23664.4 UserYanker.scala 75:23:freechips.rocketchip.system.DefaultRV32Config.fir@23669.4]
  wire [3:0] _GEN_102; // @[BundleMap.scala 248:19:freechips.rocketchip.system.DefaultRV32Config.fir@23697.4]
  wire [4:0] _T_156_3_tl_state_source; // @[UserYanker.scala 75:23:freechips.rocketchip.system.DefaultRV32Config.fir@23664.4 UserYanker.scala 75:23:freechips.rocketchip.system.DefaultRV32Config.fir@23669.4]
  wire [4:0] _GEN_103; // @[BundleMap.scala 248:19:freechips.rocketchip.system.DefaultRV32Config.fir@23697.4]
  wire [3:0] _T_156_4_tl_state_size; // @[UserYanker.scala 75:23:freechips.rocketchip.system.DefaultRV32Config.fir@23664.4 UserYanker.scala 75:23:freechips.rocketchip.system.DefaultRV32Config.fir@23670.4]
  wire [3:0] _GEN_104; // @[BundleMap.scala 248:19:freechips.rocketchip.system.DefaultRV32Config.fir@23697.4]
  wire [4:0] _T_156_4_tl_state_source; // @[UserYanker.scala 75:23:freechips.rocketchip.system.DefaultRV32Config.fir@23664.4 UserYanker.scala 75:23:freechips.rocketchip.system.DefaultRV32Config.fir@23670.4]
  wire [4:0] _GEN_105; // @[BundleMap.scala 248:19:freechips.rocketchip.system.DefaultRV32Config.fir@23697.4]
  wire [3:0] _GEN_106; // @[BundleMap.scala 248:19:freechips.rocketchip.system.DefaultRV32Config.fir@23697.4]
  wire [4:0] _GEN_107; // @[BundleMap.scala 248:19:freechips.rocketchip.system.DefaultRV32Config.fir@23697.4]
  wire [3:0] _GEN_108; // @[BundleMap.scala 248:19:freechips.rocketchip.system.DefaultRV32Config.fir@23697.4]
  wire [4:0] _GEN_109; // @[BundleMap.scala 248:19:freechips.rocketchip.system.DefaultRV32Config.fir@23697.4]
  wire [3:0] _GEN_110; // @[BundleMap.scala 248:19:freechips.rocketchip.system.DefaultRV32Config.fir@23697.4]
  wire [4:0] _GEN_111; // @[BundleMap.scala 248:19:freechips.rocketchip.system.DefaultRV32Config.fir@23697.4]
  wire [3:0] _GEN_112; // @[BundleMap.scala 248:19:freechips.rocketchip.system.DefaultRV32Config.fir@23697.4]
  wire [4:0] _GEN_113; // @[BundleMap.scala 248:19:freechips.rocketchip.system.DefaultRV32Config.fir@23697.4]
  wire [3:0] _GEN_114; // @[BundleMap.scala 248:19:freechips.rocketchip.system.DefaultRV32Config.fir@23697.4]
  wire [4:0] _GEN_115; // @[BundleMap.scala 248:19:freechips.rocketchip.system.DefaultRV32Config.fir@23697.4]
  wire [3:0] _GEN_116; // @[BundleMap.scala 248:19:freechips.rocketchip.system.DefaultRV32Config.fir@23697.4]
  wire [4:0] _GEN_117; // @[BundleMap.scala 248:19:freechips.rocketchip.system.DefaultRV32Config.fir@23697.4]
  wire [3:0] _GEN_118; // @[BundleMap.scala 248:19:freechips.rocketchip.system.DefaultRV32Config.fir@23697.4]
  wire [4:0] _GEN_119; // @[BundleMap.scala 248:19:freechips.rocketchip.system.DefaultRV32Config.fir@23697.4]
  wire [3:0] _GEN_120; // @[BundleMap.scala 248:19:freechips.rocketchip.system.DefaultRV32Config.fir@23697.4]
  wire [4:0] _GEN_121; // @[BundleMap.scala 248:19:freechips.rocketchip.system.DefaultRV32Config.fir@23697.4]
  wire [3:0] _GEN_122; // @[BundleMap.scala 248:19:freechips.rocketchip.system.DefaultRV32Config.fir@23697.4]
  wire [4:0] _GEN_123; // @[BundleMap.scala 248:19:freechips.rocketchip.system.DefaultRV32Config.fir@23697.4]
  wire [3:0] _GEN_124; // @[BundleMap.scala 248:19:freechips.rocketchip.system.DefaultRV32Config.fir@23697.4]
  wire [4:0] _GEN_125; // @[BundleMap.scala 248:19:freechips.rocketchip.system.DefaultRV32Config.fir@23697.4]
  wire [15:0] _T_163; // @[OneHot.scala 65:12:freechips.rocketchip.system.DefaultRV32Config.fir@23700.4]
  wire [15:0] _T_182; // @[OneHot.scala 65:12:freechips.rocketchip.system.DefaultRV32Config.fir@23719.4]
  wire  _T_200; // @[UserYanker.scala 83:37:freechips.rocketchip.system.DefaultRV32Config.fir@23737.4]
  wire  _T_202; // @[UserYanker.scala 84:37:freechips.rocketchip.system.DefaultRV32Config.fir@23740.4]
  QueueCompatibility QueueCompatibility ( // @[UserYanker.scala 39:17:freechips.rocketchip.system.DefaultRV32Config.fir@23263.4]
    .clock(QueueCompatibility_clock),
    .reset(QueueCompatibility_reset),
    .io_enq_ready(QueueCompatibility_io_enq_ready),
    .io_enq_valid(QueueCompatibility_io_enq_valid),
    .io_enq_bits_tl_state_size(QueueCompatibility_io_enq_bits_tl_state_size),
    .io_enq_bits_tl_state_source(QueueCompatibility_io_enq_bits_tl_state_source),
    .io_deq_ready(QueueCompatibility_io_deq_ready),
    .io_deq_valid(QueueCompatibility_io_deq_valid),
    .io_deq_bits_tl_state_size(QueueCompatibility_io_deq_bits_tl_state_size),
    .io_deq_bits_tl_state_source(QueueCompatibility_io_deq_bits_tl_state_source)
  );
  QueueCompatibility_1 QueueCompatibility_1 ( // @[UserYanker.scala 39:17:freechips.rocketchip.system.DefaultRV32Config.fir@23267.4]
    .clock(QueueCompatibility_1_clock),
    .reset(QueueCompatibility_1_reset),
    .io_enq_ready(QueueCompatibility_1_io_enq_ready),
    .io_enq_valid(QueueCompatibility_1_io_enq_valid),
    .io_enq_bits_tl_state_size(QueueCompatibility_1_io_enq_bits_tl_state_size),
    .io_enq_bits_tl_state_source(QueueCompatibility_1_io_enq_bits_tl_state_source),
    .io_deq_ready(QueueCompatibility_1_io_deq_ready),
    .io_deq_valid(QueueCompatibility_1_io_deq_valid),
    .io_deq_bits_tl_state_size(QueueCompatibility_1_io_deq_bits_tl_state_size),
    .io_deq_bits_tl_state_source(QueueCompatibility_1_io_deq_bits_tl_state_source)
  );
  QueueCompatibility_1 QueueCompatibility_2 ( // @[UserYanker.scala 39:17:freechips.rocketchip.system.DefaultRV32Config.fir@23271.4]
    .clock(QueueCompatibility_2_clock),
    .reset(QueueCompatibility_2_reset),
    .io_enq_ready(QueueCompatibility_2_io_enq_ready),
    .io_enq_valid(QueueCompatibility_2_io_enq_valid),
    .io_enq_bits_tl_state_size(QueueCompatibility_2_io_enq_bits_tl_state_size),
    .io_enq_bits_tl_state_source(QueueCompatibility_2_io_enq_bits_tl_state_source),
    .io_deq_ready(QueueCompatibility_2_io_deq_ready),
    .io_deq_valid(QueueCompatibility_2_io_deq_valid),
    .io_deq_bits_tl_state_size(QueueCompatibility_2_io_deq_bits_tl_state_size),
    .io_deq_bits_tl_state_source(QueueCompatibility_2_io_deq_bits_tl_state_source)
  );
  QueueCompatibility QueueCompatibility_3 ( // @[UserYanker.scala 39:17:freechips.rocketchip.system.DefaultRV32Config.fir@23275.4]
    .clock(QueueCompatibility_3_clock),
    .reset(QueueCompatibility_3_reset),
    .io_enq_ready(QueueCompatibility_3_io_enq_ready),
    .io_enq_valid(QueueCompatibility_3_io_enq_valid),
    .io_enq_bits_tl_state_size(QueueCompatibility_3_io_enq_bits_tl_state_size),
    .io_enq_bits_tl_state_source(QueueCompatibility_3_io_enq_bits_tl_state_source),
    .io_deq_ready(QueueCompatibility_3_io_deq_ready),
    .io_deq_valid(QueueCompatibility_3_io_deq_valid),
    .io_deq_bits_tl_state_size(QueueCompatibility_3_io_deq_bits_tl_state_size),
    .io_deq_bits_tl_state_source(QueueCompatibility_3_io_deq_bits_tl_state_source)
  );
  QueueCompatibility QueueCompatibility_4 ( // @[UserYanker.scala 39:17:freechips.rocketchip.system.DefaultRV32Config.fir@23279.4]
    .clock(QueueCompatibility_4_clock),
    .reset(QueueCompatibility_4_reset),
    .io_enq_ready(QueueCompatibility_4_io_enq_ready),
    .io_enq_valid(QueueCompatibility_4_io_enq_valid),
    .io_enq_bits_tl_state_size(QueueCompatibility_4_io_enq_bits_tl_state_size),
    .io_enq_bits_tl_state_source(QueueCompatibility_4_io_enq_bits_tl_state_source),
    .io_deq_ready(QueueCompatibility_4_io_deq_ready),
    .io_deq_valid(QueueCompatibility_4_io_deq_valid),
    .io_deq_bits_tl_state_size(QueueCompatibility_4_io_deq_bits_tl_state_size),
    .io_deq_bits_tl_state_source(QueueCompatibility_4_io_deq_bits_tl_state_source)
  );
  QueueCompatibility QueueCompatibility_5 ( // @[UserYanker.scala 39:17:freechips.rocketchip.system.DefaultRV32Config.fir@23305.4]
    .clock(QueueCompatibility_5_clock),
    .reset(QueueCompatibility_5_reset),
    .io_enq_ready(QueueCompatibility_5_io_enq_ready),
    .io_enq_valid(QueueCompatibility_5_io_enq_valid),
    .io_enq_bits_tl_state_size(QueueCompatibility_5_io_enq_bits_tl_state_size),
    .io_enq_bits_tl_state_source(QueueCompatibility_5_io_enq_bits_tl_state_source),
    .io_deq_ready(QueueCompatibility_5_io_deq_ready),
    .io_deq_valid(QueueCompatibility_5_io_deq_valid),
    .io_deq_bits_tl_state_size(QueueCompatibility_5_io_deq_bits_tl_state_size),
    .io_deq_bits_tl_state_source(QueueCompatibility_5_io_deq_bits_tl_state_source)
  );
  QueueCompatibility_1 QueueCompatibility_6 ( // @[UserYanker.scala 39:17:freechips.rocketchip.system.DefaultRV32Config.fir@23309.4]
    .clock(QueueCompatibility_6_clock),
    .reset(QueueCompatibility_6_reset),
    .io_enq_ready(QueueCompatibility_6_io_enq_ready),
    .io_enq_valid(QueueCompatibility_6_io_enq_valid),
    .io_enq_bits_tl_state_size(QueueCompatibility_6_io_enq_bits_tl_state_size),
    .io_enq_bits_tl_state_source(QueueCompatibility_6_io_enq_bits_tl_state_source),
    .io_deq_ready(QueueCompatibility_6_io_deq_ready),
    .io_deq_valid(QueueCompatibility_6_io_deq_valid),
    .io_deq_bits_tl_state_size(QueueCompatibility_6_io_deq_bits_tl_state_size),
    .io_deq_bits_tl_state_source(QueueCompatibility_6_io_deq_bits_tl_state_source)
  );
  QueueCompatibility_1 QueueCompatibility_7 ( // @[UserYanker.scala 39:17:freechips.rocketchip.system.DefaultRV32Config.fir@23313.4]
    .clock(QueueCompatibility_7_clock),
    .reset(QueueCompatibility_7_reset),
    .io_enq_ready(QueueCompatibility_7_io_enq_ready),
    .io_enq_valid(QueueCompatibility_7_io_enq_valid),
    .io_enq_bits_tl_state_size(QueueCompatibility_7_io_enq_bits_tl_state_size),
    .io_enq_bits_tl_state_source(QueueCompatibility_7_io_enq_bits_tl_state_source),
    .io_deq_ready(QueueCompatibility_7_io_deq_ready),
    .io_deq_valid(QueueCompatibility_7_io_deq_valid),
    .io_deq_bits_tl_state_size(QueueCompatibility_7_io_deq_bits_tl_state_size),
    .io_deq_bits_tl_state_source(QueueCompatibility_7_io_deq_bits_tl_state_source)
  );
  QueueCompatibility QueueCompatibility_8 ( // @[UserYanker.scala 39:17:freechips.rocketchip.system.DefaultRV32Config.fir@23317.4]
    .clock(QueueCompatibility_8_clock),
    .reset(QueueCompatibility_8_reset),
    .io_enq_ready(QueueCompatibility_8_io_enq_ready),
    .io_enq_valid(QueueCompatibility_8_io_enq_valid),
    .io_enq_bits_tl_state_size(QueueCompatibility_8_io_enq_bits_tl_state_size),
    .io_enq_bits_tl_state_source(QueueCompatibility_8_io_enq_bits_tl_state_source),
    .io_deq_ready(QueueCompatibility_8_io_deq_ready),
    .io_deq_valid(QueueCompatibility_8_io_deq_valid),
    .io_deq_bits_tl_state_size(QueueCompatibility_8_io_deq_bits_tl_state_size),
    .io_deq_bits_tl_state_source(QueueCompatibility_8_io_deq_bits_tl_state_source)
  );
  QueueCompatibility QueueCompatibility_9 ( // @[UserYanker.scala 39:17:freechips.rocketchip.system.DefaultRV32Config.fir@23321.4]
    .clock(QueueCompatibility_9_clock),
    .reset(QueueCompatibility_9_reset),
    .io_enq_ready(QueueCompatibility_9_io_enq_ready),
    .io_enq_valid(QueueCompatibility_9_io_enq_valid),
    .io_enq_bits_tl_state_size(QueueCompatibility_9_io_enq_bits_tl_state_size),
    .io_enq_bits_tl_state_source(QueueCompatibility_9_io_enq_bits_tl_state_source),
    .io_deq_ready(QueueCompatibility_9_io_deq_ready),
    .io_deq_valid(QueueCompatibility_9_io_deq_valid),
    .io_deq_bits_tl_state_size(QueueCompatibility_9_io_deq_bits_tl_state_size),
    .io_deq_bits_tl_state_source(QueueCompatibility_9_io_deq_bits_tl_state_source)
  );
  assign _T_24_0 = QueueCompatibility_io_enq_ready; // @[UserYanker.scala 47:25:freechips.rocketchip.system.DefaultRV32Config.fir@23347.4 UserYanker.scala 47:25:freechips.rocketchip.system.DefaultRV32Config.fir@23349.4]
  assign _T_24_1 = QueueCompatibility_1_io_enq_ready; // @[UserYanker.scala 47:25:freechips.rocketchip.system.DefaultRV32Config.fir@23347.4 UserYanker.scala 47:25:freechips.rocketchip.system.DefaultRV32Config.fir@23350.4]
  assign _GEN_1 = 4'h1 == auto_in_ar_bits_id ? _T_24_1 : _T_24_0; // @[UserYanker.scala 48:36:freechips.rocketchip.system.DefaultRV32Config.fir@23365.4]
  assign _T_24_2 = QueueCompatibility_2_io_enq_ready; // @[UserYanker.scala 47:25:freechips.rocketchip.system.DefaultRV32Config.fir@23347.4 UserYanker.scala 47:25:freechips.rocketchip.system.DefaultRV32Config.fir@23351.4]
  assign _GEN_2 = 4'h2 == auto_in_ar_bits_id ? _T_24_2 : _GEN_1; // @[UserYanker.scala 48:36:freechips.rocketchip.system.DefaultRV32Config.fir@23365.4]
  assign _T_24_3 = QueueCompatibility_3_io_enq_ready; // @[UserYanker.scala 47:25:freechips.rocketchip.system.DefaultRV32Config.fir@23347.4 UserYanker.scala 47:25:freechips.rocketchip.system.DefaultRV32Config.fir@23352.4]
  assign _GEN_3 = 4'h3 == auto_in_ar_bits_id ? _T_24_3 : _GEN_2; // @[UserYanker.scala 48:36:freechips.rocketchip.system.DefaultRV32Config.fir@23365.4]
  assign _T_24_4 = QueueCompatibility_4_io_enq_ready; // @[UserYanker.scala 47:25:freechips.rocketchip.system.DefaultRV32Config.fir@23347.4 UserYanker.scala 47:25:freechips.rocketchip.system.DefaultRV32Config.fir@23353.4]
  assign _GEN_4 = 4'h4 == auto_in_ar_bits_id ? _T_24_4 : _GEN_3; // @[UserYanker.scala 48:36:freechips.rocketchip.system.DefaultRV32Config.fir@23365.4]
  assign _GEN_5 = 4'h5 == auto_in_ar_bits_id ? 1'h0 : _GEN_4; // @[UserYanker.scala 48:36:freechips.rocketchip.system.DefaultRV32Config.fir@23365.4]
  assign _GEN_6 = 4'h6 == auto_in_ar_bits_id ? 1'h0 : _GEN_5; // @[UserYanker.scala 48:36:freechips.rocketchip.system.DefaultRV32Config.fir@23365.4]
  assign _GEN_7 = 4'h7 == auto_in_ar_bits_id ? 1'h0 : _GEN_6; // @[UserYanker.scala 48:36:freechips.rocketchip.system.DefaultRV32Config.fir@23365.4]
  assign _GEN_8 = 4'h8 == auto_in_ar_bits_id ? 1'h0 : _GEN_7; // @[UserYanker.scala 48:36:freechips.rocketchip.system.DefaultRV32Config.fir@23365.4]
  assign _GEN_9 = 4'h9 == auto_in_ar_bits_id ? 1'h0 : _GEN_8; // @[UserYanker.scala 48:36:freechips.rocketchip.system.DefaultRV32Config.fir@23365.4]
  assign _GEN_10 = 4'ha == auto_in_ar_bits_id ? 1'h0 : _GEN_9; // @[UserYanker.scala 48:36:freechips.rocketchip.system.DefaultRV32Config.fir@23365.4]
  assign _GEN_11 = 4'hb == auto_in_ar_bits_id ? 1'h0 : _GEN_10; // @[UserYanker.scala 48:36:freechips.rocketchip.system.DefaultRV32Config.fir@23365.4]
  assign _GEN_12 = 4'hc == auto_in_ar_bits_id ? 1'h0 : _GEN_11; // @[UserYanker.scala 48:36:freechips.rocketchip.system.DefaultRV32Config.fir@23365.4]
  assign _GEN_13 = 4'hd == auto_in_ar_bits_id ? 1'h0 : _GEN_12; // @[UserYanker.scala 48:36:freechips.rocketchip.system.DefaultRV32Config.fir@23365.4]
  assign _GEN_14 = 4'he == auto_in_ar_bits_id ? 1'h0 : _GEN_13; // @[UserYanker.scala 48:36:freechips.rocketchip.system.DefaultRV32Config.fir@23365.4]
  assign _GEN_15 = 4'hf == auto_in_ar_bits_id ? 1'h0 : _GEN_14; // @[UserYanker.scala 48:36:freechips.rocketchip.system.DefaultRV32Config.fir@23365.4]
  assign _T_29 = ~auto_out_r_valid; // @[UserYanker.scala 55:15:freechips.rocketchip.system.DefaultRV32Config.fir@23414.4]
  assign _T_27_0 = QueueCompatibility_io_deq_valid; // @[UserYanker.scala 53:24:freechips.rocketchip.system.DefaultRV32Config.fir@23378.4 UserYanker.scala 53:24:freechips.rocketchip.system.DefaultRV32Config.fir@23380.4]
  assign _T_27_1 = QueueCompatibility_1_io_deq_valid; // @[UserYanker.scala 53:24:freechips.rocketchip.system.DefaultRV32Config.fir@23378.4 UserYanker.scala 53:24:freechips.rocketchip.system.DefaultRV32Config.fir@23381.4]
  assign _GEN_17 = 4'h1 == auto_out_r_bits_id ? _T_27_1 : _T_27_0; // @[UserYanker.scala 55:28:freechips.rocketchip.system.DefaultRV32Config.fir@23415.4]
  assign _T_27_2 = QueueCompatibility_2_io_deq_valid; // @[UserYanker.scala 53:24:freechips.rocketchip.system.DefaultRV32Config.fir@23378.4 UserYanker.scala 53:24:freechips.rocketchip.system.DefaultRV32Config.fir@23382.4]
  assign _GEN_18 = 4'h2 == auto_out_r_bits_id ? _T_27_2 : _GEN_17; // @[UserYanker.scala 55:28:freechips.rocketchip.system.DefaultRV32Config.fir@23415.4]
  assign _T_27_3 = QueueCompatibility_3_io_deq_valid; // @[UserYanker.scala 53:24:freechips.rocketchip.system.DefaultRV32Config.fir@23378.4 UserYanker.scala 53:24:freechips.rocketchip.system.DefaultRV32Config.fir@23383.4]
  assign _GEN_19 = 4'h3 == auto_out_r_bits_id ? _T_27_3 : _GEN_18; // @[UserYanker.scala 55:28:freechips.rocketchip.system.DefaultRV32Config.fir@23415.4]
  assign _T_27_4 = QueueCompatibility_4_io_deq_valid; // @[UserYanker.scala 53:24:freechips.rocketchip.system.DefaultRV32Config.fir@23378.4 UserYanker.scala 53:24:freechips.rocketchip.system.DefaultRV32Config.fir@23384.4]
  assign _GEN_20 = 4'h4 == auto_out_r_bits_id ? _T_27_4 : _GEN_19; // @[UserYanker.scala 55:28:freechips.rocketchip.system.DefaultRV32Config.fir@23415.4]
  assign _GEN_21 = 4'h5 == auto_out_r_bits_id ? 1'h0 : _GEN_20; // @[UserYanker.scala 55:28:freechips.rocketchip.system.DefaultRV32Config.fir@23415.4]
  assign _GEN_22 = 4'h6 == auto_out_r_bits_id ? 1'h0 : _GEN_21; // @[UserYanker.scala 55:28:freechips.rocketchip.system.DefaultRV32Config.fir@23415.4]
  assign _GEN_23 = 4'h7 == auto_out_r_bits_id ? 1'h0 : _GEN_22; // @[UserYanker.scala 55:28:freechips.rocketchip.system.DefaultRV32Config.fir@23415.4]
  assign _GEN_24 = 4'h8 == auto_out_r_bits_id ? 1'h0 : _GEN_23; // @[UserYanker.scala 55:28:freechips.rocketchip.system.DefaultRV32Config.fir@23415.4]
  assign _GEN_25 = 4'h9 == auto_out_r_bits_id ? 1'h0 : _GEN_24; // @[UserYanker.scala 55:28:freechips.rocketchip.system.DefaultRV32Config.fir@23415.4]
  assign _GEN_26 = 4'ha == auto_out_r_bits_id ? 1'h0 : _GEN_25; // @[UserYanker.scala 55:28:freechips.rocketchip.system.DefaultRV32Config.fir@23415.4]
  assign _GEN_27 = 4'hb == auto_out_r_bits_id ? 1'h0 : _GEN_26; // @[UserYanker.scala 55:28:freechips.rocketchip.system.DefaultRV32Config.fir@23415.4]
  assign _GEN_28 = 4'hc == auto_out_r_bits_id ? 1'h0 : _GEN_27; // @[UserYanker.scala 55:28:freechips.rocketchip.system.DefaultRV32Config.fir@23415.4]
  assign _GEN_29 = 4'hd == auto_out_r_bits_id ? 1'h0 : _GEN_28; // @[UserYanker.scala 55:28:freechips.rocketchip.system.DefaultRV32Config.fir@23415.4]
  assign _GEN_30 = 4'he == auto_out_r_bits_id ? 1'h0 : _GEN_29; // @[UserYanker.scala 55:28:freechips.rocketchip.system.DefaultRV32Config.fir@23415.4]
  assign _GEN_31 = 4'hf == auto_out_r_bits_id ? 1'h0 : _GEN_30; // @[UserYanker.scala 55:28:freechips.rocketchip.system.DefaultRV32Config.fir@23415.4]
  assign _T_30 = _T_29 | _GEN_31; // @[UserYanker.scala 55:28:freechips.rocketchip.system.DefaultRV32Config.fir@23415.4]
  assign _T_32 = _T_30 | reset; // @[UserYanker.scala 55:14:freechips.rocketchip.system.DefaultRV32Config.fir@23417.4]
  assign _T_33 = ~_T_32; // @[UserYanker.scala 55:14:freechips.rocketchip.system.DefaultRV32Config.fir@23418.4]
  assign _T_28_0_tl_state_size = QueueCompatibility_io_deq_bits_tl_state_size; // @[UserYanker.scala 54:23:freechips.rocketchip.system.DefaultRV32Config.fir@23396.4 UserYanker.scala 54:23:freechips.rocketchip.system.DefaultRV32Config.fir@23398.4]
  assign _T_28_0_tl_state_source = QueueCompatibility_io_deq_bits_tl_state_source; // @[UserYanker.scala 54:23:freechips.rocketchip.system.DefaultRV32Config.fir@23396.4 UserYanker.scala 54:23:freechips.rocketchip.system.DefaultRV32Config.fir@23398.4]
  assign _T_28_1_tl_state_size = QueueCompatibility_1_io_deq_bits_tl_state_size; // @[UserYanker.scala 54:23:freechips.rocketchip.system.DefaultRV32Config.fir@23396.4 UserYanker.scala 54:23:freechips.rocketchip.system.DefaultRV32Config.fir@23399.4]
  assign _GEN_34 = 4'h1 == auto_out_r_bits_id ? _T_28_1_tl_state_size : _T_28_0_tl_state_size; // @[BundleMap.scala 248:19:freechips.rocketchip.system.DefaultRV32Config.fir@23431.4]
  assign _T_28_1_tl_state_source = QueueCompatibility_1_io_deq_bits_tl_state_source; // @[UserYanker.scala 54:23:freechips.rocketchip.system.DefaultRV32Config.fir@23396.4 UserYanker.scala 54:23:freechips.rocketchip.system.DefaultRV32Config.fir@23399.4]
  assign _GEN_35 = 4'h1 == auto_out_r_bits_id ? _T_28_1_tl_state_source : _T_28_0_tl_state_source; // @[BundleMap.scala 248:19:freechips.rocketchip.system.DefaultRV32Config.fir@23431.4]
  assign _T_28_2_tl_state_size = QueueCompatibility_2_io_deq_bits_tl_state_size; // @[UserYanker.scala 54:23:freechips.rocketchip.system.DefaultRV32Config.fir@23396.4 UserYanker.scala 54:23:freechips.rocketchip.system.DefaultRV32Config.fir@23400.4]
  assign _GEN_36 = 4'h2 == auto_out_r_bits_id ? _T_28_2_tl_state_size : _GEN_34; // @[BundleMap.scala 248:19:freechips.rocketchip.system.DefaultRV32Config.fir@23431.4]
  assign _T_28_2_tl_state_source = QueueCompatibility_2_io_deq_bits_tl_state_source; // @[UserYanker.scala 54:23:freechips.rocketchip.system.DefaultRV32Config.fir@23396.4 UserYanker.scala 54:23:freechips.rocketchip.system.DefaultRV32Config.fir@23400.4]
  assign _GEN_37 = 4'h2 == auto_out_r_bits_id ? _T_28_2_tl_state_source : _GEN_35; // @[BundleMap.scala 248:19:freechips.rocketchip.system.DefaultRV32Config.fir@23431.4]
  assign _T_28_3_tl_state_size = QueueCompatibility_3_io_deq_bits_tl_state_size; // @[UserYanker.scala 54:23:freechips.rocketchip.system.DefaultRV32Config.fir@23396.4 UserYanker.scala 54:23:freechips.rocketchip.system.DefaultRV32Config.fir@23401.4]
  assign _GEN_38 = 4'h3 == auto_out_r_bits_id ? _T_28_3_tl_state_size : _GEN_36; // @[BundleMap.scala 248:19:freechips.rocketchip.system.DefaultRV32Config.fir@23431.4]
  assign _T_28_3_tl_state_source = QueueCompatibility_3_io_deq_bits_tl_state_source; // @[UserYanker.scala 54:23:freechips.rocketchip.system.DefaultRV32Config.fir@23396.4 UserYanker.scala 54:23:freechips.rocketchip.system.DefaultRV32Config.fir@23401.4]
  assign _GEN_39 = 4'h3 == auto_out_r_bits_id ? _T_28_3_tl_state_source : _GEN_37; // @[BundleMap.scala 248:19:freechips.rocketchip.system.DefaultRV32Config.fir@23431.4]
  assign _T_28_4_tl_state_size = QueueCompatibility_4_io_deq_bits_tl_state_size; // @[UserYanker.scala 54:23:freechips.rocketchip.system.DefaultRV32Config.fir@23396.4 UserYanker.scala 54:23:freechips.rocketchip.system.DefaultRV32Config.fir@23402.4]
  assign _GEN_40 = 4'h4 == auto_out_r_bits_id ? _T_28_4_tl_state_size : _GEN_38; // @[BundleMap.scala 248:19:freechips.rocketchip.system.DefaultRV32Config.fir@23431.4]
  assign _T_28_4_tl_state_source = QueueCompatibility_4_io_deq_bits_tl_state_source; // @[UserYanker.scala 54:23:freechips.rocketchip.system.DefaultRV32Config.fir@23396.4 UserYanker.scala 54:23:freechips.rocketchip.system.DefaultRV32Config.fir@23402.4]
  assign _GEN_41 = 4'h4 == auto_out_r_bits_id ? _T_28_4_tl_state_source : _GEN_39; // @[BundleMap.scala 248:19:freechips.rocketchip.system.DefaultRV32Config.fir@23431.4]
  assign _GEN_42 = 4'h5 == auto_out_r_bits_id ? 4'h0 : _GEN_40; // @[BundleMap.scala 248:19:freechips.rocketchip.system.DefaultRV32Config.fir@23431.4]
  assign _GEN_43 = 4'h5 == auto_out_r_bits_id ? 5'h0 : _GEN_41; // @[BundleMap.scala 248:19:freechips.rocketchip.system.DefaultRV32Config.fir@23431.4]
  assign _GEN_44 = 4'h6 == auto_out_r_bits_id ? 4'h0 : _GEN_42; // @[BundleMap.scala 248:19:freechips.rocketchip.system.DefaultRV32Config.fir@23431.4]
  assign _GEN_45 = 4'h6 == auto_out_r_bits_id ? 5'h0 : _GEN_43; // @[BundleMap.scala 248:19:freechips.rocketchip.system.DefaultRV32Config.fir@23431.4]
  assign _GEN_46 = 4'h7 == auto_out_r_bits_id ? 4'h0 : _GEN_44; // @[BundleMap.scala 248:19:freechips.rocketchip.system.DefaultRV32Config.fir@23431.4]
  assign _GEN_47 = 4'h7 == auto_out_r_bits_id ? 5'h0 : _GEN_45; // @[BundleMap.scala 248:19:freechips.rocketchip.system.DefaultRV32Config.fir@23431.4]
  assign _GEN_48 = 4'h8 == auto_out_r_bits_id ? 4'h0 : _GEN_46; // @[BundleMap.scala 248:19:freechips.rocketchip.system.DefaultRV32Config.fir@23431.4]
  assign _GEN_49 = 4'h8 == auto_out_r_bits_id ? 5'h0 : _GEN_47; // @[BundleMap.scala 248:19:freechips.rocketchip.system.DefaultRV32Config.fir@23431.4]
  assign _GEN_50 = 4'h9 == auto_out_r_bits_id ? 4'h0 : _GEN_48; // @[BundleMap.scala 248:19:freechips.rocketchip.system.DefaultRV32Config.fir@23431.4]
  assign _GEN_51 = 4'h9 == auto_out_r_bits_id ? 5'h0 : _GEN_49; // @[BundleMap.scala 248:19:freechips.rocketchip.system.DefaultRV32Config.fir@23431.4]
  assign _GEN_52 = 4'ha == auto_out_r_bits_id ? 4'h0 : _GEN_50; // @[BundleMap.scala 248:19:freechips.rocketchip.system.DefaultRV32Config.fir@23431.4]
  assign _GEN_53 = 4'ha == auto_out_r_bits_id ? 5'h0 : _GEN_51; // @[BundleMap.scala 248:19:freechips.rocketchip.system.DefaultRV32Config.fir@23431.4]
  assign _GEN_54 = 4'hb == auto_out_r_bits_id ? 4'h0 : _GEN_52; // @[BundleMap.scala 248:19:freechips.rocketchip.system.DefaultRV32Config.fir@23431.4]
  assign _GEN_55 = 4'hb == auto_out_r_bits_id ? 5'h0 : _GEN_53; // @[BundleMap.scala 248:19:freechips.rocketchip.system.DefaultRV32Config.fir@23431.4]
  assign _GEN_56 = 4'hc == auto_out_r_bits_id ? 4'h0 : _GEN_54; // @[BundleMap.scala 248:19:freechips.rocketchip.system.DefaultRV32Config.fir@23431.4]
  assign _GEN_57 = 4'hc == auto_out_r_bits_id ? 5'h0 : _GEN_55; // @[BundleMap.scala 248:19:freechips.rocketchip.system.DefaultRV32Config.fir@23431.4]
  assign _GEN_58 = 4'hd == auto_out_r_bits_id ? 4'h0 : _GEN_56; // @[BundleMap.scala 248:19:freechips.rocketchip.system.DefaultRV32Config.fir@23431.4]
  assign _GEN_59 = 4'hd == auto_out_r_bits_id ? 5'h0 : _GEN_57; // @[BundleMap.scala 248:19:freechips.rocketchip.system.DefaultRV32Config.fir@23431.4]
  assign _GEN_60 = 4'he == auto_out_r_bits_id ? 4'h0 : _GEN_58; // @[BundleMap.scala 248:19:freechips.rocketchip.system.DefaultRV32Config.fir@23431.4]
  assign _GEN_61 = 4'he == auto_out_r_bits_id ? 5'h0 : _GEN_59; // @[BundleMap.scala 248:19:freechips.rocketchip.system.DefaultRV32Config.fir@23431.4]
  assign _T_35 = 16'h1 << auto_in_ar_bits_id; // @[OneHot.scala 65:12:freechips.rocketchip.system.DefaultRV32Config.fir@23434.4]
  assign _T_54 = 16'h1 << auto_out_r_bits_id; // @[OneHot.scala 65:12:freechips.rocketchip.system.DefaultRV32Config.fir@23453.4]
  assign _T_72 = auto_out_r_valid & auto_in_r_ready; // @[UserYanker.scala 62:37:freechips.rocketchip.system.DefaultRV32Config.fir@23471.4]
  assign _T_73 = _T_72 & _T_54[0]; // @[UserYanker.scala 62:53:freechips.rocketchip.system.DefaultRV32Config.fir@23472.4]
  assign _T_75 = auto_in_ar_valid & auto_out_ar_ready; // @[UserYanker.scala 63:37:freechips.rocketchip.system.DefaultRV32Config.fir@23475.4]
  assign _T_78 = _T_72 & _T_54[1]; // @[UserYanker.scala 62:53:freechips.rocketchip.system.DefaultRV32Config.fir@23481.4]
  assign _T_83 = _T_72 & _T_54[2]; // @[UserYanker.scala 62:53:freechips.rocketchip.system.DefaultRV32Config.fir@23490.4]
  assign _T_88 = _T_72 & _T_54[3]; // @[UserYanker.scala 62:53:freechips.rocketchip.system.DefaultRV32Config.fir@23499.4]
  assign _T_93 = _T_72 & _T_54[4]; // @[UserYanker.scala 62:53:freechips.rocketchip.system.DefaultRV32Config.fir@23508.4]
  assign _T_152_0 = QueueCompatibility_5_io_enq_ready; // @[UserYanker.scala 68:25:freechips.rocketchip.system.DefaultRV32Config.fir@23615.4 UserYanker.scala 68:25:freechips.rocketchip.system.DefaultRV32Config.fir@23617.4]
  assign _T_152_1 = QueueCompatibility_6_io_enq_ready; // @[UserYanker.scala 68:25:freechips.rocketchip.system.DefaultRV32Config.fir@23615.4 UserYanker.scala 68:25:freechips.rocketchip.system.DefaultRV32Config.fir@23618.4]
  assign _GEN_65 = 4'h1 == auto_in_aw_bits_id ? _T_152_1 : _T_152_0; // @[UserYanker.scala 69:36:freechips.rocketchip.system.DefaultRV32Config.fir@23633.4]
  assign _T_152_2 = QueueCompatibility_7_io_enq_ready; // @[UserYanker.scala 68:25:freechips.rocketchip.system.DefaultRV32Config.fir@23615.4 UserYanker.scala 68:25:freechips.rocketchip.system.DefaultRV32Config.fir@23619.4]
  assign _GEN_66 = 4'h2 == auto_in_aw_bits_id ? _T_152_2 : _GEN_65; // @[UserYanker.scala 69:36:freechips.rocketchip.system.DefaultRV32Config.fir@23633.4]
  assign _T_152_3 = QueueCompatibility_8_io_enq_ready; // @[UserYanker.scala 68:25:freechips.rocketchip.system.DefaultRV32Config.fir@23615.4 UserYanker.scala 68:25:freechips.rocketchip.system.DefaultRV32Config.fir@23620.4]
  assign _GEN_67 = 4'h3 == auto_in_aw_bits_id ? _T_152_3 : _GEN_66; // @[UserYanker.scala 69:36:freechips.rocketchip.system.DefaultRV32Config.fir@23633.4]
  assign _T_152_4 = QueueCompatibility_9_io_enq_ready; // @[UserYanker.scala 68:25:freechips.rocketchip.system.DefaultRV32Config.fir@23615.4 UserYanker.scala 68:25:freechips.rocketchip.system.DefaultRV32Config.fir@23621.4]
  assign _GEN_68 = 4'h4 == auto_in_aw_bits_id ? _T_152_4 : _GEN_67; // @[UserYanker.scala 69:36:freechips.rocketchip.system.DefaultRV32Config.fir@23633.4]
  assign _GEN_69 = 4'h5 == auto_in_aw_bits_id ? 1'h0 : _GEN_68; // @[UserYanker.scala 69:36:freechips.rocketchip.system.DefaultRV32Config.fir@23633.4]
  assign _GEN_70 = 4'h6 == auto_in_aw_bits_id ? 1'h0 : _GEN_69; // @[UserYanker.scala 69:36:freechips.rocketchip.system.DefaultRV32Config.fir@23633.4]
  assign _GEN_71 = 4'h7 == auto_in_aw_bits_id ? 1'h0 : _GEN_70; // @[UserYanker.scala 69:36:freechips.rocketchip.system.DefaultRV32Config.fir@23633.4]
  assign _GEN_72 = 4'h8 == auto_in_aw_bits_id ? 1'h0 : _GEN_71; // @[UserYanker.scala 69:36:freechips.rocketchip.system.DefaultRV32Config.fir@23633.4]
  assign _GEN_73 = 4'h9 == auto_in_aw_bits_id ? 1'h0 : _GEN_72; // @[UserYanker.scala 69:36:freechips.rocketchip.system.DefaultRV32Config.fir@23633.4]
  assign _GEN_74 = 4'ha == auto_in_aw_bits_id ? 1'h0 : _GEN_73; // @[UserYanker.scala 69:36:freechips.rocketchip.system.DefaultRV32Config.fir@23633.4]
  assign _GEN_75 = 4'hb == auto_in_aw_bits_id ? 1'h0 : _GEN_74; // @[UserYanker.scala 69:36:freechips.rocketchip.system.DefaultRV32Config.fir@23633.4]
  assign _GEN_76 = 4'hc == auto_in_aw_bits_id ? 1'h0 : _GEN_75; // @[UserYanker.scala 69:36:freechips.rocketchip.system.DefaultRV32Config.fir@23633.4]
  assign _GEN_77 = 4'hd == auto_in_aw_bits_id ? 1'h0 : _GEN_76; // @[UserYanker.scala 69:36:freechips.rocketchip.system.DefaultRV32Config.fir@23633.4]
  assign _GEN_78 = 4'he == auto_in_aw_bits_id ? 1'h0 : _GEN_77; // @[UserYanker.scala 69:36:freechips.rocketchip.system.DefaultRV32Config.fir@23633.4]
  assign _GEN_79 = 4'hf == auto_in_aw_bits_id ? 1'h0 : _GEN_78; // @[UserYanker.scala 69:36:freechips.rocketchip.system.DefaultRV32Config.fir@23633.4]
  assign _T_157 = ~auto_out_b_valid; // @[UserYanker.scala 76:15:freechips.rocketchip.system.DefaultRV32Config.fir@23682.4]
  assign _T_155_0 = QueueCompatibility_5_io_deq_valid; // @[UserYanker.scala 74:24:freechips.rocketchip.system.DefaultRV32Config.fir@23646.4 UserYanker.scala 74:24:freechips.rocketchip.system.DefaultRV32Config.fir@23648.4]
  assign _T_155_1 = QueueCompatibility_6_io_deq_valid; // @[UserYanker.scala 74:24:freechips.rocketchip.system.DefaultRV32Config.fir@23646.4 UserYanker.scala 74:24:freechips.rocketchip.system.DefaultRV32Config.fir@23649.4]
  assign _GEN_81 = 4'h1 == auto_out_b_bits_id ? _T_155_1 : _T_155_0; // @[UserYanker.scala 76:28:freechips.rocketchip.system.DefaultRV32Config.fir@23683.4]
  assign _T_155_2 = QueueCompatibility_7_io_deq_valid; // @[UserYanker.scala 74:24:freechips.rocketchip.system.DefaultRV32Config.fir@23646.4 UserYanker.scala 74:24:freechips.rocketchip.system.DefaultRV32Config.fir@23650.4]
  assign _GEN_82 = 4'h2 == auto_out_b_bits_id ? _T_155_2 : _GEN_81; // @[UserYanker.scala 76:28:freechips.rocketchip.system.DefaultRV32Config.fir@23683.4]
  assign _T_155_3 = QueueCompatibility_8_io_deq_valid; // @[UserYanker.scala 74:24:freechips.rocketchip.system.DefaultRV32Config.fir@23646.4 UserYanker.scala 74:24:freechips.rocketchip.system.DefaultRV32Config.fir@23651.4]
  assign _GEN_83 = 4'h3 == auto_out_b_bits_id ? _T_155_3 : _GEN_82; // @[UserYanker.scala 76:28:freechips.rocketchip.system.DefaultRV32Config.fir@23683.4]
  assign _T_155_4 = QueueCompatibility_9_io_deq_valid; // @[UserYanker.scala 74:24:freechips.rocketchip.system.DefaultRV32Config.fir@23646.4 UserYanker.scala 74:24:freechips.rocketchip.system.DefaultRV32Config.fir@23652.4]
  assign _GEN_84 = 4'h4 == auto_out_b_bits_id ? _T_155_4 : _GEN_83; // @[UserYanker.scala 76:28:freechips.rocketchip.system.DefaultRV32Config.fir@23683.4]
  assign _GEN_85 = 4'h5 == auto_out_b_bits_id ? 1'h0 : _GEN_84; // @[UserYanker.scala 76:28:freechips.rocketchip.system.DefaultRV32Config.fir@23683.4]
  assign _GEN_86 = 4'h6 == auto_out_b_bits_id ? 1'h0 : _GEN_85; // @[UserYanker.scala 76:28:freechips.rocketchip.system.DefaultRV32Config.fir@23683.4]
  assign _GEN_87 = 4'h7 == auto_out_b_bits_id ? 1'h0 : _GEN_86; // @[UserYanker.scala 76:28:freechips.rocketchip.system.DefaultRV32Config.fir@23683.4]
  assign _GEN_88 = 4'h8 == auto_out_b_bits_id ? 1'h0 : _GEN_87; // @[UserYanker.scala 76:28:freechips.rocketchip.system.DefaultRV32Config.fir@23683.4]
  assign _GEN_89 = 4'h9 == auto_out_b_bits_id ? 1'h0 : _GEN_88; // @[UserYanker.scala 76:28:freechips.rocketchip.system.DefaultRV32Config.fir@23683.4]
  assign _GEN_90 = 4'ha == auto_out_b_bits_id ? 1'h0 : _GEN_89; // @[UserYanker.scala 76:28:freechips.rocketchip.system.DefaultRV32Config.fir@23683.4]
  assign _GEN_91 = 4'hb == auto_out_b_bits_id ? 1'h0 : _GEN_90; // @[UserYanker.scala 76:28:freechips.rocketchip.system.DefaultRV32Config.fir@23683.4]
  assign _GEN_92 = 4'hc == auto_out_b_bits_id ? 1'h0 : _GEN_91; // @[UserYanker.scala 76:28:freechips.rocketchip.system.DefaultRV32Config.fir@23683.4]
  assign _GEN_93 = 4'hd == auto_out_b_bits_id ? 1'h0 : _GEN_92; // @[UserYanker.scala 76:28:freechips.rocketchip.system.DefaultRV32Config.fir@23683.4]
  assign _GEN_94 = 4'he == auto_out_b_bits_id ? 1'h0 : _GEN_93; // @[UserYanker.scala 76:28:freechips.rocketchip.system.DefaultRV32Config.fir@23683.4]
  assign _GEN_95 = 4'hf == auto_out_b_bits_id ? 1'h0 : _GEN_94; // @[UserYanker.scala 76:28:freechips.rocketchip.system.DefaultRV32Config.fir@23683.4]
  assign _T_158 = _T_157 | _GEN_95; // @[UserYanker.scala 76:28:freechips.rocketchip.system.DefaultRV32Config.fir@23683.4]
  assign _T_160 = _T_158 | reset; // @[UserYanker.scala 76:14:freechips.rocketchip.system.DefaultRV32Config.fir@23685.4]
  assign _T_161 = ~_T_160; // @[UserYanker.scala 76:14:freechips.rocketchip.system.DefaultRV32Config.fir@23686.4]
  assign _T_156_0_tl_state_size = QueueCompatibility_5_io_deq_bits_tl_state_size; // @[UserYanker.scala 75:23:freechips.rocketchip.system.DefaultRV32Config.fir@23664.4 UserYanker.scala 75:23:freechips.rocketchip.system.DefaultRV32Config.fir@23666.4]
  assign _T_156_0_tl_state_source = QueueCompatibility_5_io_deq_bits_tl_state_source; // @[UserYanker.scala 75:23:freechips.rocketchip.system.DefaultRV32Config.fir@23664.4 UserYanker.scala 75:23:freechips.rocketchip.system.DefaultRV32Config.fir@23666.4]
  assign _T_156_1_tl_state_size = QueueCompatibility_6_io_deq_bits_tl_state_size; // @[UserYanker.scala 75:23:freechips.rocketchip.system.DefaultRV32Config.fir@23664.4 UserYanker.scala 75:23:freechips.rocketchip.system.DefaultRV32Config.fir@23667.4]
  assign _GEN_98 = 4'h1 == auto_out_b_bits_id ? _T_156_1_tl_state_size : _T_156_0_tl_state_size; // @[BundleMap.scala 248:19:freechips.rocketchip.system.DefaultRV32Config.fir@23697.4]
  assign _T_156_1_tl_state_source = QueueCompatibility_6_io_deq_bits_tl_state_source; // @[UserYanker.scala 75:23:freechips.rocketchip.system.DefaultRV32Config.fir@23664.4 UserYanker.scala 75:23:freechips.rocketchip.system.DefaultRV32Config.fir@23667.4]
  assign _GEN_99 = 4'h1 == auto_out_b_bits_id ? _T_156_1_tl_state_source : _T_156_0_tl_state_source; // @[BundleMap.scala 248:19:freechips.rocketchip.system.DefaultRV32Config.fir@23697.4]
  assign _T_156_2_tl_state_size = QueueCompatibility_7_io_deq_bits_tl_state_size; // @[UserYanker.scala 75:23:freechips.rocketchip.system.DefaultRV32Config.fir@23664.4 UserYanker.scala 75:23:freechips.rocketchip.system.DefaultRV32Config.fir@23668.4]
  assign _GEN_100 = 4'h2 == auto_out_b_bits_id ? _T_156_2_tl_state_size : _GEN_98; // @[BundleMap.scala 248:19:freechips.rocketchip.system.DefaultRV32Config.fir@23697.4]
  assign _T_156_2_tl_state_source = QueueCompatibility_7_io_deq_bits_tl_state_source; // @[UserYanker.scala 75:23:freechips.rocketchip.system.DefaultRV32Config.fir@23664.4 UserYanker.scala 75:23:freechips.rocketchip.system.DefaultRV32Config.fir@23668.4]
  assign _GEN_101 = 4'h2 == auto_out_b_bits_id ? _T_156_2_tl_state_source : _GEN_99; // @[BundleMap.scala 248:19:freechips.rocketchip.system.DefaultRV32Config.fir@23697.4]
  assign _T_156_3_tl_state_size = QueueCompatibility_8_io_deq_bits_tl_state_size; // @[UserYanker.scala 75:23:freechips.rocketchip.system.DefaultRV32Config.fir@23664.4 UserYanker.scala 75:23:freechips.rocketchip.system.DefaultRV32Config.fir@23669.4]
  assign _GEN_102 = 4'h3 == auto_out_b_bits_id ? _T_156_3_tl_state_size : _GEN_100; // @[BundleMap.scala 248:19:freechips.rocketchip.system.DefaultRV32Config.fir@23697.4]
  assign _T_156_3_tl_state_source = QueueCompatibility_8_io_deq_bits_tl_state_source; // @[UserYanker.scala 75:23:freechips.rocketchip.system.DefaultRV32Config.fir@23664.4 UserYanker.scala 75:23:freechips.rocketchip.system.DefaultRV32Config.fir@23669.4]
  assign _GEN_103 = 4'h3 == auto_out_b_bits_id ? _T_156_3_tl_state_source : _GEN_101; // @[BundleMap.scala 248:19:freechips.rocketchip.system.DefaultRV32Config.fir@23697.4]
  assign _T_156_4_tl_state_size = QueueCompatibility_9_io_deq_bits_tl_state_size; // @[UserYanker.scala 75:23:freechips.rocketchip.system.DefaultRV32Config.fir@23664.4 UserYanker.scala 75:23:freechips.rocketchip.system.DefaultRV32Config.fir@23670.4]
  assign _GEN_104 = 4'h4 == auto_out_b_bits_id ? _T_156_4_tl_state_size : _GEN_102; // @[BundleMap.scala 248:19:freechips.rocketchip.system.DefaultRV32Config.fir@23697.4]
  assign _T_156_4_tl_state_source = QueueCompatibility_9_io_deq_bits_tl_state_source; // @[UserYanker.scala 75:23:freechips.rocketchip.system.DefaultRV32Config.fir@23664.4 UserYanker.scala 75:23:freechips.rocketchip.system.DefaultRV32Config.fir@23670.4]
  assign _GEN_105 = 4'h4 == auto_out_b_bits_id ? _T_156_4_tl_state_source : _GEN_103; // @[BundleMap.scala 248:19:freechips.rocketchip.system.DefaultRV32Config.fir@23697.4]
  assign _GEN_106 = 4'h5 == auto_out_b_bits_id ? 4'h0 : _GEN_104; // @[BundleMap.scala 248:19:freechips.rocketchip.system.DefaultRV32Config.fir@23697.4]
  assign _GEN_107 = 4'h5 == auto_out_b_bits_id ? 5'h0 : _GEN_105; // @[BundleMap.scala 248:19:freechips.rocketchip.system.DefaultRV32Config.fir@23697.4]
  assign _GEN_108 = 4'h6 == auto_out_b_bits_id ? 4'h0 : _GEN_106; // @[BundleMap.scala 248:19:freechips.rocketchip.system.DefaultRV32Config.fir@23697.4]
  assign _GEN_109 = 4'h6 == auto_out_b_bits_id ? 5'h0 : _GEN_107; // @[BundleMap.scala 248:19:freechips.rocketchip.system.DefaultRV32Config.fir@23697.4]
  assign _GEN_110 = 4'h7 == auto_out_b_bits_id ? 4'h0 : _GEN_108; // @[BundleMap.scala 248:19:freechips.rocketchip.system.DefaultRV32Config.fir@23697.4]
  assign _GEN_111 = 4'h7 == auto_out_b_bits_id ? 5'h0 : _GEN_109; // @[BundleMap.scala 248:19:freechips.rocketchip.system.DefaultRV32Config.fir@23697.4]
  assign _GEN_112 = 4'h8 == auto_out_b_bits_id ? 4'h0 : _GEN_110; // @[BundleMap.scala 248:19:freechips.rocketchip.system.DefaultRV32Config.fir@23697.4]
  assign _GEN_113 = 4'h8 == auto_out_b_bits_id ? 5'h0 : _GEN_111; // @[BundleMap.scala 248:19:freechips.rocketchip.system.DefaultRV32Config.fir@23697.4]
  assign _GEN_114 = 4'h9 == auto_out_b_bits_id ? 4'h0 : _GEN_112; // @[BundleMap.scala 248:19:freechips.rocketchip.system.DefaultRV32Config.fir@23697.4]
  assign _GEN_115 = 4'h9 == auto_out_b_bits_id ? 5'h0 : _GEN_113; // @[BundleMap.scala 248:19:freechips.rocketchip.system.DefaultRV32Config.fir@23697.4]
  assign _GEN_116 = 4'ha == auto_out_b_bits_id ? 4'h0 : _GEN_114; // @[BundleMap.scala 248:19:freechips.rocketchip.system.DefaultRV32Config.fir@23697.4]
  assign _GEN_117 = 4'ha == auto_out_b_bits_id ? 5'h0 : _GEN_115; // @[BundleMap.scala 248:19:freechips.rocketchip.system.DefaultRV32Config.fir@23697.4]
  assign _GEN_118 = 4'hb == auto_out_b_bits_id ? 4'h0 : _GEN_116; // @[BundleMap.scala 248:19:freechips.rocketchip.system.DefaultRV32Config.fir@23697.4]
  assign _GEN_119 = 4'hb == auto_out_b_bits_id ? 5'h0 : _GEN_117; // @[BundleMap.scala 248:19:freechips.rocketchip.system.DefaultRV32Config.fir@23697.4]
  assign _GEN_120 = 4'hc == auto_out_b_bits_id ? 4'h0 : _GEN_118; // @[BundleMap.scala 248:19:freechips.rocketchip.system.DefaultRV32Config.fir@23697.4]
  assign _GEN_121 = 4'hc == auto_out_b_bits_id ? 5'h0 : _GEN_119; // @[BundleMap.scala 248:19:freechips.rocketchip.system.DefaultRV32Config.fir@23697.4]
  assign _GEN_122 = 4'hd == auto_out_b_bits_id ? 4'h0 : _GEN_120; // @[BundleMap.scala 248:19:freechips.rocketchip.system.DefaultRV32Config.fir@23697.4]
  assign _GEN_123 = 4'hd == auto_out_b_bits_id ? 5'h0 : _GEN_121; // @[BundleMap.scala 248:19:freechips.rocketchip.system.DefaultRV32Config.fir@23697.4]
  assign _GEN_124 = 4'he == auto_out_b_bits_id ? 4'h0 : _GEN_122; // @[BundleMap.scala 248:19:freechips.rocketchip.system.DefaultRV32Config.fir@23697.4]
  assign _GEN_125 = 4'he == auto_out_b_bits_id ? 5'h0 : _GEN_123; // @[BundleMap.scala 248:19:freechips.rocketchip.system.DefaultRV32Config.fir@23697.4]
  assign _T_163 = 16'h1 << auto_in_aw_bits_id; // @[OneHot.scala 65:12:freechips.rocketchip.system.DefaultRV32Config.fir@23700.4]
  assign _T_182 = 16'h1 << auto_out_b_bits_id; // @[OneHot.scala 65:12:freechips.rocketchip.system.DefaultRV32Config.fir@23719.4]
  assign _T_200 = auto_out_b_valid & auto_in_b_ready; // @[UserYanker.scala 83:37:freechips.rocketchip.system.DefaultRV32Config.fir@23737.4]
  assign _T_202 = auto_in_aw_valid & auto_out_aw_ready; // @[UserYanker.scala 84:37:freechips.rocketchip.system.DefaultRV32Config.fir@23740.4]
  assign auto_in_aw_ready = auto_out_aw_ready & _GEN_79; // @[LazyModule.scala 303:16:freechips.rocketchip.system.DefaultRV32Config.fir@23262.4]
  assign auto_in_w_ready = auto_out_w_ready; // @[LazyModule.scala 303:16:freechips.rocketchip.system.DefaultRV32Config.fir@23262.4]
  assign auto_in_b_valid = auto_out_b_valid; // @[LazyModule.scala 303:16:freechips.rocketchip.system.DefaultRV32Config.fir@23262.4]
  assign auto_in_b_bits_id = auto_out_b_bits_id; // @[LazyModule.scala 303:16:freechips.rocketchip.system.DefaultRV32Config.fir@23262.4]
  assign auto_in_b_bits_resp = auto_out_b_bits_resp; // @[LazyModule.scala 303:16:freechips.rocketchip.system.DefaultRV32Config.fir@23262.4]
  assign auto_in_b_bits_echo_tl_state_size = 4'hf == auto_out_b_bits_id ? 4'h0 : _GEN_124; // @[LazyModule.scala 303:16:freechips.rocketchip.system.DefaultRV32Config.fir@23262.4]
  assign auto_in_b_bits_echo_tl_state_source = 4'hf == auto_out_b_bits_id ? 5'h0 : _GEN_125; // @[LazyModule.scala 303:16:freechips.rocketchip.system.DefaultRV32Config.fir@23262.4]
  assign auto_in_ar_ready = auto_out_ar_ready & _GEN_15; // @[LazyModule.scala 303:16:freechips.rocketchip.system.DefaultRV32Config.fir@23262.4]
  assign auto_in_r_valid = auto_out_r_valid; // @[LazyModule.scala 303:16:freechips.rocketchip.system.DefaultRV32Config.fir@23262.4]
  assign auto_in_r_bits_id = auto_out_r_bits_id; // @[LazyModule.scala 303:16:freechips.rocketchip.system.DefaultRV32Config.fir@23262.4]
  assign auto_in_r_bits_data = auto_out_r_bits_data; // @[LazyModule.scala 303:16:freechips.rocketchip.system.DefaultRV32Config.fir@23262.4]
  assign auto_in_r_bits_resp = auto_out_r_bits_resp; // @[LazyModule.scala 303:16:freechips.rocketchip.system.DefaultRV32Config.fir@23262.4]
  assign auto_in_r_bits_echo_tl_state_size = 4'hf == auto_out_r_bits_id ? 4'h0 : _GEN_60; // @[LazyModule.scala 303:16:freechips.rocketchip.system.DefaultRV32Config.fir@23262.4]
  assign auto_in_r_bits_echo_tl_state_source = 4'hf == auto_out_r_bits_id ? 5'h0 : _GEN_61; // @[LazyModule.scala 303:16:freechips.rocketchip.system.DefaultRV32Config.fir@23262.4]
  assign auto_in_r_bits_last = auto_out_r_bits_last; // @[LazyModule.scala 303:16:freechips.rocketchip.system.DefaultRV32Config.fir@23262.4]
  assign auto_out_aw_valid = auto_in_aw_valid & _GEN_79; // @[LazyModule.scala 305:12:freechips.rocketchip.system.DefaultRV32Config.fir@23261.4]
  assign auto_out_aw_bits_id = auto_in_aw_bits_id; // @[LazyModule.scala 305:12:freechips.rocketchip.system.DefaultRV32Config.fir@23261.4]
  assign auto_out_aw_bits_addr = auto_in_aw_bits_addr; // @[LazyModule.scala 305:12:freechips.rocketchip.system.DefaultRV32Config.fir@23261.4]
  assign auto_out_aw_bits_len = auto_in_aw_bits_len; // @[LazyModule.scala 305:12:freechips.rocketchip.system.DefaultRV32Config.fir@23261.4]
  assign auto_out_aw_bits_size = auto_in_aw_bits_size; // @[LazyModule.scala 305:12:freechips.rocketchip.system.DefaultRV32Config.fir@23261.4]
  assign auto_out_aw_bits_burst = auto_in_aw_bits_burst; // @[LazyModule.scala 305:12:freechips.rocketchip.system.DefaultRV32Config.fir@23261.4]
  assign auto_out_aw_bits_lock = auto_in_aw_bits_lock; // @[LazyModule.scala 305:12:freechips.rocketchip.system.DefaultRV32Config.fir@23261.4]
  assign auto_out_aw_bits_cache = auto_in_aw_bits_cache; // @[LazyModule.scala 305:12:freechips.rocketchip.system.DefaultRV32Config.fir@23261.4]
  assign auto_out_aw_bits_prot = auto_in_aw_bits_prot; // @[LazyModule.scala 305:12:freechips.rocketchip.system.DefaultRV32Config.fir@23261.4]
  assign auto_out_aw_bits_qos = auto_in_aw_bits_qos; // @[LazyModule.scala 305:12:freechips.rocketchip.system.DefaultRV32Config.fir@23261.4]
  assign auto_out_w_valid = auto_in_w_valid; // @[LazyModule.scala 305:12:freechips.rocketchip.system.DefaultRV32Config.fir@23261.4]
  assign auto_out_w_bits_data = auto_in_w_bits_data; // @[LazyModule.scala 305:12:freechips.rocketchip.system.DefaultRV32Config.fir@23261.4]
  assign auto_out_w_bits_strb = auto_in_w_bits_strb; // @[LazyModule.scala 305:12:freechips.rocketchip.system.DefaultRV32Config.fir@23261.4]
  assign auto_out_w_bits_last = auto_in_w_bits_last; // @[LazyModule.scala 305:12:freechips.rocketchip.system.DefaultRV32Config.fir@23261.4]
  assign auto_out_b_ready = auto_in_b_ready; // @[LazyModule.scala 305:12:freechips.rocketchip.system.DefaultRV32Config.fir@23261.4]
  assign auto_out_ar_valid = auto_in_ar_valid & _GEN_15; // @[LazyModule.scala 305:12:freechips.rocketchip.system.DefaultRV32Config.fir@23261.4]
  assign auto_out_ar_bits_id = auto_in_ar_bits_id; // @[LazyModule.scala 305:12:freechips.rocketchip.system.DefaultRV32Config.fir@23261.4]
  assign auto_out_ar_bits_addr = auto_in_ar_bits_addr; // @[LazyModule.scala 305:12:freechips.rocketchip.system.DefaultRV32Config.fir@23261.4]
  assign auto_out_ar_bits_len = auto_in_ar_bits_len; // @[LazyModule.scala 305:12:freechips.rocketchip.system.DefaultRV32Config.fir@23261.4]
  assign auto_out_ar_bits_size = auto_in_ar_bits_size; // @[LazyModule.scala 305:12:freechips.rocketchip.system.DefaultRV32Config.fir@23261.4]
  assign auto_out_ar_bits_burst = auto_in_ar_bits_burst; // @[LazyModule.scala 305:12:freechips.rocketchip.system.DefaultRV32Config.fir@23261.4]
  assign auto_out_ar_bits_lock = auto_in_ar_bits_lock; // @[LazyModule.scala 305:12:freechips.rocketchip.system.DefaultRV32Config.fir@23261.4]
  assign auto_out_ar_bits_cache = auto_in_ar_bits_cache; // @[LazyModule.scala 305:12:freechips.rocketchip.system.DefaultRV32Config.fir@23261.4]
  assign auto_out_ar_bits_prot = auto_in_ar_bits_prot; // @[LazyModule.scala 305:12:freechips.rocketchip.system.DefaultRV32Config.fir@23261.4]
  assign auto_out_ar_bits_qos = auto_in_ar_bits_qos; // @[LazyModule.scala 305:12:freechips.rocketchip.system.DefaultRV32Config.fir@23261.4]
  assign auto_out_r_ready = auto_in_r_ready; // @[LazyModule.scala 305:12:freechips.rocketchip.system.DefaultRV32Config.fir@23261.4]
  assign QueueCompatibility_clock = clock; // @[:freechips.rocketchip.system.DefaultRV32Config.fir@23265.4]
  assign QueueCompatibility_reset = reset; // @[:freechips.rocketchip.system.DefaultRV32Config.fir@23266.4]
  assign QueueCompatibility_io_enq_valid = _T_75 & _T_35[0]; // @[UserYanker.scala 63:21:freechips.rocketchip.system.DefaultRV32Config.fir@23477.4]
  assign QueueCompatibility_io_enq_bits_tl_state_size = auto_in_ar_bits_echo_tl_state_size; // @[BundleMap.scala 248:19:freechips.rocketchip.system.DefaultRV32Config.fir@23479.4]
  assign QueueCompatibility_io_enq_bits_tl_state_source = auto_in_ar_bits_echo_tl_state_source; // @[BundleMap.scala 248:19:freechips.rocketchip.system.DefaultRV32Config.fir@23478.4]
  assign QueueCompatibility_io_deq_ready = _T_73 & auto_out_r_bits_last; // @[UserYanker.scala 62:21:freechips.rocketchip.system.DefaultRV32Config.fir@23474.4]
  assign QueueCompatibility_1_clock = clock; // @[:freechips.rocketchip.system.DefaultRV32Config.fir@23269.4]
  assign QueueCompatibility_1_reset = reset; // @[:freechips.rocketchip.system.DefaultRV32Config.fir@23270.4]
  assign QueueCompatibility_1_io_enq_valid = _T_75 & _T_35[1]; // @[UserYanker.scala 63:21:freechips.rocketchip.system.DefaultRV32Config.fir@23486.4]
  assign QueueCompatibility_1_io_enq_bits_tl_state_size = auto_in_ar_bits_echo_tl_state_size; // @[BundleMap.scala 248:19:freechips.rocketchip.system.DefaultRV32Config.fir@23488.4]
  assign QueueCompatibility_1_io_enq_bits_tl_state_source = auto_in_ar_bits_echo_tl_state_source; // @[BundleMap.scala 248:19:freechips.rocketchip.system.DefaultRV32Config.fir@23487.4]
  assign QueueCompatibility_1_io_deq_ready = _T_78 & auto_out_r_bits_last; // @[UserYanker.scala 62:21:freechips.rocketchip.system.DefaultRV32Config.fir@23483.4]
  assign QueueCompatibility_2_clock = clock; // @[:freechips.rocketchip.system.DefaultRV32Config.fir@23273.4]
  assign QueueCompatibility_2_reset = reset; // @[:freechips.rocketchip.system.DefaultRV32Config.fir@23274.4]
  assign QueueCompatibility_2_io_enq_valid = _T_75 & _T_35[2]; // @[UserYanker.scala 63:21:freechips.rocketchip.system.DefaultRV32Config.fir@23495.4]
  assign QueueCompatibility_2_io_enq_bits_tl_state_size = auto_in_ar_bits_echo_tl_state_size; // @[BundleMap.scala 248:19:freechips.rocketchip.system.DefaultRV32Config.fir@23497.4]
  assign QueueCompatibility_2_io_enq_bits_tl_state_source = auto_in_ar_bits_echo_tl_state_source; // @[BundleMap.scala 248:19:freechips.rocketchip.system.DefaultRV32Config.fir@23496.4]
  assign QueueCompatibility_2_io_deq_ready = _T_83 & auto_out_r_bits_last; // @[UserYanker.scala 62:21:freechips.rocketchip.system.DefaultRV32Config.fir@23492.4]
  assign QueueCompatibility_3_clock = clock; // @[:freechips.rocketchip.system.DefaultRV32Config.fir@23277.4]
  assign QueueCompatibility_3_reset = reset; // @[:freechips.rocketchip.system.DefaultRV32Config.fir@23278.4]
  assign QueueCompatibility_3_io_enq_valid = _T_75 & _T_35[3]; // @[UserYanker.scala 63:21:freechips.rocketchip.system.DefaultRV32Config.fir@23504.4]
  assign QueueCompatibility_3_io_enq_bits_tl_state_size = auto_in_ar_bits_echo_tl_state_size; // @[BundleMap.scala 248:19:freechips.rocketchip.system.DefaultRV32Config.fir@23506.4]
  assign QueueCompatibility_3_io_enq_bits_tl_state_source = auto_in_ar_bits_echo_tl_state_source; // @[BundleMap.scala 248:19:freechips.rocketchip.system.DefaultRV32Config.fir@23505.4]
  assign QueueCompatibility_3_io_deq_ready = _T_88 & auto_out_r_bits_last; // @[UserYanker.scala 62:21:freechips.rocketchip.system.DefaultRV32Config.fir@23501.4]
  assign QueueCompatibility_4_clock = clock; // @[:freechips.rocketchip.system.DefaultRV32Config.fir@23281.4]
  assign QueueCompatibility_4_reset = reset; // @[:freechips.rocketchip.system.DefaultRV32Config.fir@23282.4]
  assign QueueCompatibility_4_io_enq_valid = _T_75 & _T_35[4]; // @[UserYanker.scala 63:21:freechips.rocketchip.system.DefaultRV32Config.fir@23513.4]
  assign QueueCompatibility_4_io_enq_bits_tl_state_size = auto_in_ar_bits_echo_tl_state_size; // @[BundleMap.scala 248:19:freechips.rocketchip.system.DefaultRV32Config.fir@23515.4]
  assign QueueCompatibility_4_io_enq_bits_tl_state_source = auto_in_ar_bits_echo_tl_state_source; // @[BundleMap.scala 248:19:freechips.rocketchip.system.DefaultRV32Config.fir@23514.4]
  assign QueueCompatibility_4_io_deq_ready = _T_93 & auto_out_r_bits_last; // @[UserYanker.scala 62:21:freechips.rocketchip.system.DefaultRV32Config.fir@23510.4]
  assign QueueCompatibility_5_clock = clock; // @[:freechips.rocketchip.system.DefaultRV32Config.fir@23307.4]
  assign QueueCompatibility_5_reset = reset; // @[:freechips.rocketchip.system.DefaultRV32Config.fir@23308.4]
  assign QueueCompatibility_5_io_enq_valid = _T_202 & _T_163[0]; // @[UserYanker.scala 84:21:freechips.rocketchip.system.DefaultRV32Config.fir@23742.4]
  assign QueueCompatibility_5_io_enq_bits_tl_state_size = auto_in_aw_bits_echo_tl_state_size; // @[BundleMap.scala 248:19:freechips.rocketchip.system.DefaultRV32Config.fir@23744.4]
  assign QueueCompatibility_5_io_enq_bits_tl_state_source = auto_in_aw_bits_echo_tl_state_source; // @[BundleMap.scala 248:19:freechips.rocketchip.system.DefaultRV32Config.fir@23743.4]
  assign QueueCompatibility_5_io_deq_ready = _T_200 & _T_182[0]; // @[UserYanker.scala 83:21:freechips.rocketchip.system.DefaultRV32Config.fir@23739.4]
  assign QueueCompatibility_6_clock = clock; // @[:freechips.rocketchip.system.DefaultRV32Config.fir@23311.4]
  assign QueueCompatibility_6_reset = reset; // @[:freechips.rocketchip.system.DefaultRV32Config.fir@23312.4]
  assign QueueCompatibility_6_io_enq_valid = _T_202 & _T_163[1]; // @[UserYanker.scala 84:21:freechips.rocketchip.system.DefaultRV32Config.fir@23750.4]
  assign QueueCompatibility_6_io_enq_bits_tl_state_size = auto_in_aw_bits_echo_tl_state_size; // @[BundleMap.scala 248:19:freechips.rocketchip.system.DefaultRV32Config.fir@23752.4]
  assign QueueCompatibility_6_io_enq_bits_tl_state_source = auto_in_aw_bits_echo_tl_state_source; // @[BundleMap.scala 248:19:freechips.rocketchip.system.DefaultRV32Config.fir@23751.4]
  assign QueueCompatibility_6_io_deq_ready = _T_200 & _T_182[1]; // @[UserYanker.scala 83:21:freechips.rocketchip.system.DefaultRV32Config.fir@23747.4]
  assign QueueCompatibility_7_clock = clock; // @[:freechips.rocketchip.system.DefaultRV32Config.fir@23315.4]
  assign QueueCompatibility_7_reset = reset; // @[:freechips.rocketchip.system.DefaultRV32Config.fir@23316.4]
  assign QueueCompatibility_7_io_enq_valid = _T_202 & _T_163[2]; // @[UserYanker.scala 84:21:freechips.rocketchip.system.DefaultRV32Config.fir@23758.4]
  assign QueueCompatibility_7_io_enq_bits_tl_state_size = auto_in_aw_bits_echo_tl_state_size; // @[BundleMap.scala 248:19:freechips.rocketchip.system.DefaultRV32Config.fir@23760.4]
  assign QueueCompatibility_7_io_enq_bits_tl_state_source = auto_in_aw_bits_echo_tl_state_source; // @[BundleMap.scala 248:19:freechips.rocketchip.system.DefaultRV32Config.fir@23759.4]
  assign QueueCompatibility_7_io_deq_ready = _T_200 & _T_182[2]; // @[UserYanker.scala 83:21:freechips.rocketchip.system.DefaultRV32Config.fir@23755.4]
  assign QueueCompatibility_8_clock = clock; // @[:freechips.rocketchip.system.DefaultRV32Config.fir@23319.4]
  assign QueueCompatibility_8_reset = reset; // @[:freechips.rocketchip.system.DefaultRV32Config.fir@23320.4]
  assign QueueCompatibility_8_io_enq_valid = _T_202 & _T_163[3]; // @[UserYanker.scala 84:21:freechips.rocketchip.system.DefaultRV32Config.fir@23766.4]
  assign QueueCompatibility_8_io_enq_bits_tl_state_size = auto_in_aw_bits_echo_tl_state_size; // @[BundleMap.scala 248:19:freechips.rocketchip.system.DefaultRV32Config.fir@23768.4]
  assign QueueCompatibility_8_io_enq_bits_tl_state_source = auto_in_aw_bits_echo_tl_state_source; // @[BundleMap.scala 248:19:freechips.rocketchip.system.DefaultRV32Config.fir@23767.4]
  assign QueueCompatibility_8_io_deq_ready = _T_200 & _T_182[3]; // @[UserYanker.scala 83:21:freechips.rocketchip.system.DefaultRV32Config.fir@23763.4]
  assign QueueCompatibility_9_clock = clock; // @[:freechips.rocketchip.system.DefaultRV32Config.fir@23323.4]
  assign QueueCompatibility_9_reset = reset; // @[:freechips.rocketchip.system.DefaultRV32Config.fir@23324.4]
  assign QueueCompatibility_9_io_enq_valid = _T_202 & _T_163[4]; // @[UserYanker.scala 84:21:freechips.rocketchip.system.DefaultRV32Config.fir@23774.4]
  assign QueueCompatibility_9_io_enq_bits_tl_state_size = auto_in_aw_bits_echo_tl_state_size; // @[BundleMap.scala 248:19:freechips.rocketchip.system.DefaultRV32Config.fir@23776.4]
  assign QueueCompatibility_9_io_enq_bits_tl_state_source = auto_in_aw_bits_echo_tl_state_source; // @[BundleMap.scala 248:19:freechips.rocketchip.system.DefaultRV32Config.fir@23775.4]
  assign QueueCompatibility_9_io_deq_ready = _T_200 & _T_182[4]; // @[UserYanker.scala 83:21:freechips.rocketchip.system.DefaultRV32Config.fir@23771.4]
  always @(posedge clock) begin
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_33) begin
          $fwrite(32'h80000002,"Assertion failed\n    at UserYanker.scala:55 assert (!out.r.valid || r_valid) // Q must be ready faster than the response\n"); // @[UserYanker.scala 55:14:freechips.rocketchip.system.DefaultRV32Config.fir@23420.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_33) begin
          $fatal; // @[UserYanker.scala 55:14:freechips.rocketchip.system.DefaultRV32Config.fir@23421.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_161) begin
          $fwrite(32'h80000002,"Assertion failed\n    at UserYanker.scala:76 assert (!out.b.valid || b_valid) // Q must be ready faster than the response\n"); // @[UserYanker.scala 76:14:freechips.rocketchip.system.DefaultRV32Config.fir@23688.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_161) begin
          $fatal; // @[UserYanker.scala 76:14:freechips.rocketchip.system.DefaultRV32Config.fir@23689.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
  end
endmodule
