module ClockGroupAggregator( // @[:freechips.rocketchip.system.DefaultRV32Config.fir@44.2]
  input   auto_in_member_5_clock, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@45.4]
  input   auto_in_member_5_reset, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@45.4]
  input   auto_in_member_4_clock, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@45.4]
  input   auto_in_member_4_reset, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@45.4]
  input   auto_in_member_3_clock, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@45.4]
  input   auto_in_member_3_reset, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@45.4]
  input   auto_in_member_2_clock, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@45.4]
  input   auto_in_member_2_reset, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@45.4]
  input   auto_in_member_1_clock, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@45.4]
  input   auto_in_member_1_reset, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@45.4]
  input   auto_in_member_0_clock, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@45.4]
  input   auto_in_member_0_reset, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@45.4]
  output  auto_out_3_member_1_clock, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@45.4]
  output  auto_out_3_member_1_reset, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@45.4]
  output  auto_out_3_member_0_clock, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@45.4]
  output  auto_out_3_member_0_reset, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@45.4]
  output  auto_out_2_member_0_clock, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@45.4]
  output  auto_out_2_member_0_reset, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@45.4]
  output  auto_out_1_member_1_clock, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@45.4]
  output  auto_out_1_member_1_reset, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@45.4]
  output  auto_out_1_member_0_clock, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@45.4]
  output  auto_out_1_member_0_reset, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@45.4]
  output  auto_out_0_member_0_clock, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@45.4]
  output  auto_out_0_member_0_reset // @[:freechips.rocketchip.system.DefaultRV32Config.fir@45.4]
);
  assign auto_out_3_member_1_clock = auto_in_member_5_clock; // @[LazyModule.scala 305:12:freechips.rocketchip.system.DefaultRV32Config.fir@68.4]
  assign auto_out_3_member_1_reset = auto_in_member_5_reset; // @[LazyModule.scala 305:12:freechips.rocketchip.system.DefaultRV32Config.fir@68.4]
  assign auto_out_3_member_0_clock = auto_in_member_4_clock; // @[LazyModule.scala 305:12:freechips.rocketchip.system.DefaultRV32Config.fir@68.4]
  assign auto_out_3_member_0_reset = auto_in_member_4_reset; // @[LazyModule.scala 305:12:freechips.rocketchip.system.DefaultRV32Config.fir@68.4]
  assign auto_out_2_member_0_clock = auto_in_member_3_clock; // @[LazyModule.scala 305:12:freechips.rocketchip.system.DefaultRV32Config.fir@67.4]
  assign auto_out_2_member_0_reset = auto_in_member_3_reset; // @[LazyModule.scala 305:12:freechips.rocketchip.system.DefaultRV32Config.fir@67.4]
  assign auto_out_1_member_1_clock = auto_in_member_2_clock; // @[LazyModule.scala 305:12:freechips.rocketchip.system.DefaultRV32Config.fir@66.4]
  assign auto_out_1_member_1_reset = auto_in_member_2_reset; // @[LazyModule.scala 305:12:freechips.rocketchip.system.DefaultRV32Config.fir@66.4]
  assign auto_out_1_member_0_clock = auto_in_member_1_clock; // @[LazyModule.scala 305:12:freechips.rocketchip.system.DefaultRV32Config.fir@66.4]
  assign auto_out_1_member_0_reset = auto_in_member_1_reset; // @[LazyModule.scala 305:12:freechips.rocketchip.system.DefaultRV32Config.fir@66.4]
  assign auto_out_0_member_0_clock = auto_in_member_0_clock; // @[LazyModule.scala 305:12:freechips.rocketchip.system.DefaultRV32Config.fir@65.4]
  assign auto_out_0_member_0_reset = auto_in_member_0_reset; // @[LazyModule.scala 305:12:freechips.rocketchip.system.DefaultRV32Config.fir@65.4]
endmodule
