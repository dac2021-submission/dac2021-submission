module PMPChecker( // @[:freechips.rocketchip.system.DefaultRV32Config.fir@175636.2]
  input  [1:0]  io_prv, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@175639.4]
  input         io_pmp_0_cfg_l, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@175639.4]
  input  [1:0]  io_pmp_0_cfg_a, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@175639.4]
  input         io_pmp_0_cfg_x, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@175639.4]
  input         io_pmp_0_cfg_w, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@175639.4]
  input         io_pmp_0_cfg_r, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@175639.4]
  input  [29:0] io_pmp_0_addr, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@175639.4]
  input  [31:0] io_pmp_0_mask, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@175639.4]
  input         io_pmp_1_cfg_l, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@175639.4]
  input  [1:0]  io_pmp_1_cfg_a, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@175639.4]
  input         io_pmp_1_cfg_x, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@175639.4]
  input         io_pmp_1_cfg_w, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@175639.4]
  input         io_pmp_1_cfg_r, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@175639.4]
  input  [29:0] io_pmp_1_addr, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@175639.4]
  input  [31:0] io_pmp_1_mask, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@175639.4]
  input         io_pmp_2_cfg_l, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@175639.4]
  input  [1:0]  io_pmp_2_cfg_a, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@175639.4]
  input         io_pmp_2_cfg_x, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@175639.4]
  input         io_pmp_2_cfg_w, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@175639.4]
  input         io_pmp_2_cfg_r, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@175639.4]
  input  [29:0] io_pmp_2_addr, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@175639.4]
  input  [31:0] io_pmp_2_mask, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@175639.4]
  input         io_pmp_3_cfg_l, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@175639.4]
  input  [1:0]  io_pmp_3_cfg_a, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@175639.4]
  input         io_pmp_3_cfg_x, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@175639.4]
  input         io_pmp_3_cfg_w, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@175639.4]
  input         io_pmp_3_cfg_r, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@175639.4]
  input  [29:0] io_pmp_3_addr, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@175639.4]
  input  [31:0] io_pmp_3_mask, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@175639.4]
  input         io_pmp_4_cfg_l, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@175639.4]
  input  [1:0]  io_pmp_4_cfg_a, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@175639.4]
  input         io_pmp_4_cfg_x, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@175639.4]
  input         io_pmp_4_cfg_w, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@175639.4]
  input         io_pmp_4_cfg_r, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@175639.4]
  input  [29:0] io_pmp_4_addr, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@175639.4]
  input  [31:0] io_pmp_4_mask, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@175639.4]
  input         io_pmp_5_cfg_l, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@175639.4]
  input  [1:0]  io_pmp_5_cfg_a, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@175639.4]
  input         io_pmp_5_cfg_x, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@175639.4]
  input         io_pmp_5_cfg_w, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@175639.4]
  input         io_pmp_5_cfg_r, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@175639.4]
  input  [29:0] io_pmp_5_addr, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@175639.4]
  input  [31:0] io_pmp_5_mask, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@175639.4]
  input         io_pmp_6_cfg_l, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@175639.4]
  input  [1:0]  io_pmp_6_cfg_a, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@175639.4]
  input         io_pmp_6_cfg_x, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@175639.4]
  input         io_pmp_6_cfg_w, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@175639.4]
  input         io_pmp_6_cfg_r, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@175639.4]
  input  [29:0] io_pmp_6_addr, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@175639.4]
  input  [31:0] io_pmp_6_mask, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@175639.4]
  input         io_pmp_7_cfg_l, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@175639.4]
  input  [1:0]  io_pmp_7_cfg_a, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@175639.4]
  input         io_pmp_7_cfg_x, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@175639.4]
  input         io_pmp_7_cfg_w, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@175639.4]
  input         io_pmp_7_cfg_r, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@175639.4]
  input  [29:0] io_pmp_7_addr, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@175639.4]
  input  [31:0] io_pmp_7_mask, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@175639.4]
  input  [31:0] io_addr, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@175639.4]
  output        io_r, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@175639.4]
  output        io_w, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@175639.4]
  output        io_x // @[:freechips.rocketchip.system.DefaultRV32Config.fir@175639.4]
);
  wire  default_; // @[PMP.scala 157:56:freechips.rocketchip.system.DefaultRV32Config.fir@175641.4]
  wire [31:0] _T_2; // @[PMP.scala 62:36:freechips.rocketchip.system.DefaultRV32Config.fir@175664.4]
  wire [31:0] _T_3; // @[PMP.scala 62:29:freechips.rocketchip.system.DefaultRV32Config.fir@175665.4]
  wire [31:0] _T_4; // @[PMP.scala 62:48:freechips.rocketchip.system.DefaultRV32Config.fir@175666.4]
  wire [31:0] _T_5; // @[PMP.scala 62:27:freechips.rocketchip.system.DefaultRV32Config.fir@175667.4]
  wire [31:0] _T_6; // @[PMP.scala 65:47:freechips.rocketchip.system.DefaultRV32Config.fir@175668.4]
  wire [31:0] _T_7; // @[PMP.scala 65:54:freechips.rocketchip.system.DefaultRV32Config.fir@175669.4]
  wire [31:0] _T_8; // @[PMP.scala 65:52:freechips.rocketchip.system.DefaultRV32Config.fir@175670.4]
  wire  _T_9; // @[PMP.scala 65:58:freechips.rocketchip.system.DefaultRV32Config.fir@175671.4]
  wire [31:0] _T_15; // @[PMP.scala 62:36:freechips.rocketchip.system.DefaultRV32Config.fir@175677.4]
  wire [31:0] _T_16; // @[PMP.scala 62:29:freechips.rocketchip.system.DefaultRV32Config.fir@175678.4]
  wire [31:0] _T_17; // @[PMP.scala 62:48:freechips.rocketchip.system.DefaultRV32Config.fir@175679.4]
  wire [31:0] _T_18; // @[PMP.scala 62:27:freechips.rocketchip.system.DefaultRV32Config.fir@175680.4]
  wire  _T_19; // @[PMP.scala 79:9:freechips.rocketchip.system.DefaultRV32Config.fir@175681.4]
  wire  _T_20; // @[PMP.scala 90:5:freechips.rocketchip.system.DefaultRV32Config.fir@175682.4]
  wire  _T_25; // @[PMP.scala 79:9:freechips.rocketchip.system.DefaultRV32Config.fir@175687.4]
  wire  _T_26; // @[PMP.scala 96:48:freechips.rocketchip.system.DefaultRV32Config.fir@175688.4]
  wire  _T_27; // @[PMP.scala 134:61:freechips.rocketchip.system.DefaultRV32Config.fir@175689.4]
  wire  _T_28; // @[PMP.scala 134:8:freechips.rocketchip.system.DefaultRV32Config.fir@175690.4]
  wire  _T_29; // @[PMP.scala 165:29:freechips.rocketchip.system.DefaultRV32Config.fir@175691.4]
  wire  _T_30; // @[PMP.scala 165:26:freechips.rocketchip.system.DefaultRV32Config.fir@175692.4]
  wire  _T_82; // @[PMP.scala 183:40:freechips.rocketchip.system.DefaultRV32Config.fir@175752.4]
  wire  _T_84; // @[PMP.scala 184:40:freechips.rocketchip.system.DefaultRV32Config.fir@175755.4]
  wire  _T_86; // @[PMP.scala 185:40:freechips.rocketchip.system.DefaultRV32Config.fir@175758.4]
  wire  _T_88_cfg_x; // @[PMP.scala 186:8:freechips.rocketchip.system.DefaultRV32Config.fir@175761.4]
  wire  _T_88_cfg_w; // @[PMP.scala 186:8:freechips.rocketchip.system.DefaultRV32Config.fir@175761.4]
  wire  _T_88_cfg_r; // @[PMP.scala 186:8:freechips.rocketchip.system.DefaultRV32Config.fir@175761.4]
  wire [31:0] _T_94; // @[PMP.scala 65:47:freechips.rocketchip.system.DefaultRV32Config.fir@175767.4]
  wire [31:0] _T_95; // @[PMP.scala 65:54:freechips.rocketchip.system.DefaultRV32Config.fir@175768.4]
  wire [31:0] _T_96; // @[PMP.scala 65:52:freechips.rocketchip.system.DefaultRV32Config.fir@175769.4]
  wire  _T_97; // @[PMP.scala 65:58:freechips.rocketchip.system.DefaultRV32Config.fir@175770.4]
  wire [31:0] _T_103; // @[PMP.scala 62:36:freechips.rocketchip.system.DefaultRV32Config.fir@175776.4]
  wire [31:0] _T_104; // @[PMP.scala 62:29:freechips.rocketchip.system.DefaultRV32Config.fir@175777.4]
  wire [31:0] _T_105; // @[PMP.scala 62:48:freechips.rocketchip.system.DefaultRV32Config.fir@175778.4]
  wire [31:0] _T_106; // @[PMP.scala 62:27:freechips.rocketchip.system.DefaultRV32Config.fir@175779.4]
  wire  _T_107; // @[PMP.scala 79:9:freechips.rocketchip.system.DefaultRV32Config.fir@175780.4]
  wire  _T_108; // @[PMP.scala 90:5:freechips.rocketchip.system.DefaultRV32Config.fir@175781.4]
  wire  _T_114; // @[PMP.scala 96:48:freechips.rocketchip.system.DefaultRV32Config.fir@175787.4]
  wire  _T_115; // @[PMP.scala 134:61:freechips.rocketchip.system.DefaultRV32Config.fir@175788.4]
  wire  _T_116; // @[PMP.scala 134:8:freechips.rocketchip.system.DefaultRV32Config.fir@175789.4]
  wire  _T_117; // @[PMP.scala 165:29:freechips.rocketchip.system.DefaultRV32Config.fir@175790.4]
  wire  _T_118; // @[PMP.scala 165:26:freechips.rocketchip.system.DefaultRV32Config.fir@175791.4]
  wire  _T_170; // @[PMP.scala 183:40:freechips.rocketchip.system.DefaultRV32Config.fir@175851.4]
  wire  _T_172; // @[PMP.scala 184:40:freechips.rocketchip.system.DefaultRV32Config.fir@175854.4]
  wire  _T_174; // @[PMP.scala 185:40:freechips.rocketchip.system.DefaultRV32Config.fir@175857.4]
  wire  _T_176_cfg_x; // @[PMP.scala 186:8:freechips.rocketchip.system.DefaultRV32Config.fir@175860.4]
  wire  _T_176_cfg_w; // @[PMP.scala 186:8:freechips.rocketchip.system.DefaultRV32Config.fir@175860.4]
  wire  _T_176_cfg_r; // @[PMP.scala 186:8:freechips.rocketchip.system.DefaultRV32Config.fir@175860.4]
  wire [31:0] _T_182; // @[PMP.scala 65:47:freechips.rocketchip.system.DefaultRV32Config.fir@175866.4]
  wire [31:0] _T_183; // @[PMP.scala 65:54:freechips.rocketchip.system.DefaultRV32Config.fir@175867.4]
  wire [31:0] _T_184; // @[PMP.scala 65:52:freechips.rocketchip.system.DefaultRV32Config.fir@175868.4]
  wire  _T_185; // @[PMP.scala 65:58:freechips.rocketchip.system.DefaultRV32Config.fir@175869.4]
  wire [31:0] _T_191; // @[PMP.scala 62:36:freechips.rocketchip.system.DefaultRV32Config.fir@175875.4]
  wire [31:0] _T_192; // @[PMP.scala 62:29:freechips.rocketchip.system.DefaultRV32Config.fir@175876.4]
  wire [31:0] _T_193; // @[PMP.scala 62:48:freechips.rocketchip.system.DefaultRV32Config.fir@175877.4]
  wire [31:0] _T_194; // @[PMP.scala 62:27:freechips.rocketchip.system.DefaultRV32Config.fir@175878.4]
  wire  _T_195; // @[PMP.scala 79:9:freechips.rocketchip.system.DefaultRV32Config.fir@175879.4]
  wire  _T_196; // @[PMP.scala 90:5:freechips.rocketchip.system.DefaultRV32Config.fir@175880.4]
  wire  _T_202; // @[PMP.scala 96:48:freechips.rocketchip.system.DefaultRV32Config.fir@175886.4]
  wire  _T_203; // @[PMP.scala 134:61:freechips.rocketchip.system.DefaultRV32Config.fir@175887.4]
  wire  _T_204; // @[PMP.scala 134:8:freechips.rocketchip.system.DefaultRV32Config.fir@175888.4]
  wire  _T_205; // @[PMP.scala 165:29:freechips.rocketchip.system.DefaultRV32Config.fir@175889.4]
  wire  _T_206; // @[PMP.scala 165:26:freechips.rocketchip.system.DefaultRV32Config.fir@175890.4]
  wire  _T_258; // @[PMP.scala 183:40:freechips.rocketchip.system.DefaultRV32Config.fir@175950.4]
  wire  _T_260; // @[PMP.scala 184:40:freechips.rocketchip.system.DefaultRV32Config.fir@175953.4]
  wire  _T_262; // @[PMP.scala 185:40:freechips.rocketchip.system.DefaultRV32Config.fir@175956.4]
  wire  _T_264_cfg_x; // @[PMP.scala 186:8:freechips.rocketchip.system.DefaultRV32Config.fir@175959.4]
  wire  _T_264_cfg_w; // @[PMP.scala 186:8:freechips.rocketchip.system.DefaultRV32Config.fir@175959.4]
  wire  _T_264_cfg_r; // @[PMP.scala 186:8:freechips.rocketchip.system.DefaultRV32Config.fir@175959.4]
  wire [31:0] _T_270; // @[PMP.scala 65:47:freechips.rocketchip.system.DefaultRV32Config.fir@175965.4]
  wire [31:0] _T_271; // @[PMP.scala 65:54:freechips.rocketchip.system.DefaultRV32Config.fir@175966.4]
  wire [31:0] _T_272; // @[PMP.scala 65:52:freechips.rocketchip.system.DefaultRV32Config.fir@175967.4]
  wire  _T_273; // @[PMP.scala 65:58:freechips.rocketchip.system.DefaultRV32Config.fir@175968.4]
  wire [31:0] _T_279; // @[PMP.scala 62:36:freechips.rocketchip.system.DefaultRV32Config.fir@175974.4]
  wire [31:0] _T_280; // @[PMP.scala 62:29:freechips.rocketchip.system.DefaultRV32Config.fir@175975.4]
  wire [31:0] _T_281; // @[PMP.scala 62:48:freechips.rocketchip.system.DefaultRV32Config.fir@175976.4]
  wire [31:0] _T_282; // @[PMP.scala 62:27:freechips.rocketchip.system.DefaultRV32Config.fir@175977.4]
  wire  _T_283; // @[PMP.scala 79:9:freechips.rocketchip.system.DefaultRV32Config.fir@175978.4]
  wire  _T_284; // @[PMP.scala 90:5:freechips.rocketchip.system.DefaultRV32Config.fir@175979.4]
  wire  _T_290; // @[PMP.scala 96:48:freechips.rocketchip.system.DefaultRV32Config.fir@175985.4]
  wire  _T_291; // @[PMP.scala 134:61:freechips.rocketchip.system.DefaultRV32Config.fir@175986.4]
  wire  _T_292; // @[PMP.scala 134:8:freechips.rocketchip.system.DefaultRV32Config.fir@175987.4]
  wire  _T_293; // @[PMP.scala 165:29:freechips.rocketchip.system.DefaultRV32Config.fir@175988.4]
  wire  _T_294; // @[PMP.scala 165:26:freechips.rocketchip.system.DefaultRV32Config.fir@175989.4]
  wire  _T_346; // @[PMP.scala 183:40:freechips.rocketchip.system.DefaultRV32Config.fir@176049.4]
  wire  _T_348; // @[PMP.scala 184:40:freechips.rocketchip.system.DefaultRV32Config.fir@176052.4]
  wire  _T_350; // @[PMP.scala 185:40:freechips.rocketchip.system.DefaultRV32Config.fir@176055.4]
  wire  _T_352_cfg_x; // @[PMP.scala 186:8:freechips.rocketchip.system.DefaultRV32Config.fir@176058.4]
  wire  _T_352_cfg_w; // @[PMP.scala 186:8:freechips.rocketchip.system.DefaultRV32Config.fir@176058.4]
  wire  _T_352_cfg_r; // @[PMP.scala 186:8:freechips.rocketchip.system.DefaultRV32Config.fir@176058.4]
  wire [31:0] _T_358; // @[PMP.scala 65:47:freechips.rocketchip.system.DefaultRV32Config.fir@176064.4]
  wire [31:0] _T_359; // @[PMP.scala 65:54:freechips.rocketchip.system.DefaultRV32Config.fir@176065.4]
  wire [31:0] _T_360; // @[PMP.scala 65:52:freechips.rocketchip.system.DefaultRV32Config.fir@176066.4]
  wire  _T_361; // @[PMP.scala 65:58:freechips.rocketchip.system.DefaultRV32Config.fir@176067.4]
  wire [31:0] _T_367; // @[PMP.scala 62:36:freechips.rocketchip.system.DefaultRV32Config.fir@176073.4]
  wire [31:0] _T_368; // @[PMP.scala 62:29:freechips.rocketchip.system.DefaultRV32Config.fir@176074.4]
  wire [31:0] _T_369; // @[PMP.scala 62:48:freechips.rocketchip.system.DefaultRV32Config.fir@176075.4]
  wire [31:0] _T_370; // @[PMP.scala 62:27:freechips.rocketchip.system.DefaultRV32Config.fir@176076.4]
  wire  _T_371; // @[PMP.scala 79:9:freechips.rocketchip.system.DefaultRV32Config.fir@176077.4]
  wire  _T_372; // @[PMP.scala 90:5:freechips.rocketchip.system.DefaultRV32Config.fir@176078.4]
  wire  _T_378; // @[PMP.scala 96:48:freechips.rocketchip.system.DefaultRV32Config.fir@176084.4]
  wire  _T_379; // @[PMP.scala 134:61:freechips.rocketchip.system.DefaultRV32Config.fir@176085.4]
  wire  _T_380; // @[PMP.scala 134:8:freechips.rocketchip.system.DefaultRV32Config.fir@176086.4]
  wire  _T_381; // @[PMP.scala 165:29:freechips.rocketchip.system.DefaultRV32Config.fir@176087.4]
  wire  _T_382; // @[PMP.scala 165:26:freechips.rocketchip.system.DefaultRV32Config.fir@176088.4]
  wire  _T_434; // @[PMP.scala 183:40:freechips.rocketchip.system.DefaultRV32Config.fir@176148.4]
  wire  _T_436; // @[PMP.scala 184:40:freechips.rocketchip.system.DefaultRV32Config.fir@176151.4]
  wire  _T_438; // @[PMP.scala 185:40:freechips.rocketchip.system.DefaultRV32Config.fir@176154.4]
  wire  _T_440_cfg_x; // @[PMP.scala 186:8:freechips.rocketchip.system.DefaultRV32Config.fir@176157.4]
  wire  _T_440_cfg_w; // @[PMP.scala 186:8:freechips.rocketchip.system.DefaultRV32Config.fir@176157.4]
  wire  _T_440_cfg_r; // @[PMP.scala 186:8:freechips.rocketchip.system.DefaultRV32Config.fir@176157.4]
  wire [31:0] _T_446; // @[PMP.scala 65:47:freechips.rocketchip.system.DefaultRV32Config.fir@176163.4]
  wire [31:0] _T_447; // @[PMP.scala 65:54:freechips.rocketchip.system.DefaultRV32Config.fir@176164.4]
  wire [31:0] _T_448; // @[PMP.scala 65:52:freechips.rocketchip.system.DefaultRV32Config.fir@176165.4]
  wire  _T_449; // @[PMP.scala 65:58:freechips.rocketchip.system.DefaultRV32Config.fir@176166.4]
  wire [31:0] _T_455; // @[PMP.scala 62:36:freechips.rocketchip.system.DefaultRV32Config.fir@176172.4]
  wire [31:0] _T_456; // @[PMP.scala 62:29:freechips.rocketchip.system.DefaultRV32Config.fir@176173.4]
  wire [31:0] _T_457; // @[PMP.scala 62:48:freechips.rocketchip.system.DefaultRV32Config.fir@176174.4]
  wire [31:0] _T_458; // @[PMP.scala 62:27:freechips.rocketchip.system.DefaultRV32Config.fir@176175.4]
  wire  _T_459; // @[PMP.scala 79:9:freechips.rocketchip.system.DefaultRV32Config.fir@176176.4]
  wire  _T_460; // @[PMP.scala 90:5:freechips.rocketchip.system.DefaultRV32Config.fir@176177.4]
  wire  _T_466; // @[PMP.scala 96:48:freechips.rocketchip.system.DefaultRV32Config.fir@176183.4]
  wire  _T_467; // @[PMP.scala 134:61:freechips.rocketchip.system.DefaultRV32Config.fir@176184.4]
  wire  _T_468; // @[PMP.scala 134:8:freechips.rocketchip.system.DefaultRV32Config.fir@176185.4]
  wire  _T_469; // @[PMP.scala 165:29:freechips.rocketchip.system.DefaultRV32Config.fir@176186.4]
  wire  _T_470; // @[PMP.scala 165:26:freechips.rocketchip.system.DefaultRV32Config.fir@176187.4]
  wire  _T_522; // @[PMP.scala 183:40:freechips.rocketchip.system.DefaultRV32Config.fir@176247.4]
  wire  _T_524; // @[PMP.scala 184:40:freechips.rocketchip.system.DefaultRV32Config.fir@176250.4]
  wire  _T_526; // @[PMP.scala 185:40:freechips.rocketchip.system.DefaultRV32Config.fir@176253.4]
  wire  _T_528_cfg_x; // @[PMP.scala 186:8:freechips.rocketchip.system.DefaultRV32Config.fir@176256.4]
  wire  _T_528_cfg_w; // @[PMP.scala 186:8:freechips.rocketchip.system.DefaultRV32Config.fir@176256.4]
  wire  _T_528_cfg_r; // @[PMP.scala 186:8:freechips.rocketchip.system.DefaultRV32Config.fir@176256.4]
  wire [31:0] _T_534; // @[PMP.scala 65:47:freechips.rocketchip.system.DefaultRV32Config.fir@176262.4]
  wire [31:0] _T_535; // @[PMP.scala 65:54:freechips.rocketchip.system.DefaultRV32Config.fir@176263.4]
  wire [31:0] _T_536; // @[PMP.scala 65:52:freechips.rocketchip.system.DefaultRV32Config.fir@176264.4]
  wire  _T_537; // @[PMP.scala 65:58:freechips.rocketchip.system.DefaultRV32Config.fir@176265.4]
  wire [31:0] _T_543; // @[PMP.scala 62:36:freechips.rocketchip.system.DefaultRV32Config.fir@176271.4]
  wire [31:0] _T_544; // @[PMP.scala 62:29:freechips.rocketchip.system.DefaultRV32Config.fir@176272.4]
  wire [31:0] _T_545; // @[PMP.scala 62:48:freechips.rocketchip.system.DefaultRV32Config.fir@176273.4]
  wire [31:0] _T_546; // @[PMP.scala 62:27:freechips.rocketchip.system.DefaultRV32Config.fir@176274.4]
  wire  _T_547; // @[PMP.scala 79:9:freechips.rocketchip.system.DefaultRV32Config.fir@176275.4]
  wire  _T_548; // @[PMP.scala 90:5:freechips.rocketchip.system.DefaultRV32Config.fir@176276.4]
  wire  _T_554; // @[PMP.scala 96:48:freechips.rocketchip.system.DefaultRV32Config.fir@176282.4]
  wire  _T_555; // @[PMP.scala 134:61:freechips.rocketchip.system.DefaultRV32Config.fir@176283.4]
  wire  _T_556; // @[PMP.scala 134:8:freechips.rocketchip.system.DefaultRV32Config.fir@176284.4]
  wire  _T_557; // @[PMP.scala 165:29:freechips.rocketchip.system.DefaultRV32Config.fir@176285.4]
  wire  _T_558; // @[PMP.scala 165:26:freechips.rocketchip.system.DefaultRV32Config.fir@176286.4]
  wire  _T_610; // @[PMP.scala 183:40:freechips.rocketchip.system.DefaultRV32Config.fir@176346.4]
  wire  _T_612; // @[PMP.scala 184:40:freechips.rocketchip.system.DefaultRV32Config.fir@176349.4]
  wire  _T_614; // @[PMP.scala 185:40:freechips.rocketchip.system.DefaultRV32Config.fir@176352.4]
  wire  _T_616_cfg_x; // @[PMP.scala 186:8:freechips.rocketchip.system.DefaultRV32Config.fir@176355.4]
  wire  _T_616_cfg_w; // @[PMP.scala 186:8:freechips.rocketchip.system.DefaultRV32Config.fir@176355.4]
  wire  _T_616_cfg_r; // @[PMP.scala 186:8:freechips.rocketchip.system.DefaultRV32Config.fir@176355.4]
  wire [31:0] _T_622; // @[PMP.scala 65:47:freechips.rocketchip.system.DefaultRV32Config.fir@176361.4]
  wire [31:0] _T_623; // @[PMP.scala 65:54:freechips.rocketchip.system.DefaultRV32Config.fir@176362.4]
  wire [31:0] _T_624; // @[PMP.scala 65:52:freechips.rocketchip.system.DefaultRV32Config.fir@176363.4]
  wire  _T_625; // @[PMP.scala 65:58:freechips.rocketchip.system.DefaultRV32Config.fir@176364.4]
  wire  _T_643; // @[PMP.scala 134:61:freechips.rocketchip.system.DefaultRV32Config.fir@176382.4]
  wire  _T_644; // @[PMP.scala 134:8:freechips.rocketchip.system.DefaultRV32Config.fir@176383.4]
  wire  _T_645; // @[PMP.scala 165:29:freechips.rocketchip.system.DefaultRV32Config.fir@176384.4]
  wire  _T_646; // @[PMP.scala 165:26:freechips.rocketchip.system.DefaultRV32Config.fir@176385.4]
  wire  _T_698; // @[PMP.scala 183:40:freechips.rocketchip.system.DefaultRV32Config.fir@176445.4]
  wire  _T_700; // @[PMP.scala 184:40:freechips.rocketchip.system.DefaultRV32Config.fir@176448.4]
  wire  _T_702; // @[PMP.scala 185:40:freechips.rocketchip.system.DefaultRV32Config.fir@176451.4]
  assign default_ = io_prv > 2'h1; // @[PMP.scala 157:56:freechips.rocketchip.system.DefaultRV32Config.fir@175641.4]
  assign _T_2 = {io_pmp_7_addr, 2'h0}; // @[PMP.scala 62:36:freechips.rocketchip.system.DefaultRV32Config.fir@175664.4]
  assign _T_3 = ~_T_2; // @[PMP.scala 62:29:freechips.rocketchip.system.DefaultRV32Config.fir@175665.4]
  assign _T_4 = _T_3 | 32'h3; // @[PMP.scala 62:48:freechips.rocketchip.system.DefaultRV32Config.fir@175666.4]
  assign _T_5 = ~_T_4; // @[PMP.scala 62:27:freechips.rocketchip.system.DefaultRV32Config.fir@175667.4]
  assign _T_6 = io_addr ^ _T_5; // @[PMP.scala 65:47:freechips.rocketchip.system.DefaultRV32Config.fir@175668.4]
  assign _T_7 = ~io_pmp_7_mask; // @[PMP.scala 65:54:freechips.rocketchip.system.DefaultRV32Config.fir@175669.4]
  assign _T_8 = _T_6 & _T_7; // @[PMP.scala 65:52:freechips.rocketchip.system.DefaultRV32Config.fir@175670.4]
  assign _T_9 = _T_8 == 32'h0; // @[PMP.scala 65:58:freechips.rocketchip.system.DefaultRV32Config.fir@175671.4]
  assign _T_15 = {io_pmp_6_addr, 2'h0}; // @[PMP.scala 62:36:freechips.rocketchip.system.DefaultRV32Config.fir@175677.4]
  assign _T_16 = ~_T_15; // @[PMP.scala 62:29:freechips.rocketchip.system.DefaultRV32Config.fir@175678.4]
  assign _T_17 = _T_16 | 32'h3; // @[PMP.scala 62:48:freechips.rocketchip.system.DefaultRV32Config.fir@175679.4]
  assign _T_18 = ~_T_17; // @[PMP.scala 62:27:freechips.rocketchip.system.DefaultRV32Config.fir@175680.4]
  assign _T_19 = io_addr < _T_18; // @[PMP.scala 79:9:freechips.rocketchip.system.DefaultRV32Config.fir@175681.4]
  assign _T_20 = ~_T_19; // @[PMP.scala 90:5:freechips.rocketchip.system.DefaultRV32Config.fir@175682.4]
  assign _T_25 = io_addr < _T_5; // @[PMP.scala 79:9:freechips.rocketchip.system.DefaultRV32Config.fir@175687.4]
  assign _T_26 = _T_20 & _T_25; // @[PMP.scala 96:48:freechips.rocketchip.system.DefaultRV32Config.fir@175688.4]
  assign _T_27 = io_pmp_7_cfg_a[0] & _T_26; // @[PMP.scala 134:61:freechips.rocketchip.system.DefaultRV32Config.fir@175689.4]
  assign _T_28 = io_pmp_7_cfg_a[1] ? _T_9 : _T_27; // @[PMP.scala 134:8:freechips.rocketchip.system.DefaultRV32Config.fir@175690.4]
  assign _T_29 = ~io_pmp_7_cfg_l; // @[PMP.scala 165:29:freechips.rocketchip.system.DefaultRV32Config.fir@175691.4]
  assign _T_30 = default_ & _T_29; // @[PMP.scala 165:26:freechips.rocketchip.system.DefaultRV32Config.fir@175692.4]
  assign _T_82 = io_pmp_7_cfg_r | _T_30; // @[PMP.scala 183:40:freechips.rocketchip.system.DefaultRV32Config.fir@175752.4]
  assign _T_84 = io_pmp_7_cfg_w | _T_30; // @[PMP.scala 184:40:freechips.rocketchip.system.DefaultRV32Config.fir@175755.4]
  assign _T_86 = io_pmp_7_cfg_x | _T_30; // @[PMP.scala 185:40:freechips.rocketchip.system.DefaultRV32Config.fir@175758.4]
  assign _T_88_cfg_x = _T_28 ? _T_86 : default_; // @[PMP.scala 186:8:freechips.rocketchip.system.DefaultRV32Config.fir@175761.4]
  assign _T_88_cfg_w = _T_28 ? _T_84 : default_; // @[PMP.scala 186:8:freechips.rocketchip.system.DefaultRV32Config.fir@175761.4]
  assign _T_88_cfg_r = _T_28 ? _T_82 : default_; // @[PMP.scala 186:8:freechips.rocketchip.system.DefaultRV32Config.fir@175761.4]
  assign _T_94 = io_addr ^ _T_18; // @[PMP.scala 65:47:freechips.rocketchip.system.DefaultRV32Config.fir@175767.4]
  assign _T_95 = ~io_pmp_6_mask; // @[PMP.scala 65:54:freechips.rocketchip.system.DefaultRV32Config.fir@175768.4]
  assign _T_96 = _T_94 & _T_95; // @[PMP.scala 65:52:freechips.rocketchip.system.DefaultRV32Config.fir@175769.4]
  assign _T_97 = _T_96 == 32'h0; // @[PMP.scala 65:58:freechips.rocketchip.system.DefaultRV32Config.fir@175770.4]
  assign _T_103 = {io_pmp_5_addr, 2'h0}; // @[PMP.scala 62:36:freechips.rocketchip.system.DefaultRV32Config.fir@175776.4]
  assign _T_104 = ~_T_103; // @[PMP.scala 62:29:freechips.rocketchip.system.DefaultRV32Config.fir@175777.4]
  assign _T_105 = _T_104 | 32'h3; // @[PMP.scala 62:48:freechips.rocketchip.system.DefaultRV32Config.fir@175778.4]
  assign _T_106 = ~_T_105; // @[PMP.scala 62:27:freechips.rocketchip.system.DefaultRV32Config.fir@175779.4]
  assign _T_107 = io_addr < _T_106; // @[PMP.scala 79:9:freechips.rocketchip.system.DefaultRV32Config.fir@175780.4]
  assign _T_108 = ~_T_107; // @[PMP.scala 90:5:freechips.rocketchip.system.DefaultRV32Config.fir@175781.4]
  assign _T_114 = _T_108 & _T_19; // @[PMP.scala 96:48:freechips.rocketchip.system.DefaultRV32Config.fir@175787.4]
  assign _T_115 = io_pmp_6_cfg_a[0] & _T_114; // @[PMP.scala 134:61:freechips.rocketchip.system.DefaultRV32Config.fir@175788.4]
  assign _T_116 = io_pmp_6_cfg_a[1] ? _T_97 : _T_115; // @[PMP.scala 134:8:freechips.rocketchip.system.DefaultRV32Config.fir@175789.4]
  assign _T_117 = ~io_pmp_6_cfg_l; // @[PMP.scala 165:29:freechips.rocketchip.system.DefaultRV32Config.fir@175790.4]
  assign _T_118 = default_ & _T_117; // @[PMP.scala 165:26:freechips.rocketchip.system.DefaultRV32Config.fir@175791.4]
  assign _T_170 = io_pmp_6_cfg_r | _T_118; // @[PMP.scala 183:40:freechips.rocketchip.system.DefaultRV32Config.fir@175851.4]
  assign _T_172 = io_pmp_6_cfg_w | _T_118; // @[PMP.scala 184:40:freechips.rocketchip.system.DefaultRV32Config.fir@175854.4]
  assign _T_174 = io_pmp_6_cfg_x | _T_118; // @[PMP.scala 185:40:freechips.rocketchip.system.DefaultRV32Config.fir@175857.4]
  assign _T_176_cfg_x = _T_116 ? _T_174 : _T_88_cfg_x; // @[PMP.scala 186:8:freechips.rocketchip.system.DefaultRV32Config.fir@175860.4]
  assign _T_176_cfg_w = _T_116 ? _T_172 : _T_88_cfg_w; // @[PMP.scala 186:8:freechips.rocketchip.system.DefaultRV32Config.fir@175860.4]
  assign _T_176_cfg_r = _T_116 ? _T_170 : _T_88_cfg_r; // @[PMP.scala 186:8:freechips.rocketchip.system.DefaultRV32Config.fir@175860.4]
  assign _T_182 = io_addr ^ _T_106; // @[PMP.scala 65:47:freechips.rocketchip.system.DefaultRV32Config.fir@175866.4]
  assign _T_183 = ~io_pmp_5_mask; // @[PMP.scala 65:54:freechips.rocketchip.system.DefaultRV32Config.fir@175867.4]
  assign _T_184 = _T_182 & _T_183; // @[PMP.scala 65:52:freechips.rocketchip.system.DefaultRV32Config.fir@175868.4]
  assign _T_185 = _T_184 == 32'h0; // @[PMP.scala 65:58:freechips.rocketchip.system.DefaultRV32Config.fir@175869.4]
  assign _T_191 = {io_pmp_4_addr, 2'h0}; // @[PMP.scala 62:36:freechips.rocketchip.system.DefaultRV32Config.fir@175875.4]
  assign _T_192 = ~_T_191; // @[PMP.scala 62:29:freechips.rocketchip.system.DefaultRV32Config.fir@175876.4]
  assign _T_193 = _T_192 | 32'h3; // @[PMP.scala 62:48:freechips.rocketchip.system.DefaultRV32Config.fir@175877.4]
  assign _T_194 = ~_T_193; // @[PMP.scala 62:27:freechips.rocketchip.system.DefaultRV32Config.fir@175878.4]
  assign _T_195 = io_addr < _T_194; // @[PMP.scala 79:9:freechips.rocketchip.system.DefaultRV32Config.fir@175879.4]
  assign _T_196 = ~_T_195; // @[PMP.scala 90:5:freechips.rocketchip.system.DefaultRV32Config.fir@175880.4]
  assign _T_202 = _T_196 & _T_107; // @[PMP.scala 96:48:freechips.rocketchip.system.DefaultRV32Config.fir@175886.4]
  assign _T_203 = io_pmp_5_cfg_a[0] & _T_202; // @[PMP.scala 134:61:freechips.rocketchip.system.DefaultRV32Config.fir@175887.4]
  assign _T_204 = io_pmp_5_cfg_a[1] ? _T_185 : _T_203; // @[PMP.scala 134:8:freechips.rocketchip.system.DefaultRV32Config.fir@175888.4]
  assign _T_205 = ~io_pmp_5_cfg_l; // @[PMP.scala 165:29:freechips.rocketchip.system.DefaultRV32Config.fir@175889.4]
  assign _T_206 = default_ & _T_205; // @[PMP.scala 165:26:freechips.rocketchip.system.DefaultRV32Config.fir@175890.4]
  assign _T_258 = io_pmp_5_cfg_r | _T_206; // @[PMP.scala 183:40:freechips.rocketchip.system.DefaultRV32Config.fir@175950.4]
  assign _T_260 = io_pmp_5_cfg_w | _T_206; // @[PMP.scala 184:40:freechips.rocketchip.system.DefaultRV32Config.fir@175953.4]
  assign _T_262 = io_pmp_5_cfg_x | _T_206; // @[PMP.scala 185:40:freechips.rocketchip.system.DefaultRV32Config.fir@175956.4]
  assign _T_264_cfg_x = _T_204 ? _T_262 : _T_176_cfg_x; // @[PMP.scala 186:8:freechips.rocketchip.system.DefaultRV32Config.fir@175959.4]
  assign _T_264_cfg_w = _T_204 ? _T_260 : _T_176_cfg_w; // @[PMP.scala 186:8:freechips.rocketchip.system.DefaultRV32Config.fir@175959.4]
  assign _T_264_cfg_r = _T_204 ? _T_258 : _T_176_cfg_r; // @[PMP.scala 186:8:freechips.rocketchip.system.DefaultRV32Config.fir@175959.4]
  assign _T_270 = io_addr ^ _T_194; // @[PMP.scala 65:47:freechips.rocketchip.system.DefaultRV32Config.fir@175965.4]
  assign _T_271 = ~io_pmp_4_mask; // @[PMP.scala 65:54:freechips.rocketchip.system.DefaultRV32Config.fir@175966.4]
  assign _T_272 = _T_270 & _T_271; // @[PMP.scala 65:52:freechips.rocketchip.system.DefaultRV32Config.fir@175967.4]
  assign _T_273 = _T_272 == 32'h0; // @[PMP.scala 65:58:freechips.rocketchip.system.DefaultRV32Config.fir@175968.4]
  assign _T_279 = {io_pmp_3_addr, 2'h0}; // @[PMP.scala 62:36:freechips.rocketchip.system.DefaultRV32Config.fir@175974.4]
  assign _T_280 = ~_T_279; // @[PMP.scala 62:29:freechips.rocketchip.system.DefaultRV32Config.fir@175975.4]
  assign _T_281 = _T_280 | 32'h3; // @[PMP.scala 62:48:freechips.rocketchip.system.DefaultRV32Config.fir@175976.4]
  assign _T_282 = ~_T_281; // @[PMP.scala 62:27:freechips.rocketchip.system.DefaultRV32Config.fir@175977.4]
  assign _T_283 = io_addr < _T_282; // @[PMP.scala 79:9:freechips.rocketchip.system.DefaultRV32Config.fir@175978.4]
  assign _T_284 = ~_T_283; // @[PMP.scala 90:5:freechips.rocketchip.system.DefaultRV32Config.fir@175979.4]
  assign _T_290 = _T_284 & _T_195; // @[PMP.scala 96:48:freechips.rocketchip.system.DefaultRV32Config.fir@175985.4]
  assign _T_291 = io_pmp_4_cfg_a[0] & _T_290; // @[PMP.scala 134:61:freechips.rocketchip.system.DefaultRV32Config.fir@175986.4]
  assign _T_292 = io_pmp_4_cfg_a[1] ? _T_273 : _T_291; // @[PMP.scala 134:8:freechips.rocketchip.system.DefaultRV32Config.fir@175987.4]
  assign _T_293 = ~io_pmp_4_cfg_l; // @[PMP.scala 165:29:freechips.rocketchip.system.DefaultRV32Config.fir@175988.4]
  assign _T_294 = default_ & _T_293; // @[PMP.scala 165:26:freechips.rocketchip.system.DefaultRV32Config.fir@175989.4]
  assign _T_346 = io_pmp_4_cfg_r | _T_294; // @[PMP.scala 183:40:freechips.rocketchip.system.DefaultRV32Config.fir@176049.4]
  assign _T_348 = io_pmp_4_cfg_w | _T_294; // @[PMP.scala 184:40:freechips.rocketchip.system.DefaultRV32Config.fir@176052.4]
  assign _T_350 = io_pmp_4_cfg_x | _T_294; // @[PMP.scala 185:40:freechips.rocketchip.system.DefaultRV32Config.fir@176055.4]
  assign _T_352_cfg_x = _T_292 ? _T_350 : _T_264_cfg_x; // @[PMP.scala 186:8:freechips.rocketchip.system.DefaultRV32Config.fir@176058.4]
  assign _T_352_cfg_w = _T_292 ? _T_348 : _T_264_cfg_w; // @[PMP.scala 186:8:freechips.rocketchip.system.DefaultRV32Config.fir@176058.4]
  assign _T_352_cfg_r = _T_292 ? _T_346 : _T_264_cfg_r; // @[PMP.scala 186:8:freechips.rocketchip.system.DefaultRV32Config.fir@176058.4]
  assign _T_358 = io_addr ^ _T_282; // @[PMP.scala 65:47:freechips.rocketchip.system.DefaultRV32Config.fir@176064.4]
  assign _T_359 = ~io_pmp_3_mask; // @[PMP.scala 65:54:freechips.rocketchip.system.DefaultRV32Config.fir@176065.4]
  assign _T_360 = _T_358 & _T_359; // @[PMP.scala 65:52:freechips.rocketchip.system.DefaultRV32Config.fir@176066.4]
  assign _T_361 = _T_360 == 32'h0; // @[PMP.scala 65:58:freechips.rocketchip.system.DefaultRV32Config.fir@176067.4]
  assign _T_367 = {io_pmp_2_addr, 2'h0}; // @[PMP.scala 62:36:freechips.rocketchip.system.DefaultRV32Config.fir@176073.4]
  assign _T_368 = ~_T_367; // @[PMP.scala 62:29:freechips.rocketchip.system.DefaultRV32Config.fir@176074.4]
  assign _T_369 = _T_368 | 32'h3; // @[PMP.scala 62:48:freechips.rocketchip.system.DefaultRV32Config.fir@176075.4]
  assign _T_370 = ~_T_369; // @[PMP.scala 62:27:freechips.rocketchip.system.DefaultRV32Config.fir@176076.4]
  assign _T_371 = io_addr < _T_370; // @[PMP.scala 79:9:freechips.rocketchip.system.DefaultRV32Config.fir@176077.4]
  assign _T_372 = ~_T_371; // @[PMP.scala 90:5:freechips.rocketchip.system.DefaultRV32Config.fir@176078.4]
  assign _T_378 = _T_372 & _T_283; // @[PMP.scala 96:48:freechips.rocketchip.system.DefaultRV32Config.fir@176084.4]
  assign _T_379 = io_pmp_3_cfg_a[0] & _T_378; // @[PMP.scala 134:61:freechips.rocketchip.system.DefaultRV32Config.fir@176085.4]
  assign _T_380 = io_pmp_3_cfg_a[1] ? _T_361 : _T_379; // @[PMP.scala 134:8:freechips.rocketchip.system.DefaultRV32Config.fir@176086.4]
  assign _T_381 = ~io_pmp_3_cfg_l; // @[PMP.scala 165:29:freechips.rocketchip.system.DefaultRV32Config.fir@176087.4]
  assign _T_382 = default_ & _T_381; // @[PMP.scala 165:26:freechips.rocketchip.system.DefaultRV32Config.fir@176088.4]
  assign _T_434 = io_pmp_3_cfg_r | _T_382; // @[PMP.scala 183:40:freechips.rocketchip.system.DefaultRV32Config.fir@176148.4]
  assign _T_436 = io_pmp_3_cfg_w | _T_382; // @[PMP.scala 184:40:freechips.rocketchip.system.DefaultRV32Config.fir@176151.4]
  assign _T_438 = io_pmp_3_cfg_x | _T_382; // @[PMP.scala 185:40:freechips.rocketchip.system.DefaultRV32Config.fir@176154.4]
  assign _T_440_cfg_x = _T_380 ? _T_438 : _T_352_cfg_x; // @[PMP.scala 186:8:freechips.rocketchip.system.DefaultRV32Config.fir@176157.4]
  assign _T_440_cfg_w = _T_380 ? _T_436 : _T_352_cfg_w; // @[PMP.scala 186:8:freechips.rocketchip.system.DefaultRV32Config.fir@176157.4]
  assign _T_440_cfg_r = _T_380 ? _T_434 : _T_352_cfg_r; // @[PMP.scala 186:8:freechips.rocketchip.system.DefaultRV32Config.fir@176157.4]
  assign _T_446 = io_addr ^ _T_370; // @[PMP.scala 65:47:freechips.rocketchip.system.DefaultRV32Config.fir@176163.4]
  assign _T_447 = ~io_pmp_2_mask; // @[PMP.scala 65:54:freechips.rocketchip.system.DefaultRV32Config.fir@176164.4]
  assign _T_448 = _T_446 & _T_447; // @[PMP.scala 65:52:freechips.rocketchip.system.DefaultRV32Config.fir@176165.4]
  assign _T_449 = _T_448 == 32'h0; // @[PMP.scala 65:58:freechips.rocketchip.system.DefaultRV32Config.fir@176166.4]
  assign _T_455 = {io_pmp_1_addr, 2'h0}; // @[PMP.scala 62:36:freechips.rocketchip.system.DefaultRV32Config.fir@176172.4]
  assign _T_456 = ~_T_455; // @[PMP.scala 62:29:freechips.rocketchip.system.DefaultRV32Config.fir@176173.4]
  assign _T_457 = _T_456 | 32'h3; // @[PMP.scala 62:48:freechips.rocketchip.system.DefaultRV32Config.fir@176174.4]
  assign _T_458 = ~_T_457; // @[PMP.scala 62:27:freechips.rocketchip.system.DefaultRV32Config.fir@176175.4]
  assign _T_459 = io_addr < _T_458; // @[PMP.scala 79:9:freechips.rocketchip.system.DefaultRV32Config.fir@176176.4]
  assign _T_460 = ~_T_459; // @[PMP.scala 90:5:freechips.rocketchip.system.DefaultRV32Config.fir@176177.4]
  assign _T_466 = _T_460 & _T_371; // @[PMP.scala 96:48:freechips.rocketchip.system.DefaultRV32Config.fir@176183.4]
  assign _T_467 = io_pmp_2_cfg_a[0] & _T_466; // @[PMP.scala 134:61:freechips.rocketchip.system.DefaultRV32Config.fir@176184.4]
  assign _T_468 = io_pmp_2_cfg_a[1] ? _T_449 : _T_467; // @[PMP.scala 134:8:freechips.rocketchip.system.DefaultRV32Config.fir@176185.4]
  assign _T_469 = ~io_pmp_2_cfg_l; // @[PMP.scala 165:29:freechips.rocketchip.system.DefaultRV32Config.fir@176186.4]
  assign _T_470 = default_ & _T_469; // @[PMP.scala 165:26:freechips.rocketchip.system.DefaultRV32Config.fir@176187.4]
  assign _T_522 = io_pmp_2_cfg_r | _T_470; // @[PMP.scala 183:40:freechips.rocketchip.system.DefaultRV32Config.fir@176247.4]
  assign _T_524 = io_pmp_2_cfg_w | _T_470; // @[PMP.scala 184:40:freechips.rocketchip.system.DefaultRV32Config.fir@176250.4]
  assign _T_526 = io_pmp_2_cfg_x | _T_470; // @[PMP.scala 185:40:freechips.rocketchip.system.DefaultRV32Config.fir@176253.4]
  assign _T_528_cfg_x = _T_468 ? _T_526 : _T_440_cfg_x; // @[PMP.scala 186:8:freechips.rocketchip.system.DefaultRV32Config.fir@176256.4]
  assign _T_528_cfg_w = _T_468 ? _T_524 : _T_440_cfg_w; // @[PMP.scala 186:8:freechips.rocketchip.system.DefaultRV32Config.fir@176256.4]
  assign _T_528_cfg_r = _T_468 ? _T_522 : _T_440_cfg_r; // @[PMP.scala 186:8:freechips.rocketchip.system.DefaultRV32Config.fir@176256.4]
  assign _T_534 = io_addr ^ _T_458; // @[PMP.scala 65:47:freechips.rocketchip.system.DefaultRV32Config.fir@176262.4]
  assign _T_535 = ~io_pmp_1_mask; // @[PMP.scala 65:54:freechips.rocketchip.system.DefaultRV32Config.fir@176263.4]
  assign _T_536 = _T_534 & _T_535; // @[PMP.scala 65:52:freechips.rocketchip.system.DefaultRV32Config.fir@176264.4]
  assign _T_537 = _T_536 == 32'h0; // @[PMP.scala 65:58:freechips.rocketchip.system.DefaultRV32Config.fir@176265.4]
  assign _T_543 = {io_pmp_0_addr, 2'h0}; // @[PMP.scala 62:36:freechips.rocketchip.system.DefaultRV32Config.fir@176271.4]
  assign _T_544 = ~_T_543; // @[PMP.scala 62:29:freechips.rocketchip.system.DefaultRV32Config.fir@176272.4]
  assign _T_545 = _T_544 | 32'h3; // @[PMP.scala 62:48:freechips.rocketchip.system.DefaultRV32Config.fir@176273.4]
  assign _T_546 = ~_T_545; // @[PMP.scala 62:27:freechips.rocketchip.system.DefaultRV32Config.fir@176274.4]
  assign _T_547 = io_addr < _T_546; // @[PMP.scala 79:9:freechips.rocketchip.system.DefaultRV32Config.fir@176275.4]
  assign _T_548 = ~_T_547; // @[PMP.scala 90:5:freechips.rocketchip.system.DefaultRV32Config.fir@176276.4]
  assign _T_554 = _T_548 & _T_459; // @[PMP.scala 96:48:freechips.rocketchip.system.DefaultRV32Config.fir@176282.4]
  assign _T_555 = io_pmp_1_cfg_a[0] & _T_554; // @[PMP.scala 134:61:freechips.rocketchip.system.DefaultRV32Config.fir@176283.4]
  assign _T_556 = io_pmp_1_cfg_a[1] ? _T_537 : _T_555; // @[PMP.scala 134:8:freechips.rocketchip.system.DefaultRV32Config.fir@176284.4]
  assign _T_557 = ~io_pmp_1_cfg_l; // @[PMP.scala 165:29:freechips.rocketchip.system.DefaultRV32Config.fir@176285.4]
  assign _T_558 = default_ & _T_557; // @[PMP.scala 165:26:freechips.rocketchip.system.DefaultRV32Config.fir@176286.4]
  assign _T_610 = io_pmp_1_cfg_r | _T_558; // @[PMP.scala 183:40:freechips.rocketchip.system.DefaultRV32Config.fir@176346.4]
  assign _T_612 = io_pmp_1_cfg_w | _T_558; // @[PMP.scala 184:40:freechips.rocketchip.system.DefaultRV32Config.fir@176349.4]
  assign _T_614 = io_pmp_1_cfg_x | _T_558; // @[PMP.scala 185:40:freechips.rocketchip.system.DefaultRV32Config.fir@176352.4]
  assign _T_616_cfg_x = _T_556 ? _T_614 : _T_528_cfg_x; // @[PMP.scala 186:8:freechips.rocketchip.system.DefaultRV32Config.fir@176355.4]
  assign _T_616_cfg_w = _T_556 ? _T_612 : _T_528_cfg_w; // @[PMP.scala 186:8:freechips.rocketchip.system.DefaultRV32Config.fir@176355.4]
  assign _T_616_cfg_r = _T_556 ? _T_610 : _T_528_cfg_r; // @[PMP.scala 186:8:freechips.rocketchip.system.DefaultRV32Config.fir@176355.4]
  assign _T_622 = io_addr ^ _T_546; // @[PMP.scala 65:47:freechips.rocketchip.system.DefaultRV32Config.fir@176361.4]
  assign _T_623 = ~io_pmp_0_mask; // @[PMP.scala 65:54:freechips.rocketchip.system.DefaultRV32Config.fir@176362.4]
  assign _T_624 = _T_622 & _T_623; // @[PMP.scala 65:52:freechips.rocketchip.system.DefaultRV32Config.fir@176363.4]
  assign _T_625 = _T_624 == 32'h0; // @[PMP.scala 65:58:freechips.rocketchip.system.DefaultRV32Config.fir@176364.4]
  assign _T_643 = io_pmp_0_cfg_a[0] & _T_547; // @[PMP.scala 134:61:freechips.rocketchip.system.DefaultRV32Config.fir@176382.4]
  assign _T_644 = io_pmp_0_cfg_a[1] ? _T_625 : _T_643; // @[PMP.scala 134:8:freechips.rocketchip.system.DefaultRV32Config.fir@176383.4]
  assign _T_645 = ~io_pmp_0_cfg_l; // @[PMP.scala 165:29:freechips.rocketchip.system.DefaultRV32Config.fir@176384.4]
  assign _T_646 = default_ & _T_645; // @[PMP.scala 165:26:freechips.rocketchip.system.DefaultRV32Config.fir@176385.4]
  assign _T_698 = io_pmp_0_cfg_r | _T_646; // @[PMP.scala 183:40:freechips.rocketchip.system.DefaultRV32Config.fir@176445.4]
  assign _T_700 = io_pmp_0_cfg_w | _T_646; // @[PMP.scala 184:40:freechips.rocketchip.system.DefaultRV32Config.fir@176448.4]
  assign _T_702 = io_pmp_0_cfg_x | _T_646; // @[PMP.scala 185:40:freechips.rocketchip.system.DefaultRV32Config.fir@176451.4]
  assign io_r = _T_644 ? _T_698 : _T_616_cfg_r; // @[PMP.scala 189:8:freechips.rocketchip.system.DefaultRV32Config.fir@176455.4]
  assign io_w = _T_644 ? _T_700 : _T_616_cfg_w; // @[PMP.scala 190:8:freechips.rocketchip.system.DefaultRV32Config.fir@176456.4]
  assign io_x = _T_644 ? _T_702 : _T_616_cfg_x; // @[PMP.scala 191:8:freechips.rocketchip.system.DefaultRV32Config.fir@176457.4]
endmodule
