module TLDebugModuleInner( // @[:freechips.rocketchip.system.DefaultRV32Config.fir@108907.2]
  input         clock, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@108908.4]
  input         reset, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@108909.4]
  output        auto_tl_in_a_ready, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@108910.4]
  input         auto_tl_in_a_valid, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@108910.4]
  input  [2:0]  auto_tl_in_a_bits_opcode, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@108910.4]
  input  [2:0]  auto_tl_in_a_bits_param, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@108910.4]
  input  [1:0]  auto_tl_in_a_bits_size, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@108910.4]
  input  [9:0]  auto_tl_in_a_bits_source, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@108910.4]
  input  [11:0] auto_tl_in_a_bits_address, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@108910.4]
  input  [3:0]  auto_tl_in_a_bits_mask, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@108910.4]
  input  [31:0] auto_tl_in_a_bits_data, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@108910.4]
  input         auto_tl_in_a_bits_corrupt, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@108910.4]
  input         auto_tl_in_d_ready, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@108910.4]
  output        auto_tl_in_d_valid, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@108910.4]
  output [2:0]  auto_tl_in_d_bits_opcode, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@108910.4]
  output [1:0]  auto_tl_in_d_bits_size, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@108910.4]
  output [9:0]  auto_tl_in_d_bits_source, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@108910.4]
  output [31:0] auto_tl_in_d_bits_data, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@108910.4]
  output        auto_dmi_in_a_ready, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@108910.4]
  input         auto_dmi_in_a_valid, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@108910.4]
  input  [2:0]  auto_dmi_in_a_bits_opcode, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@108910.4]
  input  [2:0]  auto_dmi_in_a_bits_param, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@108910.4]
  input  [1:0]  auto_dmi_in_a_bits_size, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@108910.4]
  input         auto_dmi_in_a_bits_source, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@108910.4]
  input  [8:0]  auto_dmi_in_a_bits_address, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@108910.4]
  input  [3:0]  auto_dmi_in_a_bits_mask, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@108910.4]
  input  [31:0] auto_dmi_in_a_bits_data, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@108910.4]
  input         auto_dmi_in_a_bits_corrupt, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@108910.4]
  input         auto_dmi_in_d_ready, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@108910.4]
  output        auto_dmi_in_d_valid, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@108910.4]
  output [2:0]  auto_dmi_in_d_bits_opcode, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@108910.4]
  output [1:0]  auto_dmi_in_d_bits_size, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@108910.4]
  output        auto_dmi_in_d_bits_source, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@108910.4]
  output [31:0] auto_dmi_in_d_bits_data, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@108910.4]
  input         io_dmactive, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@108911.4]
  output        io_innerCtrl_ready, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@108911.4]
  input         io_innerCtrl_valid, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@108911.4]
  input         io_innerCtrl_bits_resumereq, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@108911.4]
  input  [9:0]  io_innerCtrl_bits_hartsel, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@108911.4]
  input         io_innerCtrl_bits_ackhavereset, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@108911.4]
  input         io_innerCtrl_bits_hrmask_0, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@108911.4]
  output        io_hgDebugInt_0, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@108911.4]
  input         io_hartIsInReset_0 // @[:freechips.rocketchip.system.DefaultRV32Config.fir@108911.4]
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [31:0] _RAND_34;
  reg [31:0] _RAND_35;
  reg [31:0] _RAND_36;
  reg [31:0] _RAND_37;
  reg [31:0] _RAND_38;
  reg [31:0] _RAND_39;
  reg [31:0] _RAND_40;
  reg [31:0] _RAND_41;
  reg [31:0] _RAND_42;
  reg [31:0] _RAND_43;
  reg [31:0] _RAND_44;
  reg [31:0] _RAND_45;
  reg [31:0] _RAND_46;
  reg [31:0] _RAND_47;
  reg [31:0] _RAND_48;
  reg [31:0] _RAND_49;
  reg [31:0] _RAND_50;
  reg [31:0] _RAND_51;
  reg [31:0] _RAND_52;
  reg [31:0] _RAND_53;
  reg [31:0] _RAND_54;
  reg [31:0] _RAND_55;
  reg [31:0] _RAND_56;
  reg [31:0] _RAND_57;
  reg [31:0] _RAND_58;
  reg [31:0] _RAND_59;
  reg [31:0] _RAND_60;
  reg [31:0] _RAND_61;
  reg [31:0] _RAND_62;
  reg [31:0] _RAND_63;
  reg [31:0] _RAND_64;
  reg [31:0] _RAND_65;
  reg [31:0] _RAND_66;
  reg [31:0] _RAND_67;
  reg [31:0] _RAND_68;
  reg [31:0] _RAND_69;
  reg [31:0] _RAND_70;
  reg [31:0] _RAND_71;
  reg [31:0] _RAND_72;
  reg [31:0] _RAND_73;
  reg [31:0] _RAND_74;
  reg [31:0] _RAND_75;
  reg [31:0] _RAND_76;
  reg [31:0] _RAND_77;
  reg [31:0] _RAND_78;
  reg [31:0] _RAND_79;
  reg [31:0] _RAND_80;
  reg [31:0] _RAND_81;
`endif // RANDOMIZE_REG_INIT
  wire  TLMonitor_clock; // @[Nodes.scala 25:25:freechips.rocketchip.system.DefaultRV32Config.fir@108919.4]
  wire  TLMonitor_reset; // @[Nodes.scala 25:25:freechips.rocketchip.system.DefaultRV32Config.fir@108919.4]
  wire  TLMonitor_io_in_a_ready; // @[Nodes.scala 25:25:freechips.rocketchip.system.DefaultRV32Config.fir@108919.4]
  wire  TLMonitor_io_in_a_valid; // @[Nodes.scala 25:25:freechips.rocketchip.system.DefaultRV32Config.fir@108919.4]
  wire [2:0] TLMonitor_io_in_a_bits_opcode; // @[Nodes.scala 25:25:freechips.rocketchip.system.DefaultRV32Config.fir@108919.4]
  wire [2:0] TLMonitor_io_in_a_bits_param; // @[Nodes.scala 25:25:freechips.rocketchip.system.DefaultRV32Config.fir@108919.4]
  wire [1:0] TLMonitor_io_in_a_bits_size; // @[Nodes.scala 25:25:freechips.rocketchip.system.DefaultRV32Config.fir@108919.4]
  wire  TLMonitor_io_in_a_bits_source; // @[Nodes.scala 25:25:freechips.rocketchip.system.DefaultRV32Config.fir@108919.4]
  wire [8:0] TLMonitor_io_in_a_bits_address; // @[Nodes.scala 25:25:freechips.rocketchip.system.DefaultRV32Config.fir@108919.4]
  wire [3:0] TLMonitor_io_in_a_bits_mask; // @[Nodes.scala 25:25:freechips.rocketchip.system.DefaultRV32Config.fir@108919.4]
  wire  TLMonitor_io_in_a_bits_corrupt; // @[Nodes.scala 25:25:freechips.rocketchip.system.DefaultRV32Config.fir@108919.4]
  wire  TLMonitor_io_in_d_ready; // @[Nodes.scala 25:25:freechips.rocketchip.system.DefaultRV32Config.fir@108919.4]
  wire  TLMonitor_io_in_d_valid; // @[Nodes.scala 25:25:freechips.rocketchip.system.DefaultRV32Config.fir@108919.4]
  wire [2:0] TLMonitor_io_in_d_bits_opcode; // @[Nodes.scala 25:25:freechips.rocketchip.system.DefaultRV32Config.fir@108919.4]
  wire [1:0] TLMonitor_io_in_d_bits_size; // @[Nodes.scala 25:25:freechips.rocketchip.system.DefaultRV32Config.fir@108919.4]
  wire  TLMonitor_io_in_d_bits_source; // @[Nodes.scala 25:25:freechips.rocketchip.system.DefaultRV32Config.fir@108919.4]
  wire  TLMonitor_1_clock; // @[Nodes.scala 25:25:freechips.rocketchip.system.DefaultRV32Config.fir@108944.4]
  wire  TLMonitor_1_reset; // @[Nodes.scala 25:25:freechips.rocketchip.system.DefaultRV32Config.fir@108944.4]
  wire  TLMonitor_1_io_in_a_ready; // @[Nodes.scala 25:25:freechips.rocketchip.system.DefaultRV32Config.fir@108944.4]
  wire  TLMonitor_1_io_in_a_valid; // @[Nodes.scala 25:25:freechips.rocketchip.system.DefaultRV32Config.fir@108944.4]
  wire [2:0] TLMonitor_1_io_in_a_bits_opcode; // @[Nodes.scala 25:25:freechips.rocketchip.system.DefaultRV32Config.fir@108944.4]
  wire [2:0] TLMonitor_1_io_in_a_bits_param; // @[Nodes.scala 25:25:freechips.rocketchip.system.DefaultRV32Config.fir@108944.4]
  wire [1:0] TLMonitor_1_io_in_a_bits_size; // @[Nodes.scala 25:25:freechips.rocketchip.system.DefaultRV32Config.fir@108944.4]
  wire [9:0] TLMonitor_1_io_in_a_bits_source; // @[Nodes.scala 25:25:freechips.rocketchip.system.DefaultRV32Config.fir@108944.4]
  wire [11:0] TLMonitor_1_io_in_a_bits_address; // @[Nodes.scala 25:25:freechips.rocketchip.system.DefaultRV32Config.fir@108944.4]
  wire [3:0] TLMonitor_1_io_in_a_bits_mask; // @[Nodes.scala 25:25:freechips.rocketchip.system.DefaultRV32Config.fir@108944.4]
  wire  TLMonitor_1_io_in_a_bits_corrupt; // @[Nodes.scala 25:25:freechips.rocketchip.system.DefaultRV32Config.fir@108944.4]
  wire  TLMonitor_1_io_in_d_ready; // @[Nodes.scala 25:25:freechips.rocketchip.system.DefaultRV32Config.fir@108944.4]
  wire  TLMonitor_1_io_in_d_valid; // @[Nodes.scala 25:25:freechips.rocketchip.system.DefaultRV32Config.fir@108944.4]
  wire [2:0] TLMonitor_1_io_in_d_bits_opcode; // @[Nodes.scala 25:25:freechips.rocketchip.system.DefaultRV32Config.fir@108944.4]
  wire [1:0] TLMonitor_1_io_in_d_bits_size; // @[Nodes.scala 25:25:freechips.rocketchip.system.DefaultRV32Config.fir@108944.4]
  wire [9:0] TLMonitor_1_io_in_d_bits_source; // @[Nodes.scala 25:25:freechips.rocketchip.system.DefaultRV32Config.fir@108944.4]
  wire  debug_hartReset_0_clock; // @[ShiftReg.scala 45:23:freechips.rocketchip.system.DefaultRV32Config.fir@109292.4]
  wire  debug_hartReset_0_reset; // @[ShiftReg.scala 45:23:freechips.rocketchip.system.DefaultRV32Config.fir@109292.4]
  wire  debug_hartReset_0_io_d; // @[ShiftReg.scala 45:23:freechips.rocketchip.system.DefaultRV32Config.fir@109292.4]
  wire  debug_hartReset_0_io_q; // @[ShiftReg.scala 45:23:freechips.rocketchip.system.DefaultRV32Config.fir@109292.4]
  reg  haltedBitRegs_0; // @[Debug.scala 757:31:freechips.rocketchip.system.DefaultRV32Config.fir@108972.4]
  reg  resumeReqRegs_0; // @[Debug.scala 758:31:freechips.rocketchip.system.DefaultRV32Config.fir@108973.4]
  reg  haveResetBitRegs_0; // @[Debug.scala 759:31:freechips.rocketchip.system.DefaultRV32Config.fir@108974.4]
  wire  hamaskWrSel_0; // @[Debug.scala 820:61:freechips.rocketchip.system.DefaultRV32Config.fir@109282.4]
  reg  hrmaskReg_0; // @[Debug.scala 832:29:freechips.rocketchip.system.DefaultRV32Config.fir@109290.4]
  wire  _T_13; // @[Debug.scala 839:11:freechips.rocketchip.system.DefaultRV32Config.fir@109299.4]
  wire  _T_16; // @[Decoupled.scala 40:37:freechips.rocketchip.system.DefaultRV32Config.fir@109306.6]
  reg  hrDebugInt_0; // @[Debug.scala 846:34:freechips.rocketchip.system.DefaultRV32Config.fir@109313.4]
  wire  _T_23; // @[package.scala 62:38:freechips.rocketchip.system.DefaultRV32Config.fir@109321.6]
  wire  _T_24; // @[package.scala 57:72:freechips.rocketchip.system.DefaultRV32Config.fir@109322.6]
  wire  hartIsInResetSync_0; // @[ShiftReg.scala 48:24:freechips.rocketchip.system.DefaultRV32Config.fir@109296.4 ShiftReg.scala 48:24:freechips.rocketchip.system.DefaultRV32Config.fir@109297.4]
  wire  _T_25; // @[package.scala 58:75:freechips.rocketchip.system.DefaultRV32Config.fir@109323.6]
  wire  _T_26; // @[package.scala 57:72:freechips.rocketchip.system.DefaultRV32Config.fir@109324.6]
  wire  resumereq; // @[Debug.scala 868:41:freechips.rocketchip.system.DefaultRV32Config.fir@109373.4]
  wire  _T_306; // @[Debug.scala 1227:32:freechips.rocketchip.system.DefaultRV32Config.fir@110286.4]
  wire  _T_307; // @[Debug.scala 1227:73:freechips.rocketchip.system.DefaultRV32Config.fir@110287.4]
  wire  _T_308; // @[Debug.scala 1227:61:freechips.rocketchip.system.DefaultRV32Config.fir@110288.4]
  wire  resumeAcks_0; // @[Debug.scala 1227:58:freechips.rocketchip.system.DefaultRV32Config.fir@110289.4]
  wire  _T_64; // @[Debug.scala 902:39:freechips.rocketchip.system.DefaultRV32Config.fir@109438.8]
  wire  _T_65; // @[Debug.scala 902:73:freechips.rocketchip.system.DefaultRV32Config.fir@109439.8]
  wire  _GEN_34; // @[Debug.scala 902:100:freechips.rocketchip.system.DefaultRV32Config.fir@109440.8]
  wire  _GEN_35; // @[Debug.scala 900:49:freechips.rocketchip.system.DefaultRV32Config.fir@109433.6]
  wire [31:0] haltedStatus_0; // @[Debug.scala 1051:30:freechips.rocketchip.system.DefaultRV32Config.fir@109501.4 Debug.scala 1055:26:freechips.rocketchip.system.DefaultRV32Config.fir@109503.6 Debug.scala 1057:26:freechips.rocketchip.system.DefaultRV32Config.fir@109506.6]
  wire  haltedSummary; // @[Debug.scala 1061:48:freechips.rocketchip.system.DefaultRV32Config.fir@109508.4]
  wire [31:0] HALTSUM1RdData_haltsum1; // @[:freechips.rocketchip.system.DefaultRV32Config.fir@109510.4 :freechips.rocketchip.system.DefaultRV32Config.fir@109511.4]
  reg [2:0] ABSTRACTCSReg_cmderr; // @[Debug.scala 1075:34:freechips.rocketchip.system.DefaultRV32Config.fir@109543.4]
  wire  _T_380; // @[RegisterRouter.scala 69:36:freechips.rocketchip.system.DefaultRV32Config.fir@110366.4]
  wire [4:0] _T_2990; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@113342.4]
  wire [6:0] _T_385; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@110382.4]
  wire  _T_433; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@110430.4]
  wire  _T_389; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@110386.4]
  wire  _T_407; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@110404.4]
  wire  _T_3564; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@114522.4]
  wire  _T_3565; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@114523.4]
  wire  _T_3566; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@114524.4]
  wire [31:0] _T_3035; // @[OneHot.scala 58:35:freechips.rocketchip.system.DefaultRV32Config.fir@113387.4]
  wire  _T_3598; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@114599.4]
  wire  _T_3599; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@114600.4]
  wire [7:0] _T_465; // @[Bitwise.scala 72:12:freechips.rocketchip.system.DefaultRV32Config.fir@110466.4]
  wire [7:0] _T_463; // @[Bitwise.scala 72:12:freechips.rocketchip.system.DefaultRV32Config.fir@110464.4]
  wire [7:0] _T_461; // @[Bitwise.scala 72:12:freechips.rocketchip.system.DefaultRV32Config.fir@110462.4]
  wire [7:0] _T_459; // @[Bitwise.scala 72:12:freechips.rocketchip.system.DefaultRV32Config.fir@110460.4]
  wire [31:0] _T_468; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@110469.4]
  wire  _T_1929; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@112114.4]
  wire  ABSTRACTCSWrEnMaybe; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@112118.4]
  reg [1:0] ctrlStateReg; // @[Debug.scala 1559:27:freechips.rocketchip.system.DefaultRV32Config.fir@168657.4]
  wire  ABSTRACTCSWrEnLegal; // @[Debug.scala 1569:44:freechips.rocketchip.system.DefaultRV32Config.fir@168662.4]
  wire  ABSTRACTCSWrEn; // @[Debug.scala 1083:51:freechips.rocketchip.system.DefaultRV32Config.fir@109577.4]
  wire [2:0] ABSTRACTCSWrData_cmderr; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@112119.4]
  wire [2:0] _T_83; // @[Debug.scala 1103:58:freechips.rocketchip.system.DefaultRV32Config.fir@109617.16]
  wire [2:0] _T_84; // @[Debug.scala 1103:56:freechips.rocketchip.system.DefaultRV32Config.fir@109618.16]
  wire  _T_44818; // @[Debug.scala 1623:30:freechips.rocketchip.system.DefaultRV32Config.fir@168740.6]
  reg [7:0] COMMANDRdData_cmdtype; // @[Debug.scala 1160:25:freechips.rocketchip.system.DefaultRV32Config.fir@110144.4]
  wire  commandRegIsAccessRegister; // @[Debug.scala 1584:58:freechips.rocketchip.system.DefaultRV32Config.fir@168691.4]
  reg [23:0] COMMANDRdData_control; // @[Debug.scala 1160:25:freechips.rocketchip.system.DefaultRV32Config.fir@110144.4]
  wire [31:0] _T_3960; // @[Debug.scala 1415:62:freechips.rocketchip.system.DefaultRV32Config.fir@115544.4]
  wire  accessRegisterCommandReg_transfer; // @[Debug.scala 1415:73:freechips.rocketchip.system.DefaultRV32Config.fir@115552.4]
  wire  accessRegisterCommandReg_write; // @[Debug.scala 1415:73:freechips.rocketchip.system.DefaultRV32Config.fir@115550.4]
  wire  _T_44808; // @[Debug.scala 1602:19:freechips.rocketchip.system.DefaultRV32Config.fir@168709.8]
  wire [15:0] accessRegisterCommandReg_regno; // @[Debug.scala 1415:73:freechips.rocketchip.system.DefaultRV32Config.fir@115548.4]
  wire  _T_44803; // @[Debug.scala 1592:58:freechips.rocketchip.system.DefaultRV32Config.fir@168698.4]
  wire  _T_44804; // @[Debug.scala 1592:104:freechips.rocketchip.system.DefaultRV32Config.fir@168699.4]
  wire  accessRegIsGPR; // @[Debug.scala 1592:70:freechips.rocketchip.system.DefaultRV32Config.fir@168700.4]
  wire  _T_44809; // @[Debug.scala 1602:54:freechips.rocketchip.system.DefaultRV32Config.fir@168710.8]
  wire  _GEN_3623; // @[Debug.scala 1602:73:freechips.rocketchip.system.DefaultRV32Config.fir@168711.8]
  wire  commandRegIsUnsupported; // @[Debug.scala 1599:39:freechips.rocketchip.system.DefaultRV32Config.fir@168701.4]
  wire  _GEN_3624; // @[Debug.scala 1602:73:freechips.rocketchip.system.DefaultRV32Config.fir@168711.8]
  wire  commandRegBadHaltResume; // @[Debug.scala 1599:39:freechips.rocketchip.system.DefaultRV32Config.fir@168701.4]
  wire  _GEN_3640; // @[Debug.scala 1630:38:freechips.rocketchip.system.DefaultRV32Config.fir@168742.8]
  wire  _GEN_3653; // @[Debug.scala 1623:59:freechips.rocketchip.system.DefaultRV32Config.fir@168741.6]
  wire  errorHaltResume; // @[Debug.scala 1615:47:freechips.rocketchip.system.DefaultRV32Config.fir@168724.4]
  wire  _T_3603; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@114613.4]
  wire  _T_3604; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@114614.4]
  wire  _T_2649; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@112936.4]
  wire  COMMANDWrEnMaybe; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@112940.4]
  wire  COMMANDWrEn; // @[Debug.scala 1168:40:freechips.rocketchip.system.DefaultRV32Config.fir@110163.4]
  wire [31:0] COMMANDWrDataVal; // @[Debug.scala 265:24:freechips.rocketchip.system.DefaultRV32Config.fir@112944.4]
  wire [7:0] COMMANDWrData_cmdtype; // @[Debug.scala 1163:65:freechips.rocketchip.system.DefaultRV32Config.fir@110152.4]
  wire  commandWrIsAccessRegister; // @[Debug.scala 1583:60:freechips.rocketchip.system.DefaultRV32Config.fir@168690.4]
  wire  _T_44811; // @[Debug.scala 1608:48:freechips.rocketchip.system.DefaultRV32Config.fir@168717.4]
  wire  _T_44812; // @[Debug.scala 1608:103:freechips.rocketchip.system.DefaultRV32Config.fir@168718.4]
  wire  wrAccessRegisterCommand; // @[Debug.scala 1608:78:freechips.rocketchip.system.DefaultRV32Config.fir@168719.4]
  wire  _T_3588; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@114581.4]
  wire  _T_3589; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@114582.4]
  wire  _T_2791; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@113103.4]
  wire  dmiAbstractDataWrEnMaybe_0; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@113107.4]
  wire  _T_3400; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@114156.4]
  wire  _T_3422; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@114213.4]
  wire  _T_3423; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@114214.4]
  wire  _T_2789; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@113101.4]
  wire  dmiAbstractDataRdEn_0; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@113105.4]
  wire  dmiAbstractDataAccessVec_0; // @[Debug.scala 1141:105:freechips.rocketchip.system.DefaultRV32Config.fir@109690.4]
  reg [11:0] ABSTRACTAUTOReg_autoexecdata; // @[Debug.scala 1119:36:freechips.rocketchip.system.DefaultRV32Config.fir@109639.4]
  wire  autoexecData_0; // @[Debug.scala 1152:140:freechips.rocketchip.system.DefaultRV32Config.fir@110072.4]
  wire  _T_3648; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@114680.4]
  wire  _T_3649; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@114681.4]
  wire  dmiProgramBufferWrEnMaybe_0; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@111264.4]
  wire  _T_3482; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@114312.4]
  wire  _T_3483; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@114313.4]
  wire  dmiProgramBufferRdEn_0; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@111262.4]
  wire  dmiProgramBufferAccessVec_0; // @[Debug.scala 1144:108:freechips.rocketchip.system.DefaultRV32Config.fir@109828.4]
  reg [15:0] ABSTRACTAUTOReg_autoexecprogbuf; // @[Debug.scala 1119:36:freechips.rocketchip.system.DefaultRV32Config.fir@109639.4]
  wire  autoexecProg_0; // @[Debug.scala 1153:144:freechips.rocketchip.system.DefaultRV32Config.fir@110090.4]
  wire  _T_3653; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@114691.4]
  wire  _T_3654; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@114692.4]
  wire  dmiProgramBufferWrEnMaybe_4; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@111028.4]
  wire  _T_3487; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@114323.4]
  wire  _T_3488; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@114324.4]
  wire  dmiProgramBufferRdEn_4; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@111026.4]
  wire  dmiProgramBufferAccessVec_4; // @[Debug.scala 1144:108:freechips.rocketchip.system.DefaultRV32Config.fir@109832.4]
  wire  autoexecProg_1; // @[Debug.scala 1153:144:freechips.rocketchip.system.DefaultRV32Config.fir@110092.4]
  wire  _T_276; // @[Debug.scala 1155:73:freechips.rocketchip.system.DefaultRV32Config.fir@110122.4]
  wire  _T_3658; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@114702.4]
  wire  _T_3659; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@114703.4]
  wire  dmiProgramBufferWrEnMaybe_8; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@111382.4]
  wire  _T_3492; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@114334.4]
  wire  _T_3493; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@114335.4]
  wire  dmiProgramBufferRdEn_8; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@111380.4]
  wire  dmiProgramBufferAccessVec_8; // @[Debug.scala 1144:108:freechips.rocketchip.system.DefaultRV32Config.fir@109836.4]
  wire  autoexecProg_2; // @[Debug.scala 1153:144:freechips.rocketchip.system.DefaultRV32Config.fir@110094.4]
  wire  _T_277; // @[Debug.scala 1155:73:freechips.rocketchip.system.DefaultRV32Config.fir@110123.4]
  wire  _T_3663; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@114713.4]
  wire  _T_3664; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@114714.4]
  wire  dmiProgramBufferWrEnMaybe_12; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@112473.4]
  wire  _T_3497; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@114345.4]
  wire  _T_3498; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@114346.4]
  wire  dmiProgramBufferRdEn_12; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@112471.4]
  wire  dmiProgramBufferAccessVec_12; // @[Debug.scala 1144:108:freechips.rocketchip.system.DefaultRV32Config.fir@109840.4]
  wire  autoexecProg_3; // @[Debug.scala 1153:144:freechips.rocketchip.system.DefaultRV32Config.fir@110096.4]
  wire  _T_278; // @[Debug.scala 1155:73:freechips.rocketchip.system.DefaultRV32Config.fir@110124.4]
  wire  _T_3668; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@114724.4]
  wire  _T_3669; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@114725.4]
  wire  dmiProgramBufferWrEnMaybe_16; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@112968.4]
  wire  _T_3502; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@114356.4]
  wire  _T_3503; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@114357.4]
  wire  dmiProgramBufferRdEn_16; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@112966.4]
  wire  dmiProgramBufferAccessVec_16; // @[Debug.scala 1144:108:freechips.rocketchip.system.DefaultRV32Config.fir@109844.4]
  wire  autoexecProg_4; // @[Debug.scala 1153:144:freechips.rocketchip.system.DefaultRV32Config.fir@110098.4]
  wire  _T_279; // @[Debug.scala 1155:73:freechips.rocketchip.system.DefaultRV32Config.fir@110125.4]
  wire  _T_3673; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@114735.4]
  wire  _T_3674; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@114736.4]
  wire  dmiProgramBufferWrEnMaybe_20; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@110674.4]
  wire  _T_3507; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@114367.4]
  wire  _T_3508; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@114368.4]
  wire  dmiProgramBufferRdEn_20; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@110672.4]
  wire  dmiProgramBufferAccessVec_20; // @[Debug.scala 1144:108:freechips.rocketchip.system.DefaultRV32Config.fir@109848.4]
  wire  autoexecProg_5; // @[Debug.scala 1153:144:freechips.rocketchip.system.DefaultRV32Config.fir@110100.4]
  wire  _T_280; // @[Debug.scala 1155:73:freechips.rocketchip.system.DefaultRV32Config.fir@110126.4]
  wire  _T_3678; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@114746.4]
  wire  _T_3679; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@114747.4]
  wire  dmiProgramBufferWrEnMaybe_24; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@110910.4]
  wire  _T_3512; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@114378.4]
  wire  _T_3513; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@114379.4]
  wire  dmiProgramBufferRdEn_24; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@110908.4]
  wire  dmiProgramBufferAccessVec_24; // @[Debug.scala 1144:108:freechips.rocketchip.system.DefaultRV32Config.fir@109852.4]
  wire  autoexecProg_6; // @[Debug.scala 1153:144:freechips.rocketchip.system.DefaultRV32Config.fir@110102.4]
  wire  _T_281; // @[Debug.scala 1155:73:freechips.rocketchip.system.DefaultRV32Config.fir@110127.4]
  wire  _T_3683; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@114757.4]
  wire  _T_3684; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@114758.4]
  wire  dmiProgramBufferWrEnMaybe_28; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@112355.4]
  wire  _T_3517; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@114389.4]
  wire  _T_3518; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@114390.4]
  wire  dmiProgramBufferRdEn_28; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@112353.4]
  wire  dmiProgramBufferAccessVec_28; // @[Debug.scala 1144:108:freechips.rocketchip.system.DefaultRV32Config.fir@109856.4]
  wire  autoexecProg_7; // @[Debug.scala 1153:144:freechips.rocketchip.system.DefaultRV32Config.fir@110104.4]
  wire  _T_282; // @[Debug.scala 1155:73:freechips.rocketchip.system.DefaultRV32Config.fir@110128.4]
  wire  _T_3688; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@114768.4]
  wire  _T_3689; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@114769.4]
  wire  dmiProgramBufferWrEnMaybe_32; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@112822.4]
  wire  _T_3522; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@114400.4]
  wire  _T_3523; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@114401.4]
  wire  dmiProgramBufferRdEn_32; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@112820.4]
  wire  dmiProgramBufferAccessVec_32; // @[Debug.scala 1144:108:freechips.rocketchip.system.DefaultRV32Config.fir@109860.4]
  wire  autoexecProg_8; // @[Debug.scala 1153:144:freechips.rocketchip.system.DefaultRV32Config.fir@110106.4]
  wire  _T_283; // @[Debug.scala 1155:73:freechips.rocketchip.system.DefaultRV32Config.fir@110129.4]
  wire  _T_3693; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@114779.4]
  wire  _T_3694; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@114780.4]
  wire  dmiProgramBufferWrEnMaybe_36; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@111146.4]
  wire  _T_3527; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@114411.4]
  wire  _T_3528; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@114412.4]
  wire  dmiProgramBufferRdEn_36; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@111144.4]
  wire  dmiProgramBufferAccessVec_36; // @[Debug.scala 1144:108:freechips.rocketchip.system.DefaultRV32Config.fir@109864.4]
  wire  autoexecProg_9; // @[Debug.scala 1153:144:freechips.rocketchip.system.DefaultRV32Config.fir@110108.4]
  wire  _T_284; // @[Debug.scala 1155:73:freechips.rocketchip.system.DefaultRV32Config.fir@110130.4]
  wire  _T_3698; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@114790.4]
  wire  _T_3699; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@114791.4]
  wire  dmiProgramBufferWrEnMaybe_40; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@110481.4]
  wire  _T_3532; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@114422.4]
  wire  _T_3533; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@114423.4]
  wire  dmiProgramBufferRdEn_40; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@110479.4]
  wire  dmiProgramBufferAccessVec_40; // @[Debug.scala 1144:108:freechips.rocketchip.system.DefaultRV32Config.fir@109868.4]
  wire  autoexecProg_10; // @[Debug.scala 1153:144:freechips.rocketchip.system.DefaultRV32Config.fir@110110.4]
  wire  _T_285; // @[Debug.scala 1155:73:freechips.rocketchip.system.DefaultRV32Config.fir@110131.4]
  wire  _T_3703; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@114801.4]
  wire  _T_3704; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@114802.4]
  wire  dmiProgramBufferWrEnMaybe_44; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@112704.4]
  wire  _T_3537; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@114433.4]
  wire  _T_3538; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@114434.4]
  wire  dmiProgramBufferRdEn_44; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@112702.4]
  wire  dmiProgramBufferAccessVec_44; // @[Debug.scala 1144:108:freechips.rocketchip.system.DefaultRV32Config.fir@109872.4]
  wire  autoexecProg_11; // @[Debug.scala 1153:144:freechips.rocketchip.system.DefaultRV32Config.fir@110112.4]
  wire  _T_286; // @[Debug.scala 1155:73:freechips.rocketchip.system.DefaultRV32Config.fir@110132.4]
  wire  _T_3708; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@114812.4]
  wire  _T_3709; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@114813.4]
  wire  dmiProgramBufferWrEnMaybe_48; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@112237.4]
  wire  _T_3542; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@114444.4]
  wire  _T_3543; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@114445.4]
  wire  dmiProgramBufferRdEn_48; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@112235.4]
  wire  dmiProgramBufferAccessVec_48; // @[Debug.scala 1144:108:freechips.rocketchip.system.DefaultRV32Config.fir@109876.4]
  wire  autoexecProg_12; // @[Debug.scala 1153:144:freechips.rocketchip.system.DefaultRV32Config.fir@110114.4]
  wire  _T_287; // @[Debug.scala 1155:73:freechips.rocketchip.system.DefaultRV32Config.fir@110133.4]
  wire  _T_3713; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@114823.4]
  wire  _T_3714; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@114824.4]
  wire  dmiProgramBufferWrEnMaybe_52; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@111500.4]
  wire  _T_3547; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@114455.4]
  wire  _T_3548; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@114456.4]
  wire  dmiProgramBufferRdEn_52; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@111498.4]
  wire  dmiProgramBufferAccessVec_52; // @[Debug.scala 1144:108:freechips.rocketchip.system.DefaultRV32Config.fir@109880.4]
  wire  autoexecProg_13; // @[Debug.scala 1153:144:freechips.rocketchip.system.DefaultRV32Config.fir@110116.4]
  wire  _T_288; // @[Debug.scala 1155:73:freechips.rocketchip.system.DefaultRV32Config.fir@110134.4]
  wire  _T_3718; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@114834.4]
  wire  _T_3719; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@114835.4]
  wire  dmiProgramBufferWrEnMaybe_56; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@110792.4]
  wire  _T_3552; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@114466.4]
  wire  _T_3553; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@114467.4]
  wire  dmiProgramBufferRdEn_56; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@110790.4]
  wire  dmiProgramBufferAccessVec_56; // @[Debug.scala 1144:108:freechips.rocketchip.system.DefaultRV32Config.fir@109884.4]
  wire  autoexecProg_14; // @[Debug.scala 1153:144:freechips.rocketchip.system.DefaultRV32Config.fir@110118.4]
  wire  _T_289; // @[Debug.scala 1155:73:freechips.rocketchip.system.DefaultRV32Config.fir@110135.4]
  wire  _T_3723; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@114845.4]
  wire  _T_3724; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@114846.4]
  wire  dmiProgramBufferWrEnMaybe_60; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@113225.4]
  wire  _T_3557; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@114477.4]
  wire  _T_3558; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@114478.4]
  wire  dmiProgramBufferRdEn_60; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@113223.4]
  wire  dmiProgramBufferAccessVec_60; // @[Debug.scala 1144:108:freechips.rocketchip.system.DefaultRV32Config.fir@109888.4]
  wire  autoexecProg_15; // @[Debug.scala 1153:144:freechips.rocketchip.system.DefaultRV32Config.fir@110120.4]
  wire  _T_290; // @[Debug.scala 1155:73:freechips.rocketchip.system.DefaultRV32Config.fir@110136.4]
  wire  autoexec; // @[Debug.scala 1155:48:freechips.rocketchip.system.DefaultRV32Config.fir@110137.4]
  wire  _T_44813; // @[Debug.scala 1609:48:freechips.rocketchip.system.DefaultRV32Config.fir@168720.4]
  wire  regAccessRegisterCommand; // @[Debug.scala 1609:78:freechips.rocketchip.system.DefaultRV32Config.fir@168722.4]
  wire  _T_44816; // @[Debug.scala 1616:37:freechips.rocketchip.system.DefaultRV32Config.fir@168725.6]
  wire  _T_44802; // @[Debug.scala 1586:49:freechips.rocketchip.system.DefaultRV32Config.fir@168692.4]
  wire  commandWrIsUnsupported; // @[Debug.scala 1586:46:freechips.rocketchip.system.DefaultRV32Config.fir@168693.4]
  wire  _T_44817; // @[Debug.scala 1620:28:freechips.rocketchip.system.DefaultRV32Config.fir@168734.10]
  wire  _GEN_3630; // @[Debug.scala 1618:43:freechips.rocketchip.system.DefaultRV32Config.fir@168730.8]
  wire  _GEN_3632; // @[Debug.scala 1616:66:freechips.rocketchip.system.DefaultRV32Config.fir@168726.6]
  wire  _GEN_3651; // @[Debug.scala 1623:59:freechips.rocketchip.system.DefaultRV32Config.fir@168741.6]
  wire  errorUnsupported; // @[Debug.scala 1615:47:freechips.rocketchip.system.DefaultRV32Config.fir@168724.4]
  wire  _T_44819; // @[Debug.scala 1644:30:freechips.rocketchip.system.DefaultRV32Config.fir@168762.8]
  wire  _T_6050; // @[RegisterRouter.scala 69:36:freechips.rocketchip.system.DefaultRV32Config.fir@117696.4]
  wire [8:0] _T_33453; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@145326.4]
  wire [9:0] _T_6055; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@117712.4]
  wire  _T_6089; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@117746.4]
  wire  _T_6609; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@118266.4]
  wire  _T_42194; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@162227.4]
  wire  _T_42195; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@162228.4]
  wire  _T_42196; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@162229.4]
  wire [511:0] _T_33985; // @[OneHot.scala 58:35:freechips.rocketchip.system.DefaultRV32Config.fir@145858.4]
  wire  _T_42533; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@162788.4]
  wire  _T_42534; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@162789.4]
  wire [7:0] _T_6689; // @[Bitwise.scala 72:12:freechips.rocketchip.system.DefaultRV32Config.fir@118350.4]
  wire [7:0] _T_6687; // @[Bitwise.scala 72:12:freechips.rocketchip.system.DefaultRV32Config.fir@118348.4]
  wire [7:0] _T_6685; // @[Bitwise.scala 72:12:freechips.rocketchip.system.DefaultRV32Config.fir@118346.4]
  wire [7:0] _T_6683; // @[Bitwise.scala 72:12:freechips.rocketchip.system.DefaultRV32Config.fir@118344.4]
  wire [31:0] _T_6692; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@118353.4]
  wire  _T_25711; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@137522.4]
  wire  hartExceptionWrEn; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@137526.4]
  wire  _GEN_3649; // @[Debug.scala 1644:51:freechips.rocketchip.system.DefaultRV32Config.fir@168763.8]
  wire  _GEN_3655; // @[Debug.scala 1623:59:freechips.rocketchip.system.DefaultRV32Config.fir@168741.6]
  wire  errorException; // @[Debug.scala 1615:47:freechips.rocketchip.system.DefaultRV32Config.fir@168724.4]
  wire  _T_44785; // @[Debug.scala 1575:45:freechips.rocketchip.system.DefaultRV32Config.fir@168672.4]
  wire  _T_44786; // @[Debug.scala 1575:42:freechips.rocketchip.system.DefaultRV32Config.fir@168673.4]
  wire  _T_3608; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@114621.4]
  wire  _T_3609; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@114622.4]
  wire  _T_574; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@110595.4]
  wire  autoexecdataWrEnMaybe; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@110599.4]
  wire  _T_44788; // @[Debug.scala 1576:42:freechips.rocketchip.system.DefaultRV32Config.fir@168675.4]
  wire  _T_44789; // @[Debug.scala 1575:74:freechips.rocketchip.system.DefaultRV32Config.fir@168676.4]
  wire  _T_620; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@110643.4]
  wire  autoexecprogbufWrEnMaybe; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@110647.4]
  wire  _T_44791; // @[Debug.scala 1577:44:freechips.rocketchip.system.DefaultRV32Config.fir@168678.4]
  wire  _T_44792; // @[Debug.scala 1576:74:freechips.rocketchip.system.DefaultRV32Config.fir@168679.4]
  wire  _T_44794; // @[Debug.scala 1578:42:freechips.rocketchip.system.DefaultRV32Config.fir@168681.4]
  wire  _T_44795; // @[Debug.scala 1577:74:freechips.rocketchip.system.DefaultRV32Config.fir@168682.4]
  wire  _T_2814; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@113131.4]
  wire  dmiAbstractDataWrEnMaybe_1; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@113135.4]
  wire  _T_2812; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@113129.4]
  wire  dmiAbstractDataRdEn_1; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@113133.4]
  wire  dmiAbstractDataAccessVec_1; // @[Debug.scala 1141:105:freechips.rocketchip.system.DefaultRV32Config.fir@109691.4]
  wire  _T_165; // @[Debug.scala 1146:68:freechips.rocketchip.system.DefaultRV32Config.fir@109956.4]
  wire  _T_2839; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@113161.4]
  wire  dmiAbstractDataWrEnMaybe_2; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@113165.4]
  wire  _T_2837; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@113159.4]
  wire  dmiAbstractDataRdEn_2; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@113163.4]
  wire  dmiAbstractDataAccessVec_2; // @[Debug.scala 1141:105:freechips.rocketchip.system.DefaultRV32Config.fir@109692.4]
  wire  _T_166; // @[Debug.scala 1146:68:freechips.rocketchip.system.DefaultRV32Config.fir@109957.4]
  wire  _T_2864; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@113191.4]
  wire  dmiAbstractDataWrEnMaybe_3; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@113195.4]
  wire  _T_2862; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@113189.4]
  wire  dmiAbstractDataRdEn_3; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@113193.4]
  wire  dmiAbstractDataAccessVec_3; // @[Debug.scala 1141:105:freechips.rocketchip.system.DefaultRV32Config.fir@109693.4]
  wire  dmiAbstractDataAccess; // @[Debug.scala 1146:68:freechips.rocketchip.system.DefaultRV32Config.fir@109958.4]
  wire  _T_44797; // @[Debug.scala 1579:42:freechips.rocketchip.system.DefaultRV32Config.fir@168684.4]
  wire  _T_44798; // @[Debug.scala 1578:74:freechips.rocketchip.system.DefaultRV32Config.fir@168685.4]
  wire  dmiProgramBufferWrEnMaybe_1; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@111292.4]
  wire  dmiProgramBufferRdEn_1; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@111290.4]
  wire  dmiProgramBufferAccessVec_1; // @[Debug.scala 1144:108:freechips.rocketchip.system.DefaultRV32Config.fir@109829.4]
  wire  _T_167; // @[Debug.scala 1147:69:freechips.rocketchip.system.DefaultRV32Config.fir@109959.4]
  wire  dmiProgramBufferWrEnMaybe_2; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@111322.4]
  wire  dmiProgramBufferRdEn_2; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@111320.4]
  wire  dmiProgramBufferAccessVec_2; // @[Debug.scala 1144:108:freechips.rocketchip.system.DefaultRV32Config.fir@109830.4]
  wire  _T_168; // @[Debug.scala 1147:69:freechips.rocketchip.system.DefaultRV32Config.fir@109960.4]
  wire  dmiProgramBufferWrEnMaybe_3; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@111352.4]
  wire  dmiProgramBufferRdEn_3; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@111350.4]
  wire  dmiProgramBufferAccessVec_3; // @[Debug.scala 1144:108:freechips.rocketchip.system.DefaultRV32Config.fir@109831.4]
  wire  _T_169; // @[Debug.scala 1147:69:freechips.rocketchip.system.DefaultRV32Config.fir@109961.4]
  wire  _T_170; // @[Debug.scala 1147:69:freechips.rocketchip.system.DefaultRV32Config.fir@109962.4]
  wire  dmiProgramBufferWrEnMaybe_5; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@111056.4]
  wire  dmiProgramBufferRdEn_5; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@111054.4]
  wire  dmiProgramBufferAccessVec_5; // @[Debug.scala 1144:108:freechips.rocketchip.system.DefaultRV32Config.fir@109833.4]
  wire  _T_171; // @[Debug.scala 1147:69:freechips.rocketchip.system.DefaultRV32Config.fir@109963.4]
  wire  dmiProgramBufferWrEnMaybe_6; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@111086.4]
  wire  dmiProgramBufferRdEn_6; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@111084.4]
  wire  dmiProgramBufferAccessVec_6; // @[Debug.scala 1144:108:freechips.rocketchip.system.DefaultRV32Config.fir@109834.4]
  wire  _T_172; // @[Debug.scala 1147:69:freechips.rocketchip.system.DefaultRV32Config.fir@109964.4]
  wire  dmiProgramBufferWrEnMaybe_7; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@111116.4]
  wire  dmiProgramBufferRdEn_7; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@111114.4]
  wire  dmiProgramBufferAccessVec_7; // @[Debug.scala 1144:108:freechips.rocketchip.system.DefaultRV32Config.fir@109835.4]
  wire  _T_173; // @[Debug.scala 1147:69:freechips.rocketchip.system.DefaultRV32Config.fir@109965.4]
  wire  _T_174; // @[Debug.scala 1147:69:freechips.rocketchip.system.DefaultRV32Config.fir@109966.4]
  wire  dmiProgramBufferWrEnMaybe_9; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@111410.4]
  wire  dmiProgramBufferRdEn_9; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@111408.4]
  wire  dmiProgramBufferAccessVec_9; // @[Debug.scala 1144:108:freechips.rocketchip.system.DefaultRV32Config.fir@109837.4]
  wire  _T_175; // @[Debug.scala 1147:69:freechips.rocketchip.system.DefaultRV32Config.fir@109967.4]
  wire  dmiProgramBufferWrEnMaybe_10; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@111440.4]
  wire  dmiProgramBufferRdEn_10; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@111438.4]
  wire  dmiProgramBufferAccessVec_10; // @[Debug.scala 1144:108:freechips.rocketchip.system.DefaultRV32Config.fir@109838.4]
  wire  _T_176; // @[Debug.scala 1147:69:freechips.rocketchip.system.DefaultRV32Config.fir@109968.4]
  wire  dmiProgramBufferWrEnMaybe_11; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@111470.4]
  wire  dmiProgramBufferRdEn_11; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@111468.4]
  wire  dmiProgramBufferAccessVec_11; // @[Debug.scala 1144:108:freechips.rocketchip.system.DefaultRV32Config.fir@109839.4]
  wire  _T_177; // @[Debug.scala 1147:69:freechips.rocketchip.system.DefaultRV32Config.fir@109969.4]
  wire  _T_178; // @[Debug.scala 1147:69:freechips.rocketchip.system.DefaultRV32Config.fir@109970.4]
  wire  dmiProgramBufferWrEnMaybe_13; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@112501.4]
  wire  dmiProgramBufferRdEn_13; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@112499.4]
  wire  dmiProgramBufferAccessVec_13; // @[Debug.scala 1144:108:freechips.rocketchip.system.DefaultRV32Config.fir@109841.4]
  wire  _T_179; // @[Debug.scala 1147:69:freechips.rocketchip.system.DefaultRV32Config.fir@109971.4]
  wire  dmiProgramBufferWrEnMaybe_14; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@112531.4]
  wire  dmiProgramBufferRdEn_14; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@112529.4]
  wire  dmiProgramBufferAccessVec_14; // @[Debug.scala 1144:108:freechips.rocketchip.system.DefaultRV32Config.fir@109842.4]
  wire  _T_180; // @[Debug.scala 1147:69:freechips.rocketchip.system.DefaultRV32Config.fir@109972.4]
  wire  dmiProgramBufferWrEnMaybe_15; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@112561.4]
  wire  dmiProgramBufferRdEn_15; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@112559.4]
  wire  dmiProgramBufferAccessVec_15; // @[Debug.scala 1144:108:freechips.rocketchip.system.DefaultRV32Config.fir@109843.4]
  wire  _T_181; // @[Debug.scala 1147:69:freechips.rocketchip.system.DefaultRV32Config.fir@109973.4]
  wire  _T_182; // @[Debug.scala 1147:69:freechips.rocketchip.system.DefaultRV32Config.fir@109974.4]
  wire  dmiProgramBufferWrEnMaybe_17; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@112996.4]
  wire  dmiProgramBufferRdEn_17; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@112994.4]
  wire  dmiProgramBufferAccessVec_17; // @[Debug.scala 1144:108:freechips.rocketchip.system.DefaultRV32Config.fir@109845.4]
  wire  _T_183; // @[Debug.scala 1147:69:freechips.rocketchip.system.DefaultRV32Config.fir@109975.4]
  wire  dmiProgramBufferWrEnMaybe_18; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@113026.4]
  wire  dmiProgramBufferRdEn_18; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@113024.4]
  wire  dmiProgramBufferAccessVec_18; // @[Debug.scala 1144:108:freechips.rocketchip.system.DefaultRV32Config.fir@109846.4]
  wire  _T_184; // @[Debug.scala 1147:69:freechips.rocketchip.system.DefaultRV32Config.fir@109976.4]
  wire  dmiProgramBufferWrEnMaybe_19; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@113056.4]
  wire  dmiProgramBufferRdEn_19; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@113054.4]
  wire  dmiProgramBufferAccessVec_19; // @[Debug.scala 1144:108:freechips.rocketchip.system.DefaultRV32Config.fir@109847.4]
  wire  _T_185; // @[Debug.scala 1147:69:freechips.rocketchip.system.DefaultRV32Config.fir@109977.4]
  wire  _T_186; // @[Debug.scala 1147:69:freechips.rocketchip.system.DefaultRV32Config.fir@109978.4]
  wire  dmiProgramBufferWrEnMaybe_21; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@110702.4]
  wire  dmiProgramBufferRdEn_21; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@110700.4]
  wire  dmiProgramBufferAccessVec_21; // @[Debug.scala 1144:108:freechips.rocketchip.system.DefaultRV32Config.fir@109849.4]
  wire  _T_187; // @[Debug.scala 1147:69:freechips.rocketchip.system.DefaultRV32Config.fir@109979.4]
  wire  dmiProgramBufferWrEnMaybe_22; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@110732.4]
  wire  dmiProgramBufferRdEn_22; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@110730.4]
  wire  dmiProgramBufferAccessVec_22; // @[Debug.scala 1144:108:freechips.rocketchip.system.DefaultRV32Config.fir@109850.4]
  wire  _T_188; // @[Debug.scala 1147:69:freechips.rocketchip.system.DefaultRV32Config.fir@109980.4]
  wire  dmiProgramBufferWrEnMaybe_23; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@110762.4]
  wire  dmiProgramBufferRdEn_23; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@110760.4]
  wire  dmiProgramBufferAccessVec_23; // @[Debug.scala 1144:108:freechips.rocketchip.system.DefaultRV32Config.fir@109851.4]
  wire  _T_189; // @[Debug.scala 1147:69:freechips.rocketchip.system.DefaultRV32Config.fir@109981.4]
  wire  _T_190; // @[Debug.scala 1147:69:freechips.rocketchip.system.DefaultRV32Config.fir@109982.4]
  wire  dmiProgramBufferWrEnMaybe_25; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@110938.4]
  wire  dmiProgramBufferRdEn_25; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@110936.4]
  wire  dmiProgramBufferAccessVec_25; // @[Debug.scala 1144:108:freechips.rocketchip.system.DefaultRV32Config.fir@109853.4]
  wire  _T_191; // @[Debug.scala 1147:69:freechips.rocketchip.system.DefaultRV32Config.fir@109983.4]
  wire  dmiProgramBufferWrEnMaybe_26; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@110968.4]
  wire  dmiProgramBufferRdEn_26; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@110966.4]
  wire  dmiProgramBufferAccessVec_26; // @[Debug.scala 1144:108:freechips.rocketchip.system.DefaultRV32Config.fir@109854.4]
  wire  _T_192; // @[Debug.scala 1147:69:freechips.rocketchip.system.DefaultRV32Config.fir@109984.4]
  wire  dmiProgramBufferWrEnMaybe_27; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@110998.4]
  wire  dmiProgramBufferRdEn_27; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@110996.4]
  wire  dmiProgramBufferAccessVec_27; // @[Debug.scala 1144:108:freechips.rocketchip.system.DefaultRV32Config.fir@109855.4]
  wire  _T_193; // @[Debug.scala 1147:69:freechips.rocketchip.system.DefaultRV32Config.fir@109985.4]
  wire  _T_194; // @[Debug.scala 1147:69:freechips.rocketchip.system.DefaultRV32Config.fir@109986.4]
  wire  dmiProgramBufferWrEnMaybe_29; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@112383.4]
  wire  dmiProgramBufferRdEn_29; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@112381.4]
  wire  dmiProgramBufferAccessVec_29; // @[Debug.scala 1144:108:freechips.rocketchip.system.DefaultRV32Config.fir@109857.4]
  wire  _T_195; // @[Debug.scala 1147:69:freechips.rocketchip.system.DefaultRV32Config.fir@109987.4]
  wire  dmiProgramBufferWrEnMaybe_30; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@112413.4]
  wire  dmiProgramBufferRdEn_30; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@112411.4]
  wire  dmiProgramBufferAccessVec_30; // @[Debug.scala 1144:108:freechips.rocketchip.system.DefaultRV32Config.fir@109858.4]
  wire  _T_196; // @[Debug.scala 1147:69:freechips.rocketchip.system.DefaultRV32Config.fir@109988.4]
  wire  dmiProgramBufferWrEnMaybe_31; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@112443.4]
  wire  dmiProgramBufferRdEn_31; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@112441.4]
  wire  dmiProgramBufferAccessVec_31; // @[Debug.scala 1144:108:freechips.rocketchip.system.DefaultRV32Config.fir@109859.4]
  wire  _T_197; // @[Debug.scala 1147:69:freechips.rocketchip.system.DefaultRV32Config.fir@109989.4]
  wire  _T_198; // @[Debug.scala 1147:69:freechips.rocketchip.system.DefaultRV32Config.fir@109990.4]
  wire  dmiProgramBufferWrEnMaybe_33; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@112850.4]
  wire  dmiProgramBufferRdEn_33; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@112848.4]
  wire  dmiProgramBufferAccessVec_33; // @[Debug.scala 1144:108:freechips.rocketchip.system.DefaultRV32Config.fir@109861.4]
  wire  _T_199; // @[Debug.scala 1147:69:freechips.rocketchip.system.DefaultRV32Config.fir@109991.4]
  wire  dmiProgramBufferWrEnMaybe_34; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@112880.4]
  wire  dmiProgramBufferRdEn_34; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@112878.4]
  wire  dmiProgramBufferAccessVec_34; // @[Debug.scala 1144:108:freechips.rocketchip.system.DefaultRV32Config.fir@109862.4]
  wire  _T_200; // @[Debug.scala 1147:69:freechips.rocketchip.system.DefaultRV32Config.fir@109992.4]
  wire  dmiProgramBufferWrEnMaybe_35; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@112910.4]
  wire  dmiProgramBufferRdEn_35; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@112908.4]
  wire  dmiProgramBufferAccessVec_35; // @[Debug.scala 1144:108:freechips.rocketchip.system.DefaultRV32Config.fir@109863.4]
  wire  _T_201; // @[Debug.scala 1147:69:freechips.rocketchip.system.DefaultRV32Config.fir@109993.4]
  wire  _T_202; // @[Debug.scala 1147:69:freechips.rocketchip.system.DefaultRV32Config.fir@109994.4]
  wire  dmiProgramBufferWrEnMaybe_37; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@111174.4]
  wire  dmiProgramBufferRdEn_37; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@111172.4]
  wire  dmiProgramBufferAccessVec_37; // @[Debug.scala 1144:108:freechips.rocketchip.system.DefaultRV32Config.fir@109865.4]
  wire  _T_203; // @[Debug.scala 1147:69:freechips.rocketchip.system.DefaultRV32Config.fir@109995.4]
  wire  dmiProgramBufferWrEnMaybe_38; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@111204.4]
  wire  dmiProgramBufferRdEn_38; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@111202.4]
  wire  dmiProgramBufferAccessVec_38; // @[Debug.scala 1144:108:freechips.rocketchip.system.DefaultRV32Config.fir@109866.4]
  wire  _T_204; // @[Debug.scala 1147:69:freechips.rocketchip.system.DefaultRV32Config.fir@109996.4]
  wire  dmiProgramBufferWrEnMaybe_39; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@111234.4]
  wire  dmiProgramBufferRdEn_39; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@111232.4]
  wire  dmiProgramBufferAccessVec_39; // @[Debug.scala 1144:108:freechips.rocketchip.system.DefaultRV32Config.fir@109867.4]
  wire  _T_205; // @[Debug.scala 1147:69:freechips.rocketchip.system.DefaultRV32Config.fir@109997.4]
  wire  _T_206; // @[Debug.scala 1147:69:freechips.rocketchip.system.DefaultRV32Config.fir@109998.4]
  wire  dmiProgramBufferWrEnMaybe_41; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@110509.4]
  wire  dmiProgramBufferRdEn_41; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@110507.4]
  wire  dmiProgramBufferAccessVec_41; // @[Debug.scala 1144:108:freechips.rocketchip.system.DefaultRV32Config.fir@109869.4]
  wire  _T_207; // @[Debug.scala 1147:69:freechips.rocketchip.system.DefaultRV32Config.fir@109999.4]
  wire  dmiProgramBufferWrEnMaybe_42; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@110539.4]
  wire  dmiProgramBufferRdEn_42; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@110537.4]
  wire  dmiProgramBufferAccessVec_42; // @[Debug.scala 1144:108:freechips.rocketchip.system.DefaultRV32Config.fir@109870.4]
  wire  _T_208; // @[Debug.scala 1147:69:freechips.rocketchip.system.DefaultRV32Config.fir@110000.4]
  wire  dmiProgramBufferWrEnMaybe_43; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@110569.4]
  wire  dmiProgramBufferRdEn_43; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@110567.4]
  wire  dmiProgramBufferAccessVec_43; // @[Debug.scala 1144:108:freechips.rocketchip.system.DefaultRV32Config.fir@109871.4]
  wire  _T_209; // @[Debug.scala 1147:69:freechips.rocketchip.system.DefaultRV32Config.fir@110001.4]
  wire  _T_210; // @[Debug.scala 1147:69:freechips.rocketchip.system.DefaultRV32Config.fir@110002.4]
  wire  dmiProgramBufferWrEnMaybe_45; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@112732.4]
  wire  dmiProgramBufferRdEn_45; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@112730.4]
  wire  dmiProgramBufferAccessVec_45; // @[Debug.scala 1144:108:freechips.rocketchip.system.DefaultRV32Config.fir@109873.4]
  wire  _T_211; // @[Debug.scala 1147:69:freechips.rocketchip.system.DefaultRV32Config.fir@110003.4]
  wire  dmiProgramBufferWrEnMaybe_46; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@112762.4]
  wire  dmiProgramBufferRdEn_46; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@112760.4]
  wire  dmiProgramBufferAccessVec_46; // @[Debug.scala 1144:108:freechips.rocketchip.system.DefaultRV32Config.fir@109874.4]
  wire  _T_212; // @[Debug.scala 1147:69:freechips.rocketchip.system.DefaultRV32Config.fir@110004.4]
  wire  dmiProgramBufferWrEnMaybe_47; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@112792.4]
  wire  dmiProgramBufferRdEn_47; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@112790.4]
  wire  dmiProgramBufferAccessVec_47; // @[Debug.scala 1144:108:freechips.rocketchip.system.DefaultRV32Config.fir@109875.4]
  wire  _T_213; // @[Debug.scala 1147:69:freechips.rocketchip.system.DefaultRV32Config.fir@110005.4]
  wire  _T_214; // @[Debug.scala 1147:69:freechips.rocketchip.system.DefaultRV32Config.fir@110006.4]
  wire  dmiProgramBufferWrEnMaybe_49; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@112265.4]
  wire  dmiProgramBufferRdEn_49; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@112263.4]
  wire  dmiProgramBufferAccessVec_49; // @[Debug.scala 1144:108:freechips.rocketchip.system.DefaultRV32Config.fir@109877.4]
  wire  _T_215; // @[Debug.scala 1147:69:freechips.rocketchip.system.DefaultRV32Config.fir@110007.4]
  wire  dmiProgramBufferWrEnMaybe_50; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@112295.4]
  wire  dmiProgramBufferRdEn_50; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@112293.4]
  wire  dmiProgramBufferAccessVec_50; // @[Debug.scala 1144:108:freechips.rocketchip.system.DefaultRV32Config.fir@109878.4]
  wire  _T_216; // @[Debug.scala 1147:69:freechips.rocketchip.system.DefaultRV32Config.fir@110008.4]
  wire  dmiProgramBufferWrEnMaybe_51; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@112325.4]
  wire  dmiProgramBufferRdEn_51; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@112323.4]
  wire  dmiProgramBufferAccessVec_51; // @[Debug.scala 1144:108:freechips.rocketchip.system.DefaultRV32Config.fir@109879.4]
  wire  _T_217; // @[Debug.scala 1147:69:freechips.rocketchip.system.DefaultRV32Config.fir@110009.4]
  wire  _T_218; // @[Debug.scala 1147:69:freechips.rocketchip.system.DefaultRV32Config.fir@110010.4]
  wire  dmiProgramBufferWrEnMaybe_53; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@111528.4]
  wire  dmiProgramBufferRdEn_53; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@111526.4]
  wire  dmiProgramBufferAccessVec_53; // @[Debug.scala 1144:108:freechips.rocketchip.system.DefaultRV32Config.fir@109881.4]
  wire  _T_219; // @[Debug.scala 1147:69:freechips.rocketchip.system.DefaultRV32Config.fir@110011.4]
  wire  dmiProgramBufferWrEnMaybe_54; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@111558.4]
  wire  dmiProgramBufferRdEn_54; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@111556.4]
  wire  dmiProgramBufferAccessVec_54; // @[Debug.scala 1144:108:freechips.rocketchip.system.DefaultRV32Config.fir@109882.4]
  wire  _T_220; // @[Debug.scala 1147:69:freechips.rocketchip.system.DefaultRV32Config.fir@110012.4]
  wire  dmiProgramBufferWrEnMaybe_55; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@111588.4]
  wire  dmiProgramBufferRdEn_55; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@111586.4]
  wire  dmiProgramBufferAccessVec_55; // @[Debug.scala 1144:108:freechips.rocketchip.system.DefaultRV32Config.fir@109883.4]
  wire  _T_221; // @[Debug.scala 1147:69:freechips.rocketchip.system.DefaultRV32Config.fir@110013.4]
  wire  _T_222; // @[Debug.scala 1147:69:freechips.rocketchip.system.DefaultRV32Config.fir@110014.4]
  wire  dmiProgramBufferWrEnMaybe_57; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@110820.4]
  wire  dmiProgramBufferRdEn_57; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@110818.4]
  wire  dmiProgramBufferAccessVec_57; // @[Debug.scala 1144:108:freechips.rocketchip.system.DefaultRV32Config.fir@109885.4]
  wire  _T_223; // @[Debug.scala 1147:69:freechips.rocketchip.system.DefaultRV32Config.fir@110015.4]
  wire  dmiProgramBufferWrEnMaybe_58; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@110850.4]
  wire  dmiProgramBufferRdEn_58; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@110848.4]
  wire  dmiProgramBufferAccessVec_58; // @[Debug.scala 1144:108:freechips.rocketchip.system.DefaultRV32Config.fir@109886.4]
  wire  _T_224; // @[Debug.scala 1147:69:freechips.rocketchip.system.DefaultRV32Config.fir@110016.4]
  wire  dmiProgramBufferWrEnMaybe_59; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@110880.4]
  wire  dmiProgramBufferRdEn_59; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@110878.4]
  wire  dmiProgramBufferAccessVec_59; // @[Debug.scala 1144:108:freechips.rocketchip.system.DefaultRV32Config.fir@109887.4]
  wire  _T_225; // @[Debug.scala 1147:69:freechips.rocketchip.system.DefaultRV32Config.fir@110017.4]
  wire  _T_226; // @[Debug.scala 1147:69:freechips.rocketchip.system.DefaultRV32Config.fir@110018.4]
  wire  dmiProgramBufferWrEnMaybe_61; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@113253.4]
  wire  dmiProgramBufferRdEn_61; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@113251.4]
  wire  dmiProgramBufferAccessVec_61; // @[Debug.scala 1144:108:freechips.rocketchip.system.DefaultRV32Config.fir@109889.4]
  wire  _T_227; // @[Debug.scala 1147:69:freechips.rocketchip.system.DefaultRV32Config.fir@110019.4]
  wire  dmiProgramBufferWrEnMaybe_62; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@113283.4]
  wire  dmiProgramBufferRdEn_62; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@113281.4]
  wire  dmiProgramBufferAccessVec_62; // @[Debug.scala 1144:108:freechips.rocketchip.system.DefaultRV32Config.fir@109890.4]
  wire  _T_228; // @[Debug.scala 1147:69:freechips.rocketchip.system.DefaultRV32Config.fir@110020.4]
  wire  dmiProgramBufferWrEnMaybe_63; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@113313.4]
  wire  dmiProgramBufferRdEn_63; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@113311.4]
  wire  dmiProgramBufferAccessVec_63; // @[Debug.scala 1144:108:freechips.rocketchip.system.DefaultRV32Config.fir@109891.4]
  wire  dmiProgramBufferAccess; // @[Debug.scala 1147:69:freechips.rocketchip.system.DefaultRV32Config.fir@110021.4]
  wire  _T_44800; // @[Debug.scala 1580:42:freechips.rocketchip.system.DefaultRV32Config.fir@168687.4]
  wire  errorBusy; // @[Debug.scala 1579:74:freechips.rocketchip.system.DefaultRV32Config.fir@168688.4]
  wire  _T_91; // @[Debug.scala 1132:38:freechips.rocketchip.system.DefaultRV32Config.fir@109669.6]
  wire [15:0] ABSTRACTAUTOWrData_autoexecprogbuf; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@110648.4]
  wire  _T_93; // @[Debug.scala 1135:35:freechips.rocketchip.system.DefaultRV32Config.fir@109674.6]
  wire [11:0] ABSTRACTAUTOWrData_autoexecdata; // @[:freechips.rocketchip.system.DefaultRV32Config.fir@109644.4 :freechips.rocketchip.system.DefaultRV32Config.fir@109645.4 Debug.scala 278:12:freechips.rocketchip.system.DefaultRV32Config.fir@110602.4]
  wire [11:0] _T_94; // @[Debug.scala 1136:73:freechips.rocketchip.system.DefaultRV32Config.fir@109676.8]
  wire [23:0] COMMANDWrData_control; // @[Debug.scala 1163:65:freechips.rocketchip.system.DefaultRV32Config.fir@110150.4]
  reg [7:0] abstractDataMem_0; // @[Debug.scala 1183:36:freechips.rocketchip.system.DefaultRV32Config.fir@110177.4]
  reg [7:0] abstractDataMem_1; // @[Debug.scala 1183:36:freechips.rocketchip.system.DefaultRV32Config.fir@110177.4]
  reg [7:0] abstractDataMem_2; // @[Debug.scala 1183:36:freechips.rocketchip.system.DefaultRV32Config.fir@110177.4]
  reg [7:0] abstractDataMem_3; // @[Debug.scala 1183:36:freechips.rocketchip.system.DefaultRV32Config.fir@110177.4]
  reg [7:0] programBufferMem_0; // @[Debug.scala 1187:34:freechips.rocketchip.system.DefaultRV32Config.fir@110183.4]
  reg [7:0] programBufferMem_1; // @[Debug.scala 1187:34:freechips.rocketchip.system.DefaultRV32Config.fir@110183.4]
  reg [7:0] programBufferMem_2; // @[Debug.scala 1187:34:freechips.rocketchip.system.DefaultRV32Config.fir@110183.4]
  reg [7:0] programBufferMem_3; // @[Debug.scala 1187:34:freechips.rocketchip.system.DefaultRV32Config.fir@110183.4]
  reg [7:0] programBufferMem_4; // @[Debug.scala 1187:34:freechips.rocketchip.system.DefaultRV32Config.fir@110183.4]
  reg [7:0] programBufferMem_5; // @[Debug.scala 1187:34:freechips.rocketchip.system.DefaultRV32Config.fir@110183.4]
  reg [7:0] programBufferMem_6; // @[Debug.scala 1187:34:freechips.rocketchip.system.DefaultRV32Config.fir@110183.4]
  reg [7:0] programBufferMem_7; // @[Debug.scala 1187:34:freechips.rocketchip.system.DefaultRV32Config.fir@110183.4]
  reg [7:0] programBufferMem_8; // @[Debug.scala 1187:34:freechips.rocketchip.system.DefaultRV32Config.fir@110183.4]
  reg [7:0] programBufferMem_9; // @[Debug.scala 1187:34:freechips.rocketchip.system.DefaultRV32Config.fir@110183.4]
  reg [7:0] programBufferMem_10; // @[Debug.scala 1187:34:freechips.rocketchip.system.DefaultRV32Config.fir@110183.4]
  reg [7:0] programBufferMem_11; // @[Debug.scala 1187:34:freechips.rocketchip.system.DefaultRV32Config.fir@110183.4]
  reg [7:0] programBufferMem_12; // @[Debug.scala 1187:34:freechips.rocketchip.system.DefaultRV32Config.fir@110183.4]
  reg [7:0] programBufferMem_13; // @[Debug.scala 1187:34:freechips.rocketchip.system.DefaultRV32Config.fir@110183.4]
  reg [7:0] programBufferMem_14; // @[Debug.scala 1187:34:freechips.rocketchip.system.DefaultRV32Config.fir@110183.4]
  reg [7:0] programBufferMem_15; // @[Debug.scala 1187:34:freechips.rocketchip.system.DefaultRV32Config.fir@110183.4]
  reg [7:0] programBufferMem_16; // @[Debug.scala 1187:34:freechips.rocketchip.system.DefaultRV32Config.fir@110183.4]
  reg [7:0] programBufferMem_17; // @[Debug.scala 1187:34:freechips.rocketchip.system.DefaultRV32Config.fir@110183.4]
  reg [7:0] programBufferMem_18; // @[Debug.scala 1187:34:freechips.rocketchip.system.DefaultRV32Config.fir@110183.4]
  reg [7:0] programBufferMem_19; // @[Debug.scala 1187:34:freechips.rocketchip.system.DefaultRV32Config.fir@110183.4]
  reg [7:0] programBufferMem_20; // @[Debug.scala 1187:34:freechips.rocketchip.system.DefaultRV32Config.fir@110183.4]
  reg [7:0] programBufferMem_21; // @[Debug.scala 1187:34:freechips.rocketchip.system.DefaultRV32Config.fir@110183.4]
  reg [7:0] programBufferMem_22; // @[Debug.scala 1187:34:freechips.rocketchip.system.DefaultRV32Config.fir@110183.4]
  reg [7:0] programBufferMem_23; // @[Debug.scala 1187:34:freechips.rocketchip.system.DefaultRV32Config.fir@110183.4]
  reg [7:0] programBufferMem_24; // @[Debug.scala 1187:34:freechips.rocketchip.system.DefaultRV32Config.fir@110183.4]
  reg [7:0] programBufferMem_25; // @[Debug.scala 1187:34:freechips.rocketchip.system.DefaultRV32Config.fir@110183.4]
  reg [7:0] programBufferMem_26; // @[Debug.scala 1187:34:freechips.rocketchip.system.DefaultRV32Config.fir@110183.4]
  reg [7:0] programBufferMem_27; // @[Debug.scala 1187:34:freechips.rocketchip.system.DefaultRV32Config.fir@110183.4]
  reg [7:0] programBufferMem_28; // @[Debug.scala 1187:34:freechips.rocketchip.system.DefaultRV32Config.fir@110183.4]
  reg [7:0] programBufferMem_29; // @[Debug.scala 1187:34:freechips.rocketchip.system.DefaultRV32Config.fir@110183.4]
  reg [7:0] programBufferMem_30; // @[Debug.scala 1187:34:freechips.rocketchip.system.DefaultRV32Config.fir@110183.4]
  reg [7:0] programBufferMem_31; // @[Debug.scala 1187:34:freechips.rocketchip.system.DefaultRV32Config.fir@110183.4]
  reg [7:0] programBufferMem_32; // @[Debug.scala 1187:34:freechips.rocketchip.system.DefaultRV32Config.fir@110183.4]
  reg [7:0] programBufferMem_33; // @[Debug.scala 1187:34:freechips.rocketchip.system.DefaultRV32Config.fir@110183.4]
  reg [7:0] programBufferMem_34; // @[Debug.scala 1187:34:freechips.rocketchip.system.DefaultRV32Config.fir@110183.4]
  reg [7:0] programBufferMem_35; // @[Debug.scala 1187:34:freechips.rocketchip.system.DefaultRV32Config.fir@110183.4]
  reg [7:0] programBufferMem_36; // @[Debug.scala 1187:34:freechips.rocketchip.system.DefaultRV32Config.fir@110183.4]
  reg [7:0] programBufferMem_37; // @[Debug.scala 1187:34:freechips.rocketchip.system.DefaultRV32Config.fir@110183.4]
  reg [7:0] programBufferMem_38; // @[Debug.scala 1187:34:freechips.rocketchip.system.DefaultRV32Config.fir@110183.4]
  reg [7:0] programBufferMem_39; // @[Debug.scala 1187:34:freechips.rocketchip.system.DefaultRV32Config.fir@110183.4]
  reg [7:0] programBufferMem_40; // @[Debug.scala 1187:34:freechips.rocketchip.system.DefaultRV32Config.fir@110183.4]
  reg [7:0] programBufferMem_41; // @[Debug.scala 1187:34:freechips.rocketchip.system.DefaultRV32Config.fir@110183.4]
  reg [7:0] programBufferMem_42; // @[Debug.scala 1187:34:freechips.rocketchip.system.DefaultRV32Config.fir@110183.4]
  reg [7:0] programBufferMem_43; // @[Debug.scala 1187:34:freechips.rocketchip.system.DefaultRV32Config.fir@110183.4]
  reg [7:0] programBufferMem_44; // @[Debug.scala 1187:34:freechips.rocketchip.system.DefaultRV32Config.fir@110183.4]
  reg [7:0] programBufferMem_45; // @[Debug.scala 1187:34:freechips.rocketchip.system.DefaultRV32Config.fir@110183.4]
  reg [7:0] programBufferMem_46; // @[Debug.scala 1187:34:freechips.rocketchip.system.DefaultRV32Config.fir@110183.4]
  reg [7:0] programBufferMem_47; // @[Debug.scala 1187:34:freechips.rocketchip.system.DefaultRV32Config.fir@110183.4]
  reg [7:0] programBufferMem_48; // @[Debug.scala 1187:34:freechips.rocketchip.system.DefaultRV32Config.fir@110183.4]
  reg [7:0] programBufferMem_49; // @[Debug.scala 1187:34:freechips.rocketchip.system.DefaultRV32Config.fir@110183.4]
  reg [7:0] programBufferMem_50; // @[Debug.scala 1187:34:freechips.rocketchip.system.DefaultRV32Config.fir@110183.4]
  reg [7:0] programBufferMem_51; // @[Debug.scala 1187:34:freechips.rocketchip.system.DefaultRV32Config.fir@110183.4]
  reg [7:0] programBufferMem_52; // @[Debug.scala 1187:34:freechips.rocketchip.system.DefaultRV32Config.fir@110183.4]
  reg [7:0] programBufferMem_53; // @[Debug.scala 1187:34:freechips.rocketchip.system.DefaultRV32Config.fir@110183.4]
  reg [7:0] programBufferMem_54; // @[Debug.scala 1187:34:freechips.rocketchip.system.DefaultRV32Config.fir@110183.4]
  reg [7:0] programBufferMem_55; // @[Debug.scala 1187:34:freechips.rocketchip.system.DefaultRV32Config.fir@110183.4]
  reg [7:0] programBufferMem_56; // @[Debug.scala 1187:34:freechips.rocketchip.system.DefaultRV32Config.fir@110183.4]
  reg [7:0] programBufferMem_57; // @[Debug.scala 1187:34:freechips.rocketchip.system.DefaultRV32Config.fir@110183.4]
  reg [7:0] programBufferMem_58; // @[Debug.scala 1187:34:freechips.rocketchip.system.DefaultRV32Config.fir@110183.4]
  reg [7:0] programBufferMem_59; // @[Debug.scala 1187:34:freechips.rocketchip.system.DefaultRV32Config.fir@110183.4]
  reg [7:0] programBufferMem_60; // @[Debug.scala 1187:34:freechips.rocketchip.system.DefaultRV32Config.fir@110183.4]
  reg [7:0] programBufferMem_61; // @[Debug.scala 1187:34:freechips.rocketchip.system.DefaultRV32Config.fir@110183.4]
  reg [7:0] programBufferMem_62; // @[Debug.scala 1187:34:freechips.rocketchip.system.DefaultRV32Config.fir@110183.4]
  reg [7:0] programBufferMem_63; // @[Debug.scala 1187:34:freechips.rocketchip.system.DefaultRV32Config.fir@110183.4]
  wire  _T_42528; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@162780.4]
  wire  _T_42529; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@162781.4]
  wire  hartResumingWrEn; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@134493.4]
  wire  _GEN_68; // @[Debug.scala 1208:39:freechips.rocketchip.system.DefaultRV32Config.fir@110269.10]
  wire  _T_42518; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@162764.4]
  wire  _T_42519; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@162765.4]
  wire  hartHaltedWrEn; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@130810.4]
  wire  _GEN_69; // @[Debug.scala 1204:37:freechips.rocketchip.system.DefaultRV32Config.fir@110262.8]
  wire  _GEN_71; // @[Debug.scala 1201:45:freechips.rocketchip.system.DefaultRV32Config.fir@110257.6]
  wire  _GEN_73; // @[Debug.scala 1218:33:freechips.rocketchip.system.DefaultRV32Config.fir@110275.6]
  wire  _GEN_74; // @[Debug.scala 1223:52:freechips.rocketchip.system.DefaultRV32Config.fir@110282.6]
  wire [31:0] _T_564; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@110585.4]
  wire [1:0] _T_610; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@110633.4]
  wire [15:0] _T_611; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@110634.4]
  wire [31:0] _T_635; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@110660.4]
  wire [31:0] _T_733; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@110778.4]
  wire [31:0] _T_831; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@110896.4]
  wire [31:0] _T_929; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@111014.4]
  wire [31:0] _T_1027; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@111132.4]
  wire [31:0] _T_1125; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@111250.4]
  wire [31:0] _T_1223; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@111368.4]
  wire [31:0] _T_1321; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@111486.4]
  wire [31:0] _T_1419; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@111604.4]
  wire [16:0] _T_1760; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@111945.4]
  wire [20:0] _T_1852; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@112037.4]
  wire [21:0] _T_1853; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@112038.4]
  wire [22:0] _T_1875; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@112060.4]
  wire  abstractCommandBusy; // @[Debug.scala 1567:42:freechips.rocketchip.system.DefaultRV32Config.fir@168660.4]
  wire [13:0] _T_2013; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@112200.4]
  wire [23:0] _T_2014; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@112201.4]
  wire [28:0] _T_2036; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@112223.4]
  wire [31:0] _T_2134; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@112341.4]
  wire [31:0] _T_2232; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@112459.4]
  wire [31:0] _T_2330; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@112577.4]
  wire [31:0] _T_2541; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@112808.4]
  wire [31:0] _T_2639; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@112926.4]
  wire [31:0] _T_2760; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@113072.4]
  wire [31:0] _T_2879; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@113211.4]
  wire [31:0] _T_2977; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@113329.4]
  wire  _GEN_275; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@114936.4]
  wire  _GEN_276; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@114936.4]
  wire  _GEN_277; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@114936.4]
  wire  _GEN_278; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@114936.4]
  wire  _GEN_3664; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@114936.4]
  wire  _GEN_279; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@114936.4]
  wire  _GEN_280; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@114936.4]
  wire  _GEN_281; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@114936.4]
  wire  _GEN_282; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@114936.4]
  wire  _GEN_3665; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@114936.4]
  wire  _GEN_283; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@114936.4]
  wire  _GEN_3666; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@114936.4]
  wire  _GEN_284; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@114936.4]
  wire  _GEN_3667; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@114936.4]
  wire  _GEN_285; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@114936.4]
  wire  _GEN_3668; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@114936.4]
  wire  _GEN_286; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@114936.4]
  wire  _GEN_3669; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@114936.4]
  wire  _GEN_287; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@114936.4]
  wire  _GEN_3670; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@114936.4]
  wire  _GEN_288; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@114936.4]
  wire  _GEN_3671; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@114936.4]
  wire  _GEN_289; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@114936.4]
  wire  _GEN_290; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@114936.4]
  wire  _GEN_291; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@114936.4]
  wire  _GEN_292; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@114936.4]
  wire  _GEN_293; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@114936.4]
  wire  _GEN_294; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@114936.4]
  wire  _GEN_295; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@114936.4]
  wire  _GEN_296; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@114936.4]
  wire  _GEN_297; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@114936.4]
  wire  _GEN_298; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@114936.4]
  wire  _GEN_299; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@114936.4]
  wire  _GEN_300; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@114936.4]
  wire  _GEN_301; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@114936.4]
  wire  _GEN_302; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@114936.4]
  wire  _GEN_303; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@114936.4]
  wire  _GEN_304; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@114936.4]
  wire  _GEN_305; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@114936.4]
  wire [31:0] _T_3740_1; // @[MuxLiteral.scala 48:48:freechips.rocketchip.system.DefaultRV32Config.fir@114938.4 MuxLiteral.scala 48:48:freechips.rocketchip.system.DefaultRV32Config.fir@114941.4]
  wire [31:0] _GEN_307; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@114972.4]
  wire [31:0] _GEN_308; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@114972.4]
  wire [31:0] _GEN_309; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@114972.4]
  wire [31:0] _GEN_310; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@114972.4]
  wire [31:0] _GEN_311; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@114972.4]
  wire [31:0] _T_3740_6; // @[MuxLiteral.scala 48:48:freechips.rocketchip.system.DefaultRV32Config.fir@114938.4 MuxLiteral.scala 48:48:freechips.rocketchip.system.DefaultRV32Config.fir@114946.4]
  wire [31:0] _GEN_312; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@114972.4]
  wire [31:0] _GEN_313; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@114972.4]
  wire [31:0] _GEN_314; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@114972.4]
  wire [31:0] _GEN_315; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@114972.4]
  wire [31:0] _GEN_316; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@114972.4]
  wire [31:0] _GEN_317; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@114972.4]
  wire [31:0] _GEN_318; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@114972.4]
  wire [31:0] _GEN_319; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@114972.4]
  wire [31:0] _GEN_320; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@114972.4]
  wire [31:0] _GEN_321; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@114972.4]
  wire [31:0] _GEN_322; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@114972.4]
  wire [31:0] _GEN_323; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@114972.4]
  wire [31:0] _GEN_324; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@114972.4]
  wire [31:0] _GEN_325; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@114972.4]
  wire [31:0] _GEN_326; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@114972.4]
  wire [31:0] _GEN_327; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@114972.4]
  wire [31:0] _GEN_328; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@114972.4]
  wire [31:0] _GEN_329; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@114972.4]
  wire [31:0] _GEN_330; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@114972.4]
  wire [31:0] _GEN_331; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@114972.4]
  wire [31:0] _GEN_332; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@114972.4]
  wire [31:0] _GEN_333; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@114972.4]
  wire [31:0] _GEN_334; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@114972.4]
  wire [31:0] _GEN_335; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@114972.4]
  wire [31:0] _GEN_336; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@114972.4]
  wire [31:0] _GEN_337; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@114972.4]
  wire  _T_3749; // @[Debug.scala 1346:60:freechips.rocketchip.system.DefaultRV32Config.fir@115004.4]
  wire  _T_3751; // @[Debug.scala 1346:60:freechips.rocketchip.system.DefaultRV32Config.fir@115009.4]
  wire  _T_3753; // @[Debug.scala 1346:60:freechips.rocketchip.system.DefaultRV32Config.fir@115014.4]
  wire  _T_3755; // @[Debug.scala 1346:60:freechips.rocketchip.system.DefaultRV32Config.fir@115019.4]
  wire  _T_3757; // @[Debug.scala 1368:61:freechips.rocketchip.system.DefaultRV32Config.fir@115024.4]
  wire  _T_3759; // @[Debug.scala 1368:61:freechips.rocketchip.system.DefaultRV32Config.fir@115029.4]
  wire  _T_3761; // @[Debug.scala 1368:61:freechips.rocketchip.system.DefaultRV32Config.fir@115034.4]
  wire  _T_3763; // @[Debug.scala 1368:61:freechips.rocketchip.system.DefaultRV32Config.fir@115039.4]
  wire  _T_3765; // @[Debug.scala 1368:61:freechips.rocketchip.system.DefaultRV32Config.fir@115044.4]
  wire  _T_3767; // @[Debug.scala 1368:61:freechips.rocketchip.system.DefaultRV32Config.fir@115049.4]
  wire  _T_3769; // @[Debug.scala 1368:61:freechips.rocketchip.system.DefaultRV32Config.fir@115054.4]
  wire  _T_3771; // @[Debug.scala 1368:61:freechips.rocketchip.system.DefaultRV32Config.fir@115059.4]
  wire  _T_3773; // @[Debug.scala 1368:61:freechips.rocketchip.system.DefaultRV32Config.fir@115064.4]
  wire  _T_3775; // @[Debug.scala 1368:61:freechips.rocketchip.system.DefaultRV32Config.fir@115069.4]
  wire  _T_3777; // @[Debug.scala 1368:61:freechips.rocketchip.system.DefaultRV32Config.fir@115074.4]
  wire  _T_3779; // @[Debug.scala 1368:61:freechips.rocketchip.system.DefaultRV32Config.fir@115079.4]
  wire  _T_3781; // @[Debug.scala 1368:61:freechips.rocketchip.system.DefaultRV32Config.fir@115084.4]
  wire  _T_3783; // @[Debug.scala 1368:61:freechips.rocketchip.system.DefaultRV32Config.fir@115089.4]
  wire  _T_3785; // @[Debug.scala 1368:61:freechips.rocketchip.system.DefaultRV32Config.fir@115094.4]
  wire  _T_3787; // @[Debug.scala 1368:61:freechips.rocketchip.system.DefaultRV32Config.fir@115099.4]
  wire  _T_3789; // @[Debug.scala 1368:61:freechips.rocketchip.system.DefaultRV32Config.fir@115104.4]
  wire  _T_3791; // @[Debug.scala 1368:61:freechips.rocketchip.system.DefaultRV32Config.fir@115109.4]
  wire  _T_3793; // @[Debug.scala 1368:61:freechips.rocketchip.system.DefaultRV32Config.fir@115114.4]
  wire  _T_3795; // @[Debug.scala 1368:61:freechips.rocketchip.system.DefaultRV32Config.fir@115119.4]
  wire  _T_3797; // @[Debug.scala 1368:61:freechips.rocketchip.system.DefaultRV32Config.fir@115124.4]
  wire  _T_3799; // @[Debug.scala 1368:61:freechips.rocketchip.system.DefaultRV32Config.fir@115129.4]
  wire  _T_3801; // @[Debug.scala 1368:61:freechips.rocketchip.system.DefaultRV32Config.fir@115134.4]
  wire  _T_3803; // @[Debug.scala 1368:61:freechips.rocketchip.system.DefaultRV32Config.fir@115139.4]
  wire  _T_3805; // @[Debug.scala 1368:61:freechips.rocketchip.system.DefaultRV32Config.fir@115144.4]
  wire  _T_3807; // @[Debug.scala 1368:61:freechips.rocketchip.system.DefaultRV32Config.fir@115149.4]
  wire  _T_3809; // @[Debug.scala 1368:61:freechips.rocketchip.system.DefaultRV32Config.fir@115154.4]
  wire  _T_3811; // @[Debug.scala 1368:61:freechips.rocketchip.system.DefaultRV32Config.fir@115159.4]
  wire  _T_3813; // @[Debug.scala 1368:61:freechips.rocketchip.system.DefaultRV32Config.fir@115164.4]
  wire  _T_3815; // @[Debug.scala 1368:61:freechips.rocketchip.system.DefaultRV32Config.fir@115169.4]
  wire  _T_3817; // @[Debug.scala 1368:61:freechips.rocketchip.system.DefaultRV32Config.fir@115174.4]
  wire  _T_3819; // @[Debug.scala 1368:61:freechips.rocketchip.system.DefaultRV32Config.fir@115179.4]
  wire  _T_3821; // @[Debug.scala 1368:61:freechips.rocketchip.system.DefaultRV32Config.fir@115184.4]
  wire  _T_3823; // @[Debug.scala 1368:61:freechips.rocketchip.system.DefaultRV32Config.fir@115189.4]
  wire  _T_3825; // @[Debug.scala 1368:61:freechips.rocketchip.system.DefaultRV32Config.fir@115194.4]
  wire  _T_3827; // @[Debug.scala 1368:61:freechips.rocketchip.system.DefaultRV32Config.fir@115199.4]
  wire  _T_3829; // @[Debug.scala 1368:61:freechips.rocketchip.system.DefaultRV32Config.fir@115204.4]
  wire  _T_3831; // @[Debug.scala 1368:61:freechips.rocketchip.system.DefaultRV32Config.fir@115209.4]
  wire  _T_3833; // @[Debug.scala 1368:61:freechips.rocketchip.system.DefaultRV32Config.fir@115214.4]
  wire  _T_3835; // @[Debug.scala 1368:61:freechips.rocketchip.system.DefaultRV32Config.fir@115219.4]
  wire  _T_3837; // @[Debug.scala 1368:61:freechips.rocketchip.system.DefaultRV32Config.fir@115224.4]
  wire  _T_3839; // @[Debug.scala 1368:61:freechips.rocketchip.system.DefaultRV32Config.fir@115229.4]
  wire  _T_3841; // @[Debug.scala 1368:61:freechips.rocketchip.system.DefaultRV32Config.fir@115234.4]
  wire  _T_3843; // @[Debug.scala 1368:61:freechips.rocketchip.system.DefaultRV32Config.fir@115239.4]
  wire  _T_3845; // @[Debug.scala 1368:61:freechips.rocketchip.system.DefaultRV32Config.fir@115244.4]
  wire  _T_3847; // @[Debug.scala 1368:61:freechips.rocketchip.system.DefaultRV32Config.fir@115249.4]
  wire  _T_3849; // @[Debug.scala 1368:61:freechips.rocketchip.system.DefaultRV32Config.fir@115254.4]
  wire  _T_3851; // @[Debug.scala 1368:61:freechips.rocketchip.system.DefaultRV32Config.fir@115259.4]
  wire  _T_3853; // @[Debug.scala 1368:61:freechips.rocketchip.system.DefaultRV32Config.fir@115264.4]
  wire  _T_3855; // @[Debug.scala 1368:61:freechips.rocketchip.system.DefaultRV32Config.fir@115269.4]
  wire  _T_3857; // @[Debug.scala 1368:61:freechips.rocketchip.system.DefaultRV32Config.fir@115274.4]
  wire  _T_3859; // @[Debug.scala 1368:61:freechips.rocketchip.system.DefaultRV32Config.fir@115279.4]
  wire  _T_3861; // @[Debug.scala 1368:61:freechips.rocketchip.system.DefaultRV32Config.fir@115284.4]
  wire  _T_3863; // @[Debug.scala 1368:61:freechips.rocketchip.system.DefaultRV32Config.fir@115289.4]
  wire  _T_3865; // @[Debug.scala 1368:61:freechips.rocketchip.system.DefaultRV32Config.fir@115294.4]
  wire  _T_3867; // @[Debug.scala 1368:61:freechips.rocketchip.system.DefaultRV32Config.fir@115299.4]
  wire  _T_3869; // @[Debug.scala 1368:61:freechips.rocketchip.system.DefaultRV32Config.fir@115304.4]
  wire  _T_3871; // @[Debug.scala 1368:61:freechips.rocketchip.system.DefaultRV32Config.fir@115309.4]
  wire  _T_3873; // @[Debug.scala 1368:61:freechips.rocketchip.system.DefaultRV32Config.fir@115314.4]
  wire  _T_3875; // @[Debug.scala 1368:61:freechips.rocketchip.system.DefaultRV32Config.fir@115319.4]
  wire  _T_3877; // @[Debug.scala 1368:61:freechips.rocketchip.system.DefaultRV32Config.fir@115324.4]
  wire  _T_3879; // @[Debug.scala 1368:61:freechips.rocketchip.system.DefaultRV32Config.fir@115329.4]
  wire  _T_3881; // @[Debug.scala 1368:61:freechips.rocketchip.system.DefaultRV32Config.fir@115334.4]
  wire  _T_3883; // @[Debug.scala 1368:61:freechips.rocketchip.system.DefaultRV32Config.fir@115339.4]
  reg  goReg; // @[Debug.scala 1377:27:freechips.rocketchip.system.DefaultRV32Config.fir@115343.4]
  wire [9:0] hartGoingId; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@126788.4]
  wire  _T_3935; // @[Debug.scala 1389:28:freechips.rocketchip.system.DefaultRV32Config.fir@115468.10]
  wire  _T_3937; // @[Debug.scala 1389:15:freechips.rocketchip.system.DefaultRV32Config.fir@115470.10]
  wire  _T_3938; // @[Debug.scala 1389:15:freechips.rocketchip.system.DefaultRV32Config.fir@115471.10]
  wire  _T_42523; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@162772.4]
  wire  _T_42524; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@162773.4]
  wire  hartGoingWrEn; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@126787.4]
  wire  _GEN_406; // @[Debug.scala 1388:33:freechips.rocketchip.system.DefaultRV32Config.fir@115467.8]
  wire  _GEN_3637; // @[Debug.scala 1633:43:freechips.rocketchip.system.DefaultRV32Config.fir@168747.10]
  wire  _GEN_3641; // @[Debug.scala 1630:38:freechips.rocketchip.system.DefaultRV32Config.fir@168742.8]
  wire  _GEN_3654; // @[Debug.scala 1623:59:freechips.rocketchip.system.DefaultRV32Config.fir@168741.6]
  wire  goAbstract; // @[Debug.scala 1615:47:freechips.rocketchip.system.DefaultRV32Config.fir@168724.4]
  wire  _GEN_407; // @[Debug.scala 1386:25:freechips.rocketchip.system.DefaultRV32Config.fir@115463.6]
  wire  accessRegisterCommandReg_postexec; // @[Debug.scala 1415:73:freechips.rocketchip.system.DefaultRV32Config.fir@115554.4]
  wire [2:0] accessRegisterCommandReg_size; // @[Debug.scala 1415:73:freechips.rocketchip.system.DefaultRV32Config.fir@115558.4]
  reg [31:0] abstractGeneratedMem_0; // @[Debug.scala 1458:35:freechips.rocketchip.system.DefaultRV32Config.fir@115573.4]
  reg [31:0] abstractGeneratedMem_1; // @[Debug.scala 1458:35:freechips.rocketchip.system.DefaultRV32Config.fir@115573.4]
  wire [15:0] _T_3972; // @[Debug.scala 1464:66:freechips.rocketchip.system.DefaultRV32Config.fir@115584.4]
  wire [4:0] abstractGeneratedI_rd; // @[Debug.scala 1459:34:freechips.rocketchip.system.DefaultRV32Config.fir@115574.4 Debug.scala 1464:31:freechips.rocketchip.system.DefaultRV32Config.fir@115585.4]
  wire [31:0] _T_3979; // @[Debug.scala 1485:36:freechips.rocketchip.system.DefaultRV32Config.fir@115621.6]
  wire [31:0] _T_3984; // @[Debug.scala 1487:36:freechips.rocketchip.system.DefaultRV32Config.fir@115626.6]
  wire  _T_6696; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@118357.4]
  wire  _T_6717; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@118378.4]
  wire  _T_6740; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@118401.4]
  wire [23:0] _T_6757; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@118418.4]
  wire  _T_6763; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@118424.4]
  wire [31:0] _T_6780; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@118441.4]
  wire  _T_38152; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@153307.4]
  wire  _T_38153; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@153308.4]
  wire  _T_7603; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@119264.4]
  wire  _T_7626; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@119290.4]
  wire  _T_7651; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@119318.4]
  wire  _T_7676; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@119346.4]
  wire  _T_38147; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@153296.4]
  wire  _T_38148; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@153297.4]
  wire  _T_10671; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@122344.4]
  wire  _T_10694; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@122370.4]
  wire  _T_10719; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@122398.4]
  wire  _T_10744; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@122426.4]
  wire  _T_38122; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@153241.4]
  wire  _T_38123; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@153242.4]
  wire  _T_11219; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@122904.4]
  wire  _T_11242; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@122930.4]
  wire  _T_11267; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@122958.4]
  wire  _T_11292; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@122986.4]
  wire  _T_38172; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@153351.4]
  wire  _T_38173; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@153352.4]
  wire  _T_11947; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@123644.4]
  wire  _T_11970; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@123670.4]
  wire  _T_11995; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@123698.4]
  wire  _T_12020; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@123726.4]
  wire  _T_38167; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@153340.4]
  wire  _T_38168; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@153341.4]
  wire  _T_13686; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@125395.4]
  wire  _T_13709; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@125421.4]
  wire  _T_13734; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@125449.4]
  wire  _T_13759; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@125477.4]
  wire  _T_38187; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@153384.4]
  wire  _T_38188; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@153385.4]
  wire  _T_15806; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@127529.4]
  wire  _T_15829; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@127555.4]
  wire  _T_15854; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@127583.4]
  wire  _T_15879; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@127611.4]
  wire  _T_38127; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@153252.4]
  wire  _T_38128; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@153253.4]
  wire  _T_17254; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@128989.4]
  wire  _T_17277; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@129015.4]
  wire  _T_17302; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@129043.4]
  wire  _T_17327; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@129071.4]
  wire  _T_38162; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@153329.4]
  wire  _T_38163; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@153330.4]
  wire  _T_20793; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@132542.4]
  wire  _T_20816; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@132568.4]
  wire  _T_20841; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@132596.4]
  wire  _T_20866; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@132624.4]
  wire  _T_38107; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@153208.4]
  wire  _T_38108; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@153209.4]
  wire  _T_21791; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@133552.4]
  wire  _T_21814; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@133578.4]
  wire  _T_21839; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@133606.4]
  wire  _T_21864; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@133634.4]
  wire  _T_38132; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@153263.4]
  wire  _T_38133; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@153264.4]
  wire  _T_22429; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@134202.4]
  wire  _T_22452; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@134228.4]
  wire  _T_22477; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@134256.4]
  wire  _T_22502; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@134284.4]
  wire  _T_38182; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@153373.4]
  wire  _T_38183; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@153374.4]
  wire  _T_23268; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@135055.4]
  wire  _T_23291; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@135081.4]
  wire  _T_23316; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@135109.4]
  wire  _T_23341; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@135137.4]
  wire  _T_38112; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@153219.4]
  wire  _T_38113; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@153220.4]
  wire  _T_24446; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@136245.4]
  wire  _T_24469; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@136271.4]
  wire  _T_24494; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@136299.4]
  wire  _T_24519; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@136327.4]
  wire  _T_38157; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@153318.4]
  wire  _T_38158; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@153319.4]
  wire  _T_27445; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@139258.4]
  wire  _T_27468; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@139284.4]
  wire  _T_27493; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@139312.4]
  wire  _T_27518; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@139340.4]
  wire  _T_38137; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@153274.4]
  wire  _T_38138; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@153275.4]
  wire  _T_29094; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@140919.4]
  wire  _T_29117; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@140945.4]
  wire  _T_29142; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@140973.4]
  wire  _T_29167; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@141001.4]
  wire  _T_38117; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@153230.4]
  wire  _T_38118; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@153231.4]
  wire  _T_30272; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@142109.4]
  wire  _T_30295; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@142135.4]
  wire  _T_30320; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@142163.4]
  wire  _T_30345; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@142191.4]
  wire  _T_38142; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@153285.4]
  wire  _T_38143; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@153286.4]
  wire  _T_32890; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@144739.4]
  wire  _T_32913; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@144765.4]
  wire  _T_32938; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@144793.4]
  wire  _T_32963; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@144821.4]
  wire  _T_38177; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@153362.4]
  wire  _T_38178; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@153363.4]
  wire  _T_33078; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@144939.4]
  wire  _T_33101; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@144965.4]
  wire  _T_33126; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@144993.4]
  wire  _T_33151; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@145021.4]
  wire  _GEN_2532; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_2533; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_2534; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_2535; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_2536; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_2537; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_2538; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_2539; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_2540; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_2541; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_2542; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_2543; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_2544; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_2545; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_2546; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_2547; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_2548; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_2549; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_2550; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_2551; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_3672; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_2552; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_3673; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_2553; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_3674; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_2554; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_3675; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_2555; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_3676; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_2556; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_3677; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_2557; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_3678; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_2558; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_3679; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_2559; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_3680; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_2560; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_3681; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_2561; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_3682; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_2562; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_3683; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_2563; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_3684; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_2564; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_3685; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_2565; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_3686; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_2566; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_3687; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_2567; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_3688; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_2568; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_3689; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_2569; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_3690; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_2570; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_3691; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_2571; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_3692; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_2572; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_3693; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_2573; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_3694; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_2574; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_3695; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_2575; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_3696; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_2576; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_3697; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_2577; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_3698; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_2578; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_3699; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_2579; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_3700; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_2580; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_3701; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_2581; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_3702; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_2582; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_3703; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_2583; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_3704; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_2584; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_3705; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_2585; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_3706; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_2586; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_3707; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_2587; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_3708; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_2588; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_3709; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_2589; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_3710; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_2590; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_3711; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_2591; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_3712; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_2592; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_3713; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_2593; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_3714; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_2594; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_2595; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_2596; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_2597; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_2598; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_3715; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_2599; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_3716; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_2600; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_3717; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_2601; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_3718; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_2602; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_3719; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_2603; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_3720; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_2604; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_3721; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_2605; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_3722; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_2606; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_3723; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_2607; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_3724; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_2608; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_3725; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_2609; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_3726; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_2610; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_3727; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_2611; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_3728; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_2612; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_3729; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_2613; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_3730; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_2614; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_3731; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_2615; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_3732; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_2616; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_3733; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_2617; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_3734; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_2618; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_3735; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_2619; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_3736; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_2620; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_3737; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_2621; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_3738; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_2622; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_3739; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_2623; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_3740; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_2624; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_3741; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_2625; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_3742; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_2626; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_3743; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_2627; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_3744; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_2628; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_3745; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_2629; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_3746; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_2630; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_3747; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_2631; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_3748; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_2632; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_3749; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_2633; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_3750; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_2634; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_3751; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_2635; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_3752; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_2636; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_3753; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_2637; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_3754; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_2638; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_3755; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_2639; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_3756; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_2640; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_3757; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_2641; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_3758; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_2642; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_3759; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_2643; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_3760; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_2644; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_3761; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_2645; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_3762; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_2646; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_3763; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_2647; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_3764; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_2648; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_3765; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_2649; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_3766; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_2650; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_3767; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_2651; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_3768; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_2652; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_3769; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_2653; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_3770; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_2654; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_3771; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_2655; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_3772; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_2656; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_3773; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_2657; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_3774; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_2658; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_3775; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_2659; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_3776; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_2660; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_3777; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_2661; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_3778; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_2662; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_3779; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_2663; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_3780; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_2664; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_3781; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_2665; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_3782; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_2666; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_3783; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_2667; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_3784; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_2668; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_3785; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_2669; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_3786; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_2670; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_3787; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_2671; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_3788; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_2672; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_3789; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_2673; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_3790; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_2674; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_3791; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_2675; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_3792; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_2676; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_3793; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_2677; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_3794; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_2678; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_3795; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_2679; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_3796; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_2680; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_3797; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_2681; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_3798; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_2682; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_3799; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_2683; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_3800; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_2684; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_3801; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_2685; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_3802; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_2686; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_3803; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_2687; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_3804; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_2688; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_3805; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_2689; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_3806; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_2690; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_3807; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_2691; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_3808; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_2692; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_3809; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_2693; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_3810; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_2694; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_3811; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_2695; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_3812; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_2696; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_3813; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_2697; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_3814; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_2698; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_3815; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_2699; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_3816; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_2700; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_3817; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_2701; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_3818; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_2702; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_3819; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_2703; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_3820; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_2704; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_3821; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_2705; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_3822; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_2706; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_3823; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_2707; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_3824; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_2708; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_3825; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_2709; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_3826; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_2710; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_3827; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_2711; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_3828; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_2712; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_3829; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_2713; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_3830; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_2714; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_3831; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_2715; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_3832; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_2716; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_3833; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_2717; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_3834; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_2718; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_3835; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_2719; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_3836; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_2720; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_3837; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_2721; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_3838; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_2722; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_2723; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_3839; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_2724; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_3840; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_2725; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_3841; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_2726; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_3842; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_2727; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_3843; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_2728; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_3844; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_2729; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_3845; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_2730; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_3846; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_2731; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_3847; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_2732; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_3848; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_2733; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_3849; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_2734; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_3850; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_2735; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_3851; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_2736; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_2737; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_2738; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_2739; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_2740; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_2741; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_2742; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_2743; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_2744; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_2745; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_2746; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_2747; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_2748; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_2749; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_2750; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_2751; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_2752; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_2753; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_2754; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_2755; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_3852; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_2756; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_3853; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_2757; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_3854; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_2758; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_3855; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_2759; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_3856; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_2760; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_3857; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_2761; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_3858; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_2762; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_3859; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_2763; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_3860; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_2764; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_3861; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_2765; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_3862; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_2766; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_3863; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_2767; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_3864; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_2768; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_3865; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_2769; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_3866; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_2770; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_3867; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_2771; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_3868; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_2772; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_3869; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_2773; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_3870; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_2774; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_3871; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_2775; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_3872; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_2776; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_3873; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_2777; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_3874; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_2778; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_3875; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_2779; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_3876; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_2780; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_3877; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_2781; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_3878; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_2782; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_3879; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_2783; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_3880; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_2784; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_3881; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_2785; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_3882; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_2786; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_2787; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_2788; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_2789; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_2790; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_2791; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_2792; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_2793; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_2794; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_2795; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_2796; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_2797; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_2798; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_2799; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_2800; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_2801; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_2802; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_2803; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_2804; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_2805; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_2806; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_2807; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_2808; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_2809; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_2810; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_2811; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_2812; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_2813; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_2814; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_2815; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_2816; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_2817; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_2818; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_2819; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_2820; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_2821; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_2822; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_2823; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_2824; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_2825; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_2826; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_2827; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_2828; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_2829; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_2830; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_2831; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_2832; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_2833; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_2834; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_2835; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_2836; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_2837; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_2838; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_2839; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_2840; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_2841; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_2842; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_2843; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_2844; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_2845; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_2846; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_2847; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_2848; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_2849; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_2850; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_2851; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_2852; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_2853; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_2854; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_2855; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_2856; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_2857; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_2858; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_2859; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_2860; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_2861; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_2862; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_2863; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_2864; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_2865; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_2866; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_2867; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_2868; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_2869; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_2870; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_2871; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_2872; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_2873; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_2874; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_2875; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_2876; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_2877; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_2878; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_2879; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_2880; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_2881; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_2882; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_2883; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_2884; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_2885; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_2886; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_2887; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_2888; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_2889; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_2890; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_2891; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_2892; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_2893; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_2894; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_2895; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_2896; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_2897; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_2898; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_2899; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_2900; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_2901; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_2902; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_2903; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_2904; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_2905; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_2906; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_2907; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_2908; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_2909; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_2910; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_2911; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_2912; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_2913; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_2914; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_2915; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_2916; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_2917; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_2918; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_2919; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_2920; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_2921; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_2922; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_2923; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_2924; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_2925; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_2926; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_2927; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_2928; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_2929; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_2930; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_2931; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_2932; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_2933; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_2934; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_2935; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_2936; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_2937; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_2938; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_2939; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_2940; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_2941; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_2942; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_2943; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_2944; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_2945; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_2946; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_2947; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_2948; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_2949; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_2950; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_2951; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_2952; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_2953; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_2954; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_2955; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_2956; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_2957; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_2958; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_2959; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_2960; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_2961; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_2962; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_2963; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_2964; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_2965; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_2966; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_2967; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_2968; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_2969; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_2970; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_2971; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_2972; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_2973; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_2974; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_2975; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_2976; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_2977; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_2978; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_2979; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_2980; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_2981; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_2982; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_2983; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_2984; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_2985; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_2986; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_2987; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_2988; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_2989; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_2990; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_2991; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_2992; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_2993; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_2994; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_2995; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_2996; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_2997; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_2998; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_2999; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_3000; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_3001; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_3002; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_3003; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_3004; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_3005; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_3006; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_3007; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_3008; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_3009; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_3010; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_3011; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_3012; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_3013; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_3014; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_3015; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_3016; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_3017; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_3018; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_3019; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_3020; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_3021; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_3022; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_3023; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_3024; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_3025; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_3026; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_3027; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_3028; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_3029; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_3030; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_3031; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_3032; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_3033; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_3034; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_3035; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_3036; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_3037; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_3038; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_3039; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_3040; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_3041; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire  _GEN_3042; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  wire [31:0] _GEN_3044; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  wire [31:0] _GEN_3045; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  wire [31:0] _GEN_3046; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  wire [31:0] _GEN_3047; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  wire [31:0] _GEN_3048; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  wire [31:0] _GEN_3049; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  wire [31:0] _GEN_3050; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  wire [31:0] _GEN_3051; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  wire [31:0] _GEN_3052; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  wire [31:0] _GEN_3053; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  wire [31:0] _GEN_3054; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  wire [31:0] _GEN_3055; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  wire [31:0] _GEN_3056; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  wire [31:0] _GEN_3057; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  wire [31:0] _GEN_3058; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  wire [31:0] _GEN_3059; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  wire [31:0] _GEN_3060; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  wire [31:0] _GEN_3061; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  wire [31:0] _GEN_3062; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  wire [31:0] _GEN_3063; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  wire [31:0] _GEN_3064; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  wire [31:0] _GEN_3065; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  wire [31:0] _GEN_3066; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  wire [31:0] _GEN_3067; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  wire [31:0] _GEN_3068; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  wire [31:0] _GEN_3069; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  wire [31:0] _GEN_3070; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  wire [31:0] _GEN_3071; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  wire [31:0] _GEN_3072; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  wire [31:0] _GEN_3073; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  wire [31:0] _GEN_3074; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  wire [31:0] _GEN_3075; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  wire [31:0] _GEN_3076; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  wire [31:0] _GEN_3077; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  wire [31:0] _GEN_3078; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  wire [31:0] _GEN_3079; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  wire [31:0] _GEN_3080; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  wire [31:0] _GEN_3081; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  wire [31:0] _GEN_3082; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  wire [31:0] _GEN_3083; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  wire [31:0] _GEN_3084; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  wire [31:0] _GEN_3085; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  wire [31:0] _GEN_3086; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  wire [31:0] _GEN_3087; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  wire [31:0] _GEN_3088; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  wire [31:0] _GEN_3089; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  wire [31:0] _GEN_3090; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  wire [31:0] _GEN_3091; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  wire [31:0] _GEN_3092; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  wire [31:0] _GEN_3093; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  wire [31:0] _GEN_3094; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  wire [31:0] _GEN_3095; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  wire [31:0] _GEN_3096; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  wire [31:0] _GEN_3097; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  wire [31:0] _GEN_3098; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  wire [31:0] _GEN_3099; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  wire [31:0] _GEN_3100; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  wire [31:0] _GEN_3101; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  wire [31:0] _GEN_3102; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  wire [31:0] _GEN_3103; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  wire [31:0] _GEN_3104; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  wire [31:0] _GEN_3105; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  wire [31:0] _GEN_3106; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  wire [31:0] _GEN_3107; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  wire [31:0] _GEN_3108; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  wire [31:0] _GEN_3109; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  wire [31:0] _GEN_3110; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  wire [31:0] _GEN_3111; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  wire [31:0] _GEN_3112; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  wire [31:0] _GEN_3113; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  wire [31:0] _GEN_3114; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  wire [31:0] _GEN_3115; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  wire [31:0] _GEN_3116; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  wire [31:0] _GEN_3117; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  wire [31:0] _GEN_3118; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  wire [31:0] _GEN_3119; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  wire [31:0] _GEN_3120; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  wire [31:0] _GEN_3121; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  wire [31:0] _GEN_3122; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  wire [31:0] _GEN_3123; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  wire [31:0] _GEN_3124; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  wire [31:0] _GEN_3125; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  wire [31:0] _GEN_3126; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  wire [31:0] _GEN_3127; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  wire [31:0] _GEN_3128; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  wire [31:0] _GEN_3129; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  wire [31:0] _GEN_3130; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  wire [31:0] _GEN_3131; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  wire [31:0] _GEN_3132; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  wire [31:0] _GEN_3133; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  wire [31:0] _GEN_3134; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  wire [31:0] _GEN_3135; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  wire [31:0] _GEN_3136; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  wire [31:0] _GEN_3137; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  wire [31:0] _GEN_3138; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  wire [31:0] _GEN_3139; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  wire [31:0] _GEN_3140; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  wire [31:0] _GEN_3141; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  wire [31:0] _GEN_3142; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  wire [31:0] _GEN_3143; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  wire [31:0] _GEN_3144; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  wire [31:0] _GEN_3145; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  wire [31:0] _GEN_3146; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  wire [31:0] _GEN_3147; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  wire [31:0] _GEN_3148; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  wire [31:0] _GEN_3149; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  wire [31:0] _GEN_3150; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  wire [31:0] _GEN_3151; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  wire [31:0] _GEN_3152; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  wire [31:0] _GEN_3153; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  wire [31:0] _GEN_3154; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  wire [31:0] _GEN_3155; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  wire [31:0] _GEN_3156; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  wire [31:0] _GEN_3157; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  wire [31:0] _GEN_3158; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  wire [31:0] _GEN_3159; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  wire [31:0] _GEN_3160; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  wire [31:0] _GEN_3161; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  wire [31:0] _GEN_3162; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  wire [31:0] _GEN_3163; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  wire [31:0] _GEN_3164; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  wire [31:0] _GEN_3165; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  wire [31:0] _GEN_3166; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  wire [31:0] _GEN_3167; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  wire [31:0] _GEN_3168; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  wire [31:0] _GEN_3169; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  wire [31:0] _GEN_3170; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  wire [31:0] _GEN_3171; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  wire [31:0] _GEN_3172; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  wire [31:0] _GEN_3173; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  wire [31:0] _GEN_3174; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  wire [31:0] _GEN_3175; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  wire [31:0] _GEN_3176; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  wire [31:0] _GEN_3177; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  wire [31:0] _GEN_3178; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  wire [31:0] _GEN_3179; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  wire [31:0] _GEN_3180; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  wire [31:0] _GEN_3181; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  wire [31:0] _GEN_3182; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  wire [31:0] _GEN_3183; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  wire [31:0] _GEN_3184; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  wire [31:0] _GEN_3185; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  wire [31:0] _GEN_3186; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  wire [31:0] _GEN_3187; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  wire [31:0] _GEN_3188; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  wire [31:0] _GEN_3189; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  wire [31:0] _GEN_3190; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  wire [31:0] _GEN_3191; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  wire [31:0] _GEN_3192; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  wire [31:0] _GEN_3193; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  wire [31:0] _GEN_3194; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  wire [31:0] _GEN_3195; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  wire [31:0] _GEN_3196; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  wire [31:0] _GEN_3197; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  wire [31:0] _GEN_3198; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  wire [31:0] _GEN_3199; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  wire [31:0] _GEN_3200; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  wire [31:0] _GEN_3201; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  wire [31:0] _GEN_3202; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  wire [31:0] _GEN_3203; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  wire [31:0] _GEN_3204; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  wire [31:0] _GEN_3205; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  wire [31:0] _GEN_3206; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  wire [31:0] _GEN_3207; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  wire [31:0] _GEN_3208; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  wire [31:0] _GEN_3209; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  wire [31:0] _GEN_3210; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  wire [31:0] _GEN_3211; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  wire [31:0] _GEN_3212; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  wire [31:0] _GEN_3213; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  wire [31:0] _GEN_3214; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  wire [31:0] _GEN_3215; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  wire [31:0] _GEN_3216; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  wire [31:0] _GEN_3217; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  wire [31:0] _GEN_3218; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  wire [31:0] _GEN_3219; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  wire [31:0] _GEN_3220; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  wire [31:0] _GEN_3221; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  wire [31:0] _GEN_3222; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  wire [31:0] _GEN_3223; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  wire [31:0] _GEN_3224; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  wire [31:0] _GEN_3225; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  wire [31:0] _GEN_3226; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  wire [31:0] _GEN_3227; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  wire [31:0] _GEN_3228; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  wire [31:0] _GEN_3229; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  wire [31:0] _GEN_3230; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  wire [31:0] _GEN_3231; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  wire [31:0] _GEN_3232; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  wire [31:0] _GEN_3233; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  wire [31:0] _GEN_3234; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  wire [31:0] _GEN_3235; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  wire [31:0] _GEN_3236; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  wire [31:0] _GEN_3237; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  wire [31:0] _GEN_3238; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  wire [31:0] _GEN_3239; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  wire [31:0] _GEN_3240; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  wire [31:0] _GEN_3241; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  wire [31:0] _GEN_3242; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  wire [31:0] _GEN_3243; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  wire [31:0] _GEN_3244; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  wire [31:0] _GEN_3245; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  wire [31:0] _GEN_3246; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  wire [31:0] _GEN_3247; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  wire [31:0] _GEN_3248; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  wire [31:0] _GEN_3249; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  wire [31:0] _GEN_3250; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  wire [31:0] _GEN_3251; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  wire [31:0] _GEN_3252; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  wire [31:0] _GEN_3253; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  wire [31:0] _GEN_3254; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  wire [31:0] _GEN_3255; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  wire [31:0] _GEN_3256; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  wire [31:0] _GEN_3257; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  wire [31:0] _GEN_3258; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  wire [31:0] _GEN_3259; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  wire [31:0] _GEN_3260; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  wire [31:0] _GEN_3261; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  wire [31:0] _GEN_3262; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  wire [31:0] _GEN_3263; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  wire [31:0] _GEN_3264; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  wire [31:0] _GEN_3265; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  wire [31:0] _GEN_3266; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  wire [31:0] _GEN_3267; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  wire [31:0] _GEN_3268; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  wire [31:0] _GEN_3269; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  wire [31:0] _GEN_3270; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  wire [31:0] _GEN_3271; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  wire [31:0] _GEN_3272; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  wire [31:0] _GEN_3273; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  wire [31:0] _GEN_3274; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  wire [31:0] _GEN_3275; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  wire [31:0] _GEN_3276; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  wire [31:0] _GEN_3277; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  wire [31:0] _GEN_3278; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  wire [31:0] _GEN_3279; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  wire [31:0] _GEN_3280; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  wire [31:0] _GEN_3281; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  wire [31:0] _GEN_3282; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  wire [31:0] _GEN_3283; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  wire [31:0] _GEN_3284; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  wire [31:0] _GEN_3285; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  wire [31:0] _GEN_3286; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  wire [31:0] _GEN_3287; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  wire [31:0] _GEN_3288; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  wire [31:0] _GEN_3289; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  wire [31:0] _GEN_3290; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  wire [31:0] _GEN_3291; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  wire [31:0] _GEN_3292; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  wire [31:0] _GEN_3293; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  wire [31:0] _GEN_3294; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  wire [31:0] _GEN_3295; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  wire [31:0] _GEN_3296; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  wire [31:0] _GEN_3297; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  wire [31:0] _GEN_3298; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  wire [31:0] _GEN_3299; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  wire [31:0] _GEN_3300; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  wire [31:0] _GEN_3301; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  wire [31:0] _GEN_3302; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  wire [31:0] _GEN_3303; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  wire [31:0] _GEN_3304; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  wire [31:0] _GEN_3305; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  wire [31:0] _GEN_3306; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  wire [31:0] _GEN_3307; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  wire [31:0] _GEN_3308; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  wire [31:0] _GEN_3309; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  wire [31:0] _GEN_3310; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  wire [31:0] _GEN_3311; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  wire [31:0] _GEN_3312; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  wire [31:0] _GEN_3313; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  wire [31:0] _GEN_3314; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  wire [31:0] _GEN_3315; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  wire [31:0] _GEN_3316; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  wire [31:0] _GEN_3317; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  wire [31:0] _GEN_3318; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  wire [31:0] _GEN_3319; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  wire [31:0] _GEN_3320; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  wire [31:0] _GEN_3321; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  wire [31:0] _GEN_3322; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  wire [31:0] _GEN_3323; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  wire [31:0] _GEN_3324; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  wire [31:0] _GEN_3325; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  wire [31:0] _GEN_3326; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  wire [31:0] _GEN_3327; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  wire [31:0] _GEN_3328; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  wire [31:0] _GEN_3329; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  wire [31:0] _GEN_3330; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  wire [31:0] _GEN_3331; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  wire [31:0] _GEN_3332; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  wire [31:0] _GEN_3333; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  wire [31:0] _GEN_3334; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  wire [31:0] _GEN_3335; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  wire [31:0] _GEN_3336; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  wire [31:0] _GEN_3337; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  wire [31:0] _GEN_3338; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  wire [31:0] _GEN_3339; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  wire [31:0] _GEN_3340; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  wire [31:0] _GEN_3341; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  wire [31:0] _GEN_3342; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  wire [31:0] _GEN_3343; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  wire [31:0] _GEN_3344; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  wire [31:0] _GEN_3345; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  wire [31:0] _GEN_3346; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  wire [31:0] _GEN_3347; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  wire [31:0] _GEN_3348; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  wire [31:0] _GEN_3349; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  wire [31:0] _GEN_3350; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  wire [31:0] _GEN_3351; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  wire [31:0] _GEN_3352; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  wire [31:0] _GEN_3353; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  wire [31:0] _GEN_3354; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  wire [31:0] _GEN_3355; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  wire [31:0] _GEN_3356; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  wire [31:0] _GEN_3357; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  wire [31:0] _GEN_3358; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  wire [31:0] _GEN_3359; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  wire [31:0] _GEN_3360; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  wire [31:0] _GEN_3361; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  wire [31:0] _GEN_3362; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  wire [31:0] _GEN_3363; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  wire [31:0] _GEN_3364; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  wire [31:0] _GEN_3365; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  wire [31:0] _GEN_3366; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  wire [31:0] _GEN_3367; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  wire [31:0] _GEN_3368; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  wire [31:0] _GEN_3369; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  wire [31:0] _GEN_3370; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  wire [31:0] _GEN_3371; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  wire [31:0] _GEN_3372; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  wire [31:0] _GEN_3373; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  wire [31:0] _GEN_3374; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  wire [31:0] _GEN_3375; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  wire [31:0] _GEN_3376; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  wire [31:0] _GEN_3377; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  wire [31:0] _GEN_3378; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  wire [31:0] _GEN_3379; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  wire [31:0] _GEN_3380; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  wire [31:0] _GEN_3381; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  wire [31:0] _GEN_3382; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  wire [31:0] _GEN_3383; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  wire [31:0] _GEN_3384; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  wire [31:0] _GEN_3385; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  wire [31:0] _GEN_3386; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  wire [31:0] _GEN_3387; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  wire [31:0] _GEN_3388; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  wire [31:0] _GEN_3389; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  wire [31:0] _GEN_3390; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  wire [31:0] _GEN_3391; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  wire [31:0] _GEN_3392; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  wire [31:0] _GEN_3393; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  wire [31:0] _GEN_3394; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  wire [31:0] _GEN_3395; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  wire [31:0] _GEN_3396; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  wire [31:0] _GEN_3397; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  wire [31:0] _GEN_3398; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  wire [31:0] _GEN_3399; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  wire [31:0] _GEN_3400; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  wire [31:0] _GEN_3401; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  wire [31:0] _GEN_3402; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  wire [31:0] _GEN_3403; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  wire [31:0] _GEN_3404; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  wire [31:0] _GEN_3405; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  wire [31:0] _GEN_3406; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  wire [31:0] _GEN_3407; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  wire [31:0] _GEN_3408; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  wire [31:0] _GEN_3409; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  wire [31:0] _GEN_3410; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  wire [31:0] _GEN_3411; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  wire [31:0] _GEN_3412; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  wire [31:0] _GEN_3413; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  wire [31:0] _GEN_3414; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  wire [31:0] _GEN_3415; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  wire [31:0] _GEN_3416; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  wire [31:0] _GEN_3417; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  wire [31:0] _GEN_3418; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  wire [31:0] _GEN_3419; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  wire [31:0] _GEN_3420; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  wire [31:0] _GEN_3421; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  wire [31:0] _GEN_3422; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  wire [31:0] _GEN_3423; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  wire [31:0] _GEN_3424; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  wire [31:0] _GEN_3425; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  wire [31:0] _GEN_3426; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  wire [31:0] _GEN_3427; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  wire [31:0] _GEN_3428; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  wire [31:0] _GEN_3429; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  wire [31:0] _GEN_3430; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  wire [31:0] _GEN_3431; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  wire [31:0] _GEN_3432; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  wire [31:0] _GEN_3433; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  wire [31:0] _GEN_3434; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  wire [31:0] _GEN_3435; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  wire [31:0] _GEN_3436; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  wire [31:0] _GEN_3437; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  wire [31:0] _GEN_3438; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  wire [31:0] _GEN_3439; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  wire [31:0] _GEN_3440; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  wire [31:0] _GEN_3441; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  wire [31:0] _GEN_3442; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  wire [31:0] _GEN_3443; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  wire [31:0] _GEN_3444; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  wire [31:0] _GEN_3445; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  wire [31:0] _GEN_3446; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  wire [31:0] _GEN_3447; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  wire [31:0] _GEN_3448; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  wire [31:0] _GEN_3449; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  wire [31:0] _GEN_3450; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  wire [31:0] _GEN_3451; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  wire [31:0] _GEN_3452; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  wire [31:0] _GEN_3453; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  wire [31:0] _GEN_3454; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  wire [31:0] _GEN_3455; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  wire [31:0] _GEN_3456; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  wire [31:0] _GEN_3457; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  wire [31:0] _GEN_3458; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  wire [31:0] _GEN_3459; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  wire [31:0] _GEN_3460; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  wire [31:0] _GEN_3461; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  wire [31:0] _GEN_3462; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  wire [31:0] _GEN_3463; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  wire [31:0] _GEN_3464; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  wire [31:0] _GEN_3465; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  wire [31:0] _GEN_3466; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  wire [31:0] _GEN_3467; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  wire [31:0] _GEN_3468; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  wire [31:0] _GEN_3469; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  wire [31:0] _GEN_3470; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  wire [31:0] _GEN_3471; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  wire [31:0] _GEN_3472; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  wire [31:0] _GEN_3473; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  wire [31:0] _GEN_3474; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  wire [31:0] _GEN_3475; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  wire [31:0] _GEN_3476; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  wire [31:0] _GEN_3477; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  wire [31:0] _GEN_3478; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  wire [31:0] _GEN_3479; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  wire [31:0] _GEN_3480; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  wire [31:0] _GEN_3481; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  wire [31:0] _GEN_3482; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  wire [31:0] _GEN_3483; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  wire [31:0] _GEN_3484; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  wire [31:0] _GEN_3485; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  wire [31:0] _GEN_3486; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  wire [31:0] _GEN_3487; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  wire [31:0] _GEN_3488; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  wire [31:0] _GEN_3489; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  wire [31:0] _GEN_3490; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  wire [31:0] _GEN_3491; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  wire [31:0] _GEN_3492; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  wire [31:0] _GEN_3493; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  wire [31:0] _GEN_3494; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  wire [31:0] _GEN_3495; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  wire [31:0] _GEN_3496; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  wire [31:0] _GEN_3497; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  wire [31:0] _GEN_3498; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  wire [31:0] _GEN_3499; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  wire [31:0] _GEN_3500; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  wire [31:0] _GEN_3501; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  wire [31:0] _GEN_3502; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  wire [31:0] _GEN_3503; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  wire [31:0] _GEN_3504; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  wire [31:0] _GEN_3505; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  wire [31:0] _GEN_3506; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  wire [31:0] _GEN_3507; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  wire [31:0] _GEN_3508; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  wire [31:0] _GEN_3509; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  wire [31:0] _GEN_3510; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  wire [31:0] _GEN_3511; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  wire [31:0] _GEN_3512; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  wire [31:0] _GEN_3513; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  wire [31:0] _GEN_3514; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  wire [31:0] _GEN_3515; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  wire [31:0] _GEN_3516; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  wire [31:0] _GEN_3517; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  wire [31:0] _GEN_3518; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  wire [31:0] _GEN_3519; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  wire [31:0] _GEN_3520; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  wire [31:0] _GEN_3521; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  wire [31:0] _GEN_3522; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  wire [31:0] _GEN_3523; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  wire [31:0] _GEN_3524; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  wire [31:0] _GEN_3525; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  wire [31:0] _GEN_3526; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  wire [31:0] _GEN_3527; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  wire [31:0] _GEN_3528; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  wire [31:0] _GEN_3529; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  wire [31:0] _GEN_3530; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  wire [31:0] _GEN_3531; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  wire [31:0] _GEN_3532; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  wire [31:0] _GEN_3533; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  wire [31:0] _GEN_3534; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  wire [31:0] _GEN_3535; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  wire [31:0] _GEN_3536; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  wire [31:0] _GEN_3537; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  wire [31:0] _GEN_3538; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  wire [31:0] _GEN_3539; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  wire [31:0] _GEN_3540; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  wire [31:0] _GEN_3541; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  wire [31:0] _GEN_3542; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  wire [31:0] _GEN_3543; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  wire [31:0] _GEN_3544; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  wire [31:0] _GEN_3545; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  wire [31:0] _GEN_3546; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  wire [31:0] _GEN_3547; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  wire [31:0] _GEN_3548; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  wire [31:0] _GEN_3549; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  wire [31:0] _GEN_3550; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  wire [31:0] _GEN_3551; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  wire [31:0] _GEN_3552; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  wire [31:0] _GEN_3553; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  wire [31:0] _GEN_3554; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  wire  _T_44820; // @[Debug.scala 1649:18:freechips.rocketchip.system.DefaultRV32Config.fir@168764.10]
  wire  _T_44821; // @[Debug.scala 1649:30:freechips.rocketchip.system.DefaultRV32Config.fir@168765.10]
  wire  _T_44828; // @[Debug.scala 1657:30:freechips.rocketchip.system.DefaultRV32Config.fir@168785.10]
  wire  _T_44831; // @[Debug.scala 1658:13:freechips.rocketchip.system.DefaultRV32Config.fir@168789.12]
  wire  _T_44837; // @[Debug.scala 1671:30:freechips.rocketchip.system.DefaultRV32Config.fir@168810.4]
  wire  _T_44838; // @[Debug.scala 1671:27:freechips.rocketchip.system.DefaultRV32Config.fir@168811.4]
  wire  _T_44840; // @[Debug.scala 1671:49:freechips.rocketchip.system.DefaultRV32Config.fir@168813.4]
  wire  _T_44842; // @[Debug.scala 1671:12:freechips.rocketchip.system.DefaultRV32Config.fir@168815.4]
  wire  _T_44843; // @[Debug.scala 1671:12:freechips.rocketchip.system.DefaultRV32Config.fir@168816.4]
  wire  _GEN_3883; // @[Debug.scala 1389:15:freechips.rocketchip.system.DefaultRV32Config.fir@115473.12]
  wire  _GEN_3884; // @[Debug.scala 1389:15:freechips.rocketchip.system.DefaultRV32Config.fir@115473.12]
  wire  _GEN_3885; // @[Debug.scala 1389:15:freechips.rocketchip.system.DefaultRV32Config.fir@115473.12]
  wire  _GEN_3886; // @[Debug.scala 1389:15:freechips.rocketchip.system.DefaultRV32Config.fir@115473.12]
  wire  _GEN_3892; // @[Debug.scala 1653:15:freechips.rocketchip.system.DefaultRV32Config.fir@168777.14]
  wire  _GEN_3893; // @[Debug.scala 1653:15:freechips.rocketchip.system.DefaultRV32Config.fir@168777.14]
  wire  _GEN_3894; // @[Debug.scala 1653:15:freechips.rocketchip.system.DefaultRV32Config.fir@168777.14]
  wire  _GEN_3895; // @[Debug.scala 1653:15:freechips.rocketchip.system.DefaultRV32Config.fir@168777.14]
  wire  _GEN_3904; // @[Debug.scala 1658:13:freechips.rocketchip.system.DefaultRV32Config.fir@168791.14]
  wire  _GEN_3905; // @[Debug.scala 1658:13:freechips.rocketchip.system.DefaultRV32Config.fir@168791.14]
  wire  _GEN_3906; // @[Debug.scala 1658:13:freechips.rocketchip.system.DefaultRV32Config.fir@168791.14]
  TLMonitor_44 TLMonitor ( // @[Nodes.scala 25:25:freechips.rocketchip.system.DefaultRV32Config.fir@108919.4]
    .clock(TLMonitor_clock),
    .reset(TLMonitor_reset),
    .io_in_a_ready(TLMonitor_io_in_a_ready),
    .io_in_a_valid(TLMonitor_io_in_a_valid),
    .io_in_a_bits_opcode(TLMonitor_io_in_a_bits_opcode),
    .io_in_a_bits_param(TLMonitor_io_in_a_bits_param),
    .io_in_a_bits_size(TLMonitor_io_in_a_bits_size),
    .io_in_a_bits_source(TLMonitor_io_in_a_bits_source),
    .io_in_a_bits_address(TLMonitor_io_in_a_bits_address),
    .io_in_a_bits_mask(TLMonitor_io_in_a_bits_mask),
    .io_in_a_bits_corrupt(TLMonitor_io_in_a_bits_corrupt),
    .io_in_d_ready(TLMonitor_io_in_d_ready),
    .io_in_d_valid(TLMonitor_io_in_d_valid),
    .io_in_d_bits_opcode(TLMonitor_io_in_d_bits_opcode),
    .io_in_d_bits_size(TLMonitor_io_in_d_bits_size),
    .io_in_d_bits_source(TLMonitor_io_in_d_bits_source)
  );
  TLMonitor_45 TLMonitor_1 ( // @[Nodes.scala 25:25:freechips.rocketchip.system.DefaultRV32Config.fir@108944.4]
    .clock(TLMonitor_1_clock),
    .reset(TLMonitor_1_reset),
    .io_in_a_ready(TLMonitor_1_io_in_a_ready),
    .io_in_a_valid(TLMonitor_1_io_in_a_valid),
    .io_in_a_bits_opcode(TLMonitor_1_io_in_a_bits_opcode),
    .io_in_a_bits_param(TLMonitor_1_io_in_a_bits_param),
    .io_in_a_bits_size(TLMonitor_1_io_in_a_bits_size),
    .io_in_a_bits_source(TLMonitor_1_io_in_a_bits_source),
    .io_in_a_bits_address(TLMonitor_1_io_in_a_bits_address),
    .io_in_a_bits_mask(TLMonitor_1_io_in_a_bits_mask),
    .io_in_a_bits_corrupt(TLMonitor_1_io_in_a_bits_corrupt),
    .io_in_d_ready(TLMonitor_1_io_in_d_ready),
    .io_in_d_valid(TLMonitor_1_io_in_d_valid),
    .io_in_d_bits_opcode(TLMonitor_1_io_in_d_bits_opcode),
    .io_in_d_bits_size(TLMonitor_1_io_in_d_bits_size),
    .io_in_d_bits_source(TLMonitor_1_io_in_d_bits_source)
  );
  AsyncResetSynchronizerShiftReg_w1_d3_i0 debug_hartReset_0 ( // @[ShiftReg.scala 45:23:freechips.rocketchip.system.DefaultRV32Config.fir@109292.4]
    .clock(debug_hartReset_0_clock),
    .reset(debug_hartReset_0_reset),
    .io_d(debug_hartReset_0_io_d),
    .io_q(debug_hartReset_0_io_q)
  );
  assign hamaskWrSel_0 = io_innerCtrl_bits_hartsel == 10'h0; // @[Debug.scala 820:61:freechips.rocketchip.system.DefaultRV32Config.fir@109282.4]
  assign _T_13 = ~io_dmactive; // @[Debug.scala 839:11:freechips.rocketchip.system.DefaultRV32Config.fir@109299.4]
  assign _T_16 = io_innerCtrl_ready & io_innerCtrl_valid; // @[Decoupled.scala 40:37:freechips.rocketchip.system.DefaultRV32Config.fir@109306.6]
  assign _T_23 = ~haltedBitRegs_0; // @[package.scala 62:38:freechips.rocketchip.system.DefaultRV32Config.fir@109321.6]
  assign _T_24 = hrDebugInt_0 & _T_23; // @[package.scala 57:72:freechips.rocketchip.system.DefaultRV32Config.fir@109322.6]
  assign hartIsInResetSync_0 = debug_hartReset_0_io_q; // @[ShiftReg.scala 48:24:freechips.rocketchip.system.DefaultRV32Config.fir@109296.4 ShiftReg.scala 48:24:freechips.rocketchip.system.DefaultRV32Config.fir@109297.4]
  assign _T_25 = hartIsInResetSync_0 | _T_24; // @[package.scala 58:75:freechips.rocketchip.system.DefaultRV32Config.fir@109323.6]
  assign _T_26 = hrmaskReg_0 & _T_25; // @[package.scala 57:72:freechips.rocketchip.system.DefaultRV32Config.fir@109324.6]
  assign resumereq = _T_16 & io_innerCtrl_bits_resumereq; // @[Debug.scala 868:41:freechips.rocketchip.system.DefaultRV32Config.fir@109373.4]
  assign _T_306 = ~resumeReqRegs_0; // @[Debug.scala 1227:32:freechips.rocketchip.system.DefaultRV32Config.fir@110286.4]
  assign _T_307 = resumereq & hamaskWrSel_0; // @[Debug.scala 1227:73:freechips.rocketchip.system.DefaultRV32Config.fir@110287.4]
  assign _T_308 = ~_T_307; // @[Debug.scala 1227:61:freechips.rocketchip.system.DefaultRV32Config.fir@110288.4]
  assign resumeAcks_0 = _T_306 & _T_308; // @[Debug.scala 1227:58:freechips.rocketchip.system.DefaultRV32Config.fir@110289.4]
  assign _T_64 = _T_16 & io_innerCtrl_bits_ackhavereset; // @[Debug.scala 902:39:freechips.rocketchip.system.DefaultRV32Config.fir@109438.8]
  assign _T_65 = _T_64 & hamaskWrSel_0; // @[Debug.scala 902:73:freechips.rocketchip.system.DefaultRV32Config.fir@109439.8]
  assign _GEN_34 = _T_65 ? 1'h0 : haveResetBitRegs_0; // @[Debug.scala 902:100:freechips.rocketchip.system.DefaultRV32Config.fir@109440.8]
  assign _GEN_35 = hartIsInResetSync_0 | _GEN_34; // @[Debug.scala 900:49:freechips.rocketchip.system.DefaultRV32Config.fir@109433.6]
  assign haltedStatus_0 = {{31'd0}, haltedBitRegs_0}; // @[Debug.scala 1051:30:freechips.rocketchip.system.DefaultRV32Config.fir@109501.4 Debug.scala 1055:26:freechips.rocketchip.system.DefaultRV32Config.fir@109503.6 Debug.scala 1057:26:freechips.rocketchip.system.DefaultRV32Config.fir@109506.6]
  assign haltedSummary = |haltedStatus_0; // @[Debug.scala 1061:48:freechips.rocketchip.system.DefaultRV32Config.fir@109508.4]
  assign HALTSUM1RdData_haltsum1 = {{31'd0}, haltedSummary}; // @[:freechips.rocketchip.system.DefaultRV32Config.fir@109510.4 :freechips.rocketchip.system.DefaultRV32Config.fir@109511.4]
  assign _T_380 = auto_dmi_in_a_bits_opcode == 3'h4; // @[RegisterRouter.scala 69:36:freechips.rocketchip.system.DefaultRV32Config.fir@110366.4]
  assign _T_2990 = {auto_dmi_in_a_bits_address[7],auto_dmi_in_a_bits_address[5],auto_dmi_in_a_bits_address[4],auto_dmi_in_a_bits_address[3],auto_dmi_in_a_bits_address[2]}; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@113342.4]
  assign _T_385 = auto_dmi_in_a_bits_address[8:2] & 7'h50; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@110382.4]
  assign _T_433 = _T_385 == 7'h0; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@110430.4]
  assign _T_389 = _T_385 == 7'h10; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@110386.4]
  assign _T_407 = _T_385 == 7'h40; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@110404.4]
  assign _T_3564 = auto_dmi_in_a_valid & auto_dmi_in_d_ready; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@114522.4]
  assign _T_3565 = ~_T_380; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@114523.4]
  assign _T_3566 = _T_3564 & _T_3565; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@114524.4]
  assign _T_3035 = 32'h1 << _T_2990; // @[OneHot.scala 58:35:freechips.rocketchip.system.DefaultRV32Config.fir@113387.4]
  assign _T_3598 = _T_3566 & _T_3035[6]; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@114599.4]
  assign _T_3599 = _T_3598 & _T_389; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@114600.4]
  assign _T_465 = auto_dmi_in_a_bits_mask[3] ? 8'hff : 8'h0; // @[Bitwise.scala 72:12:freechips.rocketchip.system.DefaultRV32Config.fir@110466.4]
  assign _T_463 = auto_dmi_in_a_bits_mask[2] ? 8'hff : 8'h0; // @[Bitwise.scala 72:12:freechips.rocketchip.system.DefaultRV32Config.fir@110464.4]
  assign _T_461 = auto_dmi_in_a_bits_mask[1] ? 8'hff : 8'h0; // @[Bitwise.scala 72:12:freechips.rocketchip.system.DefaultRV32Config.fir@110462.4]
  assign _T_459 = auto_dmi_in_a_bits_mask[0] ? 8'hff : 8'h0; // @[Bitwise.scala 72:12:freechips.rocketchip.system.DefaultRV32Config.fir@110460.4]
  assign _T_468 = {_T_465,_T_463,_T_461,_T_459}; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@110469.4]
  assign _T_1929 = &_T_468[10:8]; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@112114.4]
  assign ABSTRACTCSWrEnMaybe = _T_3599 & _T_1929; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@112118.4]
  assign ABSTRACTCSWrEnLegal = ctrlStateReg == 2'h0; // @[Debug.scala 1569:44:freechips.rocketchip.system.DefaultRV32Config.fir@168662.4]
  assign ABSTRACTCSWrEn = ABSTRACTCSWrEnMaybe & ABSTRACTCSWrEnLegal; // @[Debug.scala 1083:51:freechips.rocketchip.system.DefaultRV32Config.fir@109577.4]
  assign ABSTRACTCSWrData_cmderr = auto_dmi_in_a_bits_data[10:8]; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@112119.4]
  assign _T_83 = ~ABSTRACTCSWrData_cmderr; // @[Debug.scala 1103:58:freechips.rocketchip.system.DefaultRV32Config.fir@109617.16]
  assign _T_84 = ABSTRACTCSReg_cmderr & _T_83; // @[Debug.scala 1103:56:freechips.rocketchip.system.DefaultRV32Config.fir@109618.16]
  assign _T_44818 = ctrlStateReg == 2'h1; // @[Debug.scala 1623:30:freechips.rocketchip.system.DefaultRV32Config.fir@168740.6]
  assign commandRegIsAccessRegister = COMMANDRdData_cmdtype == 8'h0; // @[Debug.scala 1584:58:freechips.rocketchip.system.DefaultRV32Config.fir@168691.4]
  assign _T_3960 = {COMMANDRdData_cmdtype,COMMANDRdData_control}; // @[Debug.scala 1415:62:freechips.rocketchip.system.DefaultRV32Config.fir@115544.4]
  assign accessRegisterCommandReg_transfer = _T_3960[17]; // @[Debug.scala 1415:73:freechips.rocketchip.system.DefaultRV32Config.fir@115552.4]
  assign accessRegisterCommandReg_write = _T_3960[16]; // @[Debug.scala 1415:73:freechips.rocketchip.system.DefaultRV32Config.fir@115550.4]
  assign _T_44808 = ~accessRegisterCommandReg_transfer; // @[Debug.scala 1602:19:freechips.rocketchip.system.DefaultRV32Config.fir@168709.8]
  assign accessRegisterCommandReg_regno = _T_3960[15:0]; // @[Debug.scala 1415:73:freechips.rocketchip.system.DefaultRV32Config.fir@115548.4]
  assign _T_44803 = accessRegisterCommandReg_regno >= 16'h1000; // @[Debug.scala 1592:58:freechips.rocketchip.system.DefaultRV32Config.fir@168698.4]
  assign _T_44804 = accessRegisterCommandReg_regno <= 16'h101f; // @[Debug.scala 1592:104:freechips.rocketchip.system.DefaultRV32Config.fir@168699.4]
  assign accessRegIsGPR = _T_44803 & _T_44804; // @[Debug.scala 1592:70:freechips.rocketchip.system.DefaultRV32Config.fir@168700.4]
  assign _T_44809 = _T_44808 | accessRegIsGPR; // @[Debug.scala 1602:54:freechips.rocketchip.system.DefaultRV32Config.fir@168710.8]
  assign _GEN_3623 = _T_44809 ? 1'h0 : 1'h1; // @[Debug.scala 1602:73:freechips.rocketchip.system.DefaultRV32Config.fir@168711.8]
  assign commandRegIsUnsupported = commandRegIsAccessRegister ? _GEN_3623 : 1'h1; // @[Debug.scala 1599:39:freechips.rocketchip.system.DefaultRV32Config.fir@168701.4]
  assign _GEN_3624 = _T_44809 & _T_23; // @[Debug.scala 1602:73:freechips.rocketchip.system.DefaultRV32Config.fir@168711.8]
  assign commandRegBadHaltResume = commandRegIsAccessRegister & _GEN_3624; // @[Debug.scala 1599:39:freechips.rocketchip.system.DefaultRV32Config.fir@168701.4]
  assign _GEN_3640 = commandRegIsUnsupported ? 1'h0 : commandRegBadHaltResume; // @[Debug.scala 1630:38:freechips.rocketchip.system.DefaultRV32Config.fir@168742.8]
  assign _GEN_3653 = _T_44818 & _GEN_3640; // @[Debug.scala 1623:59:freechips.rocketchip.system.DefaultRV32Config.fir@168741.6]
  assign errorHaltResume = ABSTRACTCSWrEnLegal ? 1'h0 : _GEN_3653; // @[Debug.scala 1615:47:freechips.rocketchip.system.DefaultRV32Config.fir@168724.4]
  assign _T_3603 = _T_3566 & _T_3035[7]; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@114613.4]
  assign _T_3604 = _T_3603 & _T_389; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@114614.4]
  assign _T_2649 = &_T_468; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@112936.4]
  assign COMMANDWrEnMaybe = _T_3604 & _T_2649; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@112940.4]
  assign COMMANDWrEn = COMMANDWrEnMaybe & ABSTRACTCSWrEnLegal; // @[Debug.scala 1168:40:freechips.rocketchip.system.DefaultRV32Config.fir@110163.4]
  assign COMMANDWrDataVal = COMMANDWrEnMaybe ? auto_dmi_in_a_bits_data : 32'h0; // @[Debug.scala 265:24:freechips.rocketchip.system.DefaultRV32Config.fir@112944.4]
  assign COMMANDWrData_cmdtype = COMMANDWrDataVal[31:24]; // @[Debug.scala 1163:65:freechips.rocketchip.system.DefaultRV32Config.fir@110152.4]
  assign commandWrIsAccessRegister = COMMANDWrData_cmdtype == 8'h0; // @[Debug.scala 1583:60:freechips.rocketchip.system.DefaultRV32Config.fir@168690.4]
  assign _T_44811 = COMMANDWrEn & commandWrIsAccessRegister; // @[Debug.scala 1608:48:freechips.rocketchip.system.DefaultRV32Config.fir@168717.4]
  assign _T_44812 = ABSTRACTCSReg_cmderr == 3'h0; // @[Debug.scala 1608:103:freechips.rocketchip.system.DefaultRV32Config.fir@168718.4]
  assign wrAccessRegisterCommand = _T_44811 & _T_44812; // @[Debug.scala 1608:78:freechips.rocketchip.system.DefaultRV32Config.fir@168719.4]
  assign _T_3588 = _T_3566 & _T_3035[4]; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@114581.4]
  assign _T_3589 = _T_3588 & _T_433; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@114582.4]
  assign _T_2791 = &_T_468[7:0]; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@113103.4]
  assign dmiAbstractDataWrEnMaybe_0 = _T_3589 & _T_2791; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@113107.4]
  assign _T_3400 = _T_3564 & _T_380; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@114156.4]
  assign _T_3422 = _T_3400 & _T_3035[4]; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@114213.4]
  assign _T_3423 = _T_3422 & _T_433; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@114214.4]
  assign _T_2789 = |_T_468[7:0]; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@113101.4]
  assign dmiAbstractDataRdEn_0 = _T_3423 & _T_2789; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@113105.4]
  assign dmiAbstractDataAccessVec_0 = dmiAbstractDataWrEnMaybe_0 | dmiAbstractDataRdEn_0; // @[Debug.scala 1141:105:freechips.rocketchip.system.DefaultRV32Config.fir@109690.4]
  assign autoexecData_0 = dmiAbstractDataAccessVec_0 & ABSTRACTAUTOReg_autoexecdata[0]; // @[Debug.scala 1152:140:freechips.rocketchip.system.DefaultRV32Config.fir@110072.4]
  assign _T_3648 = _T_3566 & _T_3035[16]; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@114680.4]
  assign _T_3649 = _T_3648 & _T_433; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@114681.4]
  assign dmiProgramBufferWrEnMaybe_0 = _T_3649 & _T_2791; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@111264.4]
  assign _T_3482 = _T_3400 & _T_3035[16]; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@114312.4]
  assign _T_3483 = _T_3482 & _T_433; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@114313.4]
  assign dmiProgramBufferRdEn_0 = _T_3483 & _T_2789; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@111262.4]
  assign dmiProgramBufferAccessVec_0 = dmiProgramBufferWrEnMaybe_0 | dmiProgramBufferRdEn_0; // @[Debug.scala 1144:108:freechips.rocketchip.system.DefaultRV32Config.fir@109828.4]
  assign autoexecProg_0 = dmiProgramBufferAccessVec_0 & ABSTRACTAUTOReg_autoexecprogbuf[0]; // @[Debug.scala 1153:144:freechips.rocketchip.system.DefaultRV32Config.fir@110090.4]
  assign _T_3653 = _T_3566 & _T_3035[17]; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@114691.4]
  assign _T_3654 = _T_3653 & _T_433; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@114692.4]
  assign dmiProgramBufferWrEnMaybe_4 = _T_3654 & _T_2791; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@111028.4]
  assign _T_3487 = _T_3400 & _T_3035[17]; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@114323.4]
  assign _T_3488 = _T_3487 & _T_433; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@114324.4]
  assign dmiProgramBufferRdEn_4 = _T_3488 & _T_2789; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@111026.4]
  assign dmiProgramBufferAccessVec_4 = dmiProgramBufferWrEnMaybe_4 | dmiProgramBufferRdEn_4; // @[Debug.scala 1144:108:freechips.rocketchip.system.DefaultRV32Config.fir@109832.4]
  assign autoexecProg_1 = dmiProgramBufferAccessVec_4 & ABSTRACTAUTOReg_autoexecprogbuf[1]; // @[Debug.scala 1153:144:freechips.rocketchip.system.DefaultRV32Config.fir@110092.4]
  assign _T_276 = autoexecProg_0 | autoexecProg_1; // @[Debug.scala 1155:73:freechips.rocketchip.system.DefaultRV32Config.fir@110122.4]
  assign _T_3658 = _T_3566 & _T_3035[18]; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@114702.4]
  assign _T_3659 = _T_3658 & _T_433; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@114703.4]
  assign dmiProgramBufferWrEnMaybe_8 = _T_3659 & _T_2791; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@111382.4]
  assign _T_3492 = _T_3400 & _T_3035[18]; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@114334.4]
  assign _T_3493 = _T_3492 & _T_433; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@114335.4]
  assign dmiProgramBufferRdEn_8 = _T_3493 & _T_2789; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@111380.4]
  assign dmiProgramBufferAccessVec_8 = dmiProgramBufferWrEnMaybe_8 | dmiProgramBufferRdEn_8; // @[Debug.scala 1144:108:freechips.rocketchip.system.DefaultRV32Config.fir@109836.4]
  assign autoexecProg_2 = dmiProgramBufferAccessVec_8 & ABSTRACTAUTOReg_autoexecprogbuf[2]; // @[Debug.scala 1153:144:freechips.rocketchip.system.DefaultRV32Config.fir@110094.4]
  assign _T_277 = _T_276 | autoexecProg_2; // @[Debug.scala 1155:73:freechips.rocketchip.system.DefaultRV32Config.fir@110123.4]
  assign _T_3663 = _T_3566 & _T_3035[19]; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@114713.4]
  assign _T_3664 = _T_3663 & _T_433; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@114714.4]
  assign dmiProgramBufferWrEnMaybe_12 = _T_3664 & _T_2791; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@112473.4]
  assign _T_3497 = _T_3400 & _T_3035[19]; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@114345.4]
  assign _T_3498 = _T_3497 & _T_433; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@114346.4]
  assign dmiProgramBufferRdEn_12 = _T_3498 & _T_2789; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@112471.4]
  assign dmiProgramBufferAccessVec_12 = dmiProgramBufferWrEnMaybe_12 | dmiProgramBufferRdEn_12; // @[Debug.scala 1144:108:freechips.rocketchip.system.DefaultRV32Config.fir@109840.4]
  assign autoexecProg_3 = dmiProgramBufferAccessVec_12 & ABSTRACTAUTOReg_autoexecprogbuf[3]; // @[Debug.scala 1153:144:freechips.rocketchip.system.DefaultRV32Config.fir@110096.4]
  assign _T_278 = _T_277 | autoexecProg_3; // @[Debug.scala 1155:73:freechips.rocketchip.system.DefaultRV32Config.fir@110124.4]
  assign _T_3668 = _T_3566 & _T_3035[20]; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@114724.4]
  assign _T_3669 = _T_3668 & _T_433; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@114725.4]
  assign dmiProgramBufferWrEnMaybe_16 = _T_3669 & _T_2791; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@112968.4]
  assign _T_3502 = _T_3400 & _T_3035[20]; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@114356.4]
  assign _T_3503 = _T_3502 & _T_433; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@114357.4]
  assign dmiProgramBufferRdEn_16 = _T_3503 & _T_2789; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@112966.4]
  assign dmiProgramBufferAccessVec_16 = dmiProgramBufferWrEnMaybe_16 | dmiProgramBufferRdEn_16; // @[Debug.scala 1144:108:freechips.rocketchip.system.DefaultRV32Config.fir@109844.4]
  assign autoexecProg_4 = dmiProgramBufferAccessVec_16 & ABSTRACTAUTOReg_autoexecprogbuf[4]; // @[Debug.scala 1153:144:freechips.rocketchip.system.DefaultRV32Config.fir@110098.4]
  assign _T_279 = _T_278 | autoexecProg_4; // @[Debug.scala 1155:73:freechips.rocketchip.system.DefaultRV32Config.fir@110125.4]
  assign _T_3673 = _T_3566 & _T_3035[21]; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@114735.4]
  assign _T_3674 = _T_3673 & _T_433; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@114736.4]
  assign dmiProgramBufferWrEnMaybe_20 = _T_3674 & _T_2791; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@110674.4]
  assign _T_3507 = _T_3400 & _T_3035[21]; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@114367.4]
  assign _T_3508 = _T_3507 & _T_433; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@114368.4]
  assign dmiProgramBufferRdEn_20 = _T_3508 & _T_2789; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@110672.4]
  assign dmiProgramBufferAccessVec_20 = dmiProgramBufferWrEnMaybe_20 | dmiProgramBufferRdEn_20; // @[Debug.scala 1144:108:freechips.rocketchip.system.DefaultRV32Config.fir@109848.4]
  assign autoexecProg_5 = dmiProgramBufferAccessVec_20 & ABSTRACTAUTOReg_autoexecprogbuf[5]; // @[Debug.scala 1153:144:freechips.rocketchip.system.DefaultRV32Config.fir@110100.4]
  assign _T_280 = _T_279 | autoexecProg_5; // @[Debug.scala 1155:73:freechips.rocketchip.system.DefaultRV32Config.fir@110126.4]
  assign _T_3678 = _T_3566 & _T_3035[22]; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@114746.4]
  assign _T_3679 = _T_3678 & _T_433; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@114747.4]
  assign dmiProgramBufferWrEnMaybe_24 = _T_3679 & _T_2791; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@110910.4]
  assign _T_3512 = _T_3400 & _T_3035[22]; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@114378.4]
  assign _T_3513 = _T_3512 & _T_433; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@114379.4]
  assign dmiProgramBufferRdEn_24 = _T_3513 & _T_2789; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@110908.4]
  assign dmiProgramBufferAccessVec_24 = dmiProgramBufferWrEnMaybe_24 | dmiProgramBufferRdEn_24; // @[Debug.scala 1144:108:freechips.rocketchip.system.DefaultRV32Config.fir@109852.4]
  assign autoexecProg_6 = dmiProgramBufferAccessVec_24 & ABSTRACTAUTOReg_autoexecprogbuf[6]; // @[Debug.scala 1153:144:freechips.rocketchip.system.DefaultRV32Config.fir@110102.4]
  assign _T_281 = _T_280 | autoexecProg_6; // @[Debug.scala 1155:73:freechips.rocketchip.system.DefaultRV32Config.fir@110127.4]
  assign _T_3683 = _T_3566 & _T_3035[23]; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@114757.4]
  assign _T_3684 = _T_3683 & _T_433; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@114758.4]
  assign dmiProgramBufferWrEnMaybe_28 = _T_3684 & _T_2791; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@112355.4]
  assign _T_3517 = _T_3400 & _T_3035[23]; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@114389.4]
  assign _T_3518 = _T_3517 & _T_433; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@114390.4]
  assign dmiProgramBufferRdEn_28 = _T_3518 & _T_2789; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@112353.4]
  assign dmiProgramBufferAccessVec_28 = dmiProgramBufferWrEnMaybe_28 | dmiProgramBufferRdEn_28; // @[Debug.scala 1144:108:freechips.rocketchip.system.DefaultRV32Config.fir@109856.4]
  assign autoexecProg_7 = dmiProgramBufferAccessVec_28 & ABSTRACTAUTOReg_autoexecprogbuf[7]; // @[Debug.scala 1153:144:freechips.rocketchip.system.DefaultRV32Config.fir@110104.4]
  assign _T_282 = _T_281 | autoexecProg_7; // @[Debug.scala 1155:73:freechips.rocketchip.system.DefaultRV32Config.fir@110128.4]
  assign _T_3688 = _T_3566 & _T_3035[24]; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@114768.4]
  assign _T_3689 = _T_3688 & _T_433; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@114769.4]
  assign dmiProgramBufferWrEnMaybe_32 = _T_3689 & _T_2791; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@112822.4]
  assign _T_3522 = _T_3400 & _T_3035[24]; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@114400.4]
  assign _T_3523 = _T_3522 & _T_433; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@114401.4]
  assign dmiProgramBufferRdEn_32 = _T_3523 & _T_2789; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@112820.4]
  assign dmiProgramBufferAccessVec_32 = dmiProgramBufferWrEnMaybe_32 | dmiProgramBufferRdEn_32; // @[Debug.scala 1144:108:freechips.rocketchip.system.DefaultRV32Config.fir@109860.4]
  assign autoexecProg_8 = dmiProgramBufferAccessVec_32 & ABSTRACTAUTOReg_autoexecprogbuf[8]; // @[Debug.scala 1153:144:freechips.rocketchip.system.DefaultRV32Config.fir@110106.4]
  assign _T_283 = _T_282 | autoexecProg_8; // @[Debug.scala 1155:73:freechips.rocketchip.system.DefaultRV32Config.fir@110129.4]
  assign _T_3693 = _T_3566 & _T_3035[25]; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@114779.4]
  assign _T_3694 = _T_3693 & _T_433; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@114780.4]
  assign dmiProgramBufferWrEnMaybe_36 = _T_3694 & _T_2791; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@111146.4]
  assign _T_3527 = _T_3400 & _T_3035[25]; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@114411.4]
  assign _T_3528 = _T_3527 & _T_433; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@114412.4]
  assign dmiProgramBufferRdEn_36 = _T_3528 & _T_2789; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@111144.4]
  assign dmiProgramBufferAccessVec_36 = dmiProgramBufferWrEnMaybe_36 | dmiProgramBufferRdEn_36; // @[Debug.scala 1144:108:freechips.rocketchip.system.DefaultRV32Config.fir@109864.4]
  assign autoexecProg_9 = dmiProgramBufferAccessVec_36 & ABSTRACTAUTOReg_autoexecprogbuf[9]; // @[Debug.scala 1153:144:freechips.rocketchip.system.DefaultRV32Config.fir@110108.4]
  assign _T_284 = _T_283 | autoexecProg_9; // @[Debug.scala 1155:73:freechips.rocketchip.system.DefaultRV32Config.fir@110130.4]
  assign _T_3698 = _T_3566 & _T_3035[26]; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@114790.4]
  assign _T_3699 = _T_3698 & _T_433; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@114791.4]
  assign dmiProgramBufferWrEnMaybe_40 = _T_3699 & _T_2791; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@110481.4]
  assign _T_3532 = _T_3400 & _T_3035[26]; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@114422.4]
  assign _T_3533 = _T_3532 & _T_433; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@114423.4]
  assign dmiProgramBufferRdEn_40 = _T_3533 & _T_2789; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@110479.4]
  assign dmiProgramBufferAccessVec_40 = dmiProgramBufferWrEnMaybe_40 | dmiProgramBufferRdEn_40; // @[Debug.scala 1144:108:freechips.rocketchip.system.DefaultRV32Config.fir@109868.4]
  assign autoexecProg_10 = dmiProgramBufferAccessVec_40 & ABSTRACTAUTOReg_autoexecprogbuf[10]; // @[Debug.scala 1153:144:freechips.rocketchip.system.DefaultRV32Config.fir@110110.4]
  assign _T_285 = _T_284 | autoexecProg_10; // @[Debug.scala 1155:73:freechips.rocketchip.system.DefaultRV32Config.fir@110131.4]
  assign _T_3703 = _T_3566 & _T_3035[27]; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@114801.4]
  assign _T_3704 = _T_3703 & _T_433; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@114802.4]
  assign dmiProgramBufferWrEnMaybe_44 = _T_3704 & _T_2791; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@112704.4]
  assign _T_3537 = _T_3400 & _T_3035[27]; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@114433.4]
  assign _T_3538 = _T_3537 & _T_433; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@114434.4]
  assign dmiProgramBufferRdEn_44 = _T_3538 & _T_2789; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@112702.4]
  assign dmiProgramBufferAccessVec_44 = dmiProgramBufferWrEnMaybe_44 | dmiProgramBufferRdEn_44; // @[Debug.scala 1144:108:freechips.rocketchip.system.DefaultRV32Config.fir@109872.4]
  assign autoexecProg_11 = dmiProgramBufferAccessVec_44 & ABSTRACTAUTOReg_autoexecprogbuf[11]; // @[Debug.scala 1153:144:freechips.rocketchip.system.DefaultRV32Config.fir@110112.4]
  assign _T_286 = _T_285 | autoexecProg_11; // @[Debug.scala 1155:73:freechips.rocketchip.system.DefaultRV32Config.fir@110132.4]
  assign _T_3708 = _T_3566 & _T_3035[28]; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@114812.4]
  assign _T_3709 = _T_3708 & _T_433; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@114813.4]
  assign dmiProgramBufferWrEnMaybe_48 = _T_3709 & _T_2791; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@112237.4]
  assign _T_3542 = _T_3400 & _T_3035[28]; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@114444.4]
  assign _T_3543 = _T_3542 & _T_433; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@114445.4]
  assign dmiProgramBufferRdEn_48 = _T_3543 & _T_2789; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@112235.4]
  assign dmiProgramBufferAccessVec_48 = dmiProgramBufferWrEnMaybe_48 | dmiProgramBufferRdEn_48; // @[Debug.scala 1144:108:freechips.rocketchip.system.DefaultRV32Config.fir@109876.4]
  assign autoexecProg_12 = dmiProgramBufferAccessVec_48 & ABSTRACTAUTOReg_autoexecprogbuf[12]; // @[Debug.scala 1153:144:freechips.rocketchip.system.DefaultRV32Config.fir@110114.4]
  assign _T_287 = _T_286 | autoexecProg_12; // @[Debug.scala 1155:73:freechips.rocketchip.system.DefaultRV32Config.fir@110133.4]
  assign _T_3713 = _T_3566 & _T_3035[29]; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@114823.4]
  assign _T_3714 = _T_3713 & _T_433; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@114824.4]
  assign dmiProgramBufferWrEnMaybe_52 = _T_3714 & _T_2791; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@111500.4]
  assign _T_3547 = _T_3400 & _T_3035[29]; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@114455.4]
  assign _T_3548 = _T_3547 & _T_433; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@114456.4]
  assign dmiProgramBufferRdEn_52 = _T_3548 & _T_2789; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@111498.4]
  assign dmiProgramBufferAccessVec_52 = dmiProgramBufferWrEnMaybe_52 | dmiProgramBufferRdEn_52; // @[Debug.scala 1144:108:freechips.rocketchip.system.DefaultRV32Config.fir@109880.4]
  assign autoexecProg_13 = dmiProgramBufferAccessVec_52 & ABSTRACTAUTOReg_autoexecprogbuf[13]; // @[Debug.scala 1153:144:freechips.rocketchip.system.DefaultRV32Config.fir@110116.4]
  assign _T_288 = _T_287 | autoexecProg_13; // @[Debug.scala 1155:73:freechips.rocketchip.system.DefaultRV32Config.fir@110134.4]
  assign _T_3718 = _T_3566 & _T_3035[30]; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@114834.4]
  assign _T_3719 = _T_3718 & _T_433; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@114835.4]
  assign dmiProgramBufferWrEnMaybe_56 = _T_3719 & _T_2791; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@110792.4]
  assign _T_3552 = _T_3400 & _T_3035[30]; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@114466.4]
  assign _T_3553 = _T_3552 & _T_433; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@114467.4]
  assign dmiProgramBufferRdEn_56 = _T_3553 & _T_2789; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@110790.4]
  assign dmiProgramBufferAccessVec_56 = dmiProgramBufferWrEnMaybe_56 | dmiProgramBufferRdEn_56; // @[Debug.scala 1144:108:freechips.rocketchip.system.DefaultRV32Config.fir@109884.4]
  assign autoexecProg_14 = dmiProgramBufferAccessVec_56 & ABSTRACTAUTOReg_autoexecprogbuf[14]; // @[Debug.scala 1153:144:freechips.rocketchip.system.DefaultRV32Config.fir@110118.4]
  assign _T_289 = _T_288 | autoexecProg_14; // @[Debug.scala 1155:73:freechips.rocketchip.system.DefaultRV32Config.fir@110135.4]
  assign _T_3723 = _T_3566 & _T_3035[31]; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@114845.4]
  assign _T_3724 = _T_3723 & _T_433; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@114846.4]
  assign dmiProgramBufferWrEnMaybe_60 = _T_3724 & _T_2791; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@113225.4]
  assign _T_3557 = _T_3400 & _T_3035[31]; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@114477.4]
  assign _T_3558 = _T_3557 & _T_433; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@114478.4]
  assign dmiProgramBufferRdEn_60 = _T_3558 & _T_2789; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@113223.4]
  assign dmiProgramBufferAccessVec_60 = dmiProgramBufferWrEnMaybe_60 | dmiProgramBufferRdEn_60; // @[Debug.scala 1144:108:freechips.rocketchip.system.DefaultRV32Config.fir@109888.4]
  assign autoexecProg_15 = dmiProgramBufferAccessVec_60 & ABSTRACTAUTOReg_autoexecprogbuf[15]; // @[Debug.scala 1153:144:freechips.rocketchip.system.DefaultRV32Config.fir@110120.4]
  assign _T_290 = _T_289 | autoexecProg_15; // @[Debug.scala 1155:73:freechips.rocketchip.system.DefaultRV32Config.fir@110136.4]
  assign autoexec = autoexecData_0 | _T_290; // @[Debug.scala 1155:48:freechips.rocketchip.system.DefaultRV32Config.fir@110137.4]
  assign _T_44813 = autoexec & commandRegIsAccessRegister; // @[Debug.scala 1609:48:freechips.rocketchip.system.DefaultRV32Config.fir@168720.4]
  assign regAccessRegisterCommand = _T_44813 & _T_44812; // @[Debug.scala 1609:78:freechips.rocketchip.system.DefaultRV32Config.fir@168722.4]
  assign _T_44816 = wrAccessRegisterCommand | regAccessRegisterCommand; // @[Debug.scala 1616:37:freechips.rocketchip.system.DefaultRV32Config.fir@168725.6]
  assign _T_44802 = ~commandWrIsAccessRegister; // @[Debug.scala 1586:49:freechips.rocketchip.system.DefaultRV32Config.fir@168692.4]
  assign commandWrIsUnsupported = COMMANDWrEn & _T_44802; // @[Debug.scala 1586:46:freechips.rocketchip.system.DefaultRV32Config.fir@168693.4]
  assign _T_44817 = autoexec & commandRegIsUnsupported; // @[Debug.scala 1620:28:freechips.rocketchip.system.DefaultRV32Config.fir@168734.10]
  assign _GEN_3630 = commandWrIsUnsupported | _T_44817; // @[Debug.scala 1618:43:freechips.rocketchip.system.DefaultRV32Config.fir@168730.8]
  assign _GEN_3632 = _T_44816 ? 1'h0 : _GEN_3630; // @[Debug.scala 1616:66:freechips.rocketchip.system.DefaultRV32Config.fir@168726.6]
  assign _GEN_3651 = _T_44818 & commandRegIsUnsupported; // @[Debug.scala 1623:59:freechips.rocketchip.system.DefaultRV32Config.fir@168741.6]
  assign errorUnsupported = ABSTRACTCSWrEnLegal ? _GEN_3632 : _GEN_3651; // @[Debug.scala 1615:47:freechips.rocketchip.system.DefaultRV32Config.fir@168724.4]
  assign _T_44819 = ctrlStateReg == 2'h2; // @[Debug.scala 1644:30:freechips.rocketchip.system.DefaultRV32Config.fir@168762.8]
  assign _T_6050 = auto_tl_in_a_bits_opcode == 3'h4; // @[RegisterRouter.scala 69:36:freechips.rocketchip.system.DefaultRV32Config.fir@117696.4]
  assign _T_33453 = {auto_tl_in_a_bits_address[10],auto_tl_in_a_bits_address[9],auto_tl_in_a_bits_address[8],auto_tl_in_a_bits_address[7],auto_tl_in_a_bits_address[6],auto_tl_in_a_bits_address[5],auto_tl_in_a_bits_address[4],auto_tl_in_a_bits_address[3],auto_tl_in_a_bits_address[2]}; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@145326.4]
  assign _T_6055 = auto_tl_in_a_bits_address[11:2] & 10'h200; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@117712.4]
  assign _T_6089 = _T_6055 == 10'h0; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@117746.4]
  assign _T_6609 = _T_6055 == 10'h200; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@118266.4]
  assign _T_42194 = auto_tl_in_a_valid & auto_tl_in_d_ready; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@162227.4]
  assign _T_42195 = ~_T_6050; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@162228.4]
  assign _T_42196 = _T_42194 & _T_42195; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@162229.4]
  assign _T_33985 = 512'h1 << _T_33453; // @[OneHot.scala 58:35:freechips.rocketchip.system.DefaultRV32Config.fir@145858.4]
  assign _T_42533 = _T_42196 & _T_33985[67]; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@162788.4]
  assign _T_42534 = _T_42533 & _T_6089; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@162789.4]
  assign _T_6689 = auto_tl_in_a_bits_mask[3] ? 8'hff : 8'h0; // @[Bitwise.scala 72:12:freechips.rocketchip.system.DefaultRV32Config.fir@118350.4]
  assign _T_6687 = auto_tl_in_a_bits_mask[2] ? 8'hff : 8'h0; // @[Bitwise.scala 72:12:freechips.rocketchip.system.DefaultRV32Config.fir@118348.4]
  assign _T_6685 = auto_tl_in_a_bits_mask[1] ? 8'hff : 8'h0; // @[Bitwise.scala 72:12:freechips.rocketchip.system.DefaultRV32Config.fir@118346.4]
  assign _T_6683 = auto_tl_in_a_bits_mask[0] ? 8'hff : 8'h0; // @[Bitwise.scala 72:12:freechips.rocketchip.system.DefaultRV32Config.fir@118344.4]
  assign _T_6692 = {_T_6689,_T_6687,_T_6685,_T_6683}; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@118353.4]
  assign _T_25711 = &_T_6692[9:0]; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@137522.4]
  assign hartExceptionWrEn = _T_42534 & _T_25711; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@137526.4]
  assign _GEN_3649 = _T_44819 & hartExceptionWrEn; // @[Debug.scala 1644:51:freechips.rocketchip.system.DefaultRV32Config.fir@168763.8]
  assign _GEN_3655 = _T_44818 ? 1'h0 : _GEN_3649; // @[Debug.scala 1623:59:freechips.rocketchip.system.DefaultRV32Config.fir@168741.6]
  assign errorException = ABSTRACTCSWrEnLegal ? 1'h0 : _GEN_3655; // @[Debug.scala 1615:47:freechips.rocketchip.system.DefaultRV32Config.fir@168724.4]
  assign _T_44785 = ~ABSTRACTCSWrEnLegal; // @[Debug.scala 1575:45:freechips.rocketchip.system.DefaultRV32Config.fir@168672.4]
  assign _T_44786 = ABSTRACTCSWrEnMaybe & _T_44785; // @[Debug.scala 1575:42:freechips.rocketchip.system.DefaultRV32Config.fir@168673.4]
  assign _T_3608 = _T_3566 & _T_3035[8]; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@114621.4]
  assign _T_3609 = _T_3608 & _T_389; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@114622.4]
  assign _T_574 = &_T_468[0]; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@110595.4]
  assign autoexecdataWrEnMaybe = _T_3609 & _T_574; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@110599.4]
  assign _T_44788 = autoexecdataWrEnMaybe & _T_44785; // @[Debug.scala 1576:42:freechips.rocketchip.system.DefaultRV32Config.fir@168675.4]
  assign _T_44789 = _T_44786 | _T_44788; // @[Debug.scala 1575:74:freechips.rocketchip.system.DefaultRV32Config.fir@168676.4]
  assign _T_620 = &_T_468[31:16]; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@110643.4]
  assign autoexecprogbufWrEnMaybe = _T_3609 & _T_620; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@110647.4]
  assign _T_44791 = autoexecprogbufWrEnMaybe & _T_44785; // @[Debug.scala 1577:44:freechips.rocketchip.system.DefaultRV32Config.fir@168678.4]
  assign _T_44792 = _T_44789 | _T_44791; // @[Debug.scala 1576:74:freechips.rocketchip.system.DefaultRV32Config.fir@168679.4]
  assign _T_44794 = COMMANDWrEnMaybe & _T_44785; // @[Debug.scala 1578:42:freechips.rocketchip.system.DefaultRV32Config.fir@168681.4]
  assign _T_44795 = _T_44792 | _T_44794; // @[Debug.scala 1577:74:freechips.rocketchip.system.DefaultRV32Config.fir@168682.4]
  assign _T_2814 = &_T_468[15:8]; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@113131.4]
  assign dmiAbstractDataWrEnMaybe_1 = _T_3589 & _T_2814; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@113135.4]
  assign _T_2812 = |_T_468[15:8]; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@113129.4]
  assign dmiAbstractDataRdEn_1 = _T_3423 & _T_2812; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@113133.4]
  assign dmiAbstractDataAccessVec_1 = dmiAbstractDataWrEnMaybe_1 | dmiAbstractDataRdEn_1; // @[Debug.scala 1141:105:freechips.rocketchip.system.DefaultRV32Config.fir@109691.4]
  assign _T_165 = dmiAbstractDataAccessVec_0 | dmiAbstractDataAccessVec_1; // @[Debug.scala 1146:68:freechips.rocketchip.system.DefaultRV32Config.fir@109956.4]
  assign _T_2839 = &_T_468[23:16]; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@113161.4]
  assign dmiAbstractDataWrEnMaybe_2 = _T_3589 & _T_2839; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@113165.4]
  assign _T_2837 = |_T_468[23:16]; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@113159.4]
  assign dmiAbstractDataRdEn_2 = _T_3423 & _T_2837; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@113163.4]
  assign dmiAbstractDataAccessVec_2 = dmiAbstractDataWrEnMaybe_2 | dmiAbstractDataRdEn_2; // @[Debug.scala 1141:105:freechips.rocketchip.system.DefaultRV32Config.fir@109692.4]
  assign _T_166 = _T_165 | dmiAbstractDataAccessVec_2; // @[Debug.scala 1146:68:freechips.rocketchip.system.DefaultRV32Config.fir@109957.4]
  assign _T_2864 = &_T_468[31:24]; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@113191.4]
  assign dmiAbstractDataWrEnMaybe_3 = _T_3589 & _T_2864; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@113195.4]
  assign _T_2862 = |_T_468[31:24]; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@113189.4]
  assign dmiAbstractDataRdEn_3 = _T_3423 & _T_2862; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@113193.4]
  assign dmiAbstractDataAccessVec_3 = dmiAbstractDataWrEnMaybe_3 | dmiAbstractDataRdEn_3; // @[Debug.scala 1141:105:freechips.rocketchip.system.DefaultRV32Config.fir@109693.4]
  assign dmiAbstractDataAccess = _T_166 | dmiAbstractDataAccessVec_3; // @[Debug.scala 1146:68:freechips.rocketchip.system.DefaultRV32Config.fir@109958.4]
  assign _T_44797 = dmiAbstractDataAccess & _T_44785; // @[Debug.scala 1579:42:freechips.rocketchip.system.DefaultRV32Config.fir@168684.4]
  assign _T_44798 = _T_44795 | _T_44797; // @[Debug.scala 1578:74:freechips.rocketchip.system.DefaultRV32Config.fir@168685.4]
  assign dmiProgramBufferWrEnMaybe_1 = _T_3649 & _T_2814; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@111292.4]
  assign dmiProgramBufferRdEn_1 = _T_3483 & _T_2812; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@111290.4]
  assign dmiProgramBufferAccessVec_1 = dmiProgramBufferWrEnMaybe_1 | dmiProgramBufferRdEn_1; // @[Debug.scala 1144:108:freechips.rocketchip.system.DefaultRV32Config.fir@109829.4]
  assign _T_167 = dmiProgramBufferAccessVec_0 | dmiProgramBufferAccessVec_1; // @[Debug.scala 1147:69:freechips.rocketchip.system.DefaultRV32Config.fir@109959.4]
  assign dmiProgramBufferWrEnMaybe_2 = _T_3649 & _T_2839; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@111322.4]
  assign dmiProgramBufferRdEn_2 = _T_3483 & _T_2837; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@111320.4]
  assign dmiProgramBufferAccessVec_2 = dmiProgramBufferWrEnMaybe_2 | dmiProgramBufferRdEn_2; // @[Debug.scala 1144:108:freechips.rocketchip.system.DefaultRV32Config.fir@109830.4]
  assign _T_168 = _T_167 | dmiProgramBufferAccessVec_2; // @[Debug.scala 1147:69:freechips.rocketchip.system.DefaultRV32Config.fir@109960.4]
  assign dmiProgramBufferWrEnMaybe_3 = _T_3649 & _T_2864; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@111352.4]
  assign dmiProgramBufferRdEn_3 = _T_3483 & _T_2862; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@111350.4]
  assign dmiProgramBufferAccessVec_3 = dmiProgramBufferWrEnMaybe_3 | dmiProgramBufferRdEn_3; // @[Debug.scala 1144:108:freechips.rocketchip.system.DefaultRV32Config.fir@109831.4]
  assign _T_169 = _T_168 | dmiProgramBufferAccessVec_3; // @[Debug.scala 1147:69:freechips.rocketchip.system.DefaultRV32Config.fir@109961.4]
  assign _T_170 = _T_169 | dmiProgramBufferAccessVec_4; // @[Debug.scala 1147:69:freechips.rocketchip.system.DefaultRV32Config.fir@109962.4]
  assign dmiProgramBufferWrEnMaybe_5 = _T_3654 & _T_2814; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@111056.4]
  assign dmiProgramBufferRdEn_5 = _T_3488 & _T_2812; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@111054.4]
  assign dmiProgramBufferAccessVec_5 = dmiProgramBufferWrEnMaybe_5 | dmiProgramBufferRdEn_5; // @[Debug.scala 1144:108:freechips.rocketchip.system.DefaultRV32Config.fir@109833.4]
  assign _T_171 = _T_170 | dmiProgramBufferAccessVec_5; // @[Debug.scala 1147:69:freechips.rocketchip.system.DefaultRV32Config.fir@109963.4]
  assign dmiProgramBufferWrEnMaybe_6 = _T_3654 & _T_2839; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@111086.4]
  assign dmiProgramBufferRdEn_6 = _T_3488 & _T_2837; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@111084.4]
  assign dmiProgramBufferAccessVec_6 = dmiProgramBufferWrEnMaybe_6 | dmiProgramBufferRdEn_6; // @[Debug.scala 1144:108:freechips.rocketchip.system.DefaultRV32Config.fir@109834.4]
  assign _T_172 = _T_171 | dmiProgramBufferAccessVec_6; // @[Debug.scala 1147:69:freechips.rocketchip.system.DefaultRV32Config.fir@109964.4]
  assign dmiProgramBufferWrEnMaybe_7 = _T_3654 & _T_2864; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@111116.4]
  assign dmiProgramBufferRdEn_7 = _T_3488 & _T_2862; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@111114.4]
  assign dmiProgramBufferAccessVec_7 = dmiProgramBufferWrEnMaybe_7 | dmiProgramBufferRdEn_7; // @[Debug.scala 1144:108:freechips.rocketchip.system.DefaultRV32Config.fir@109835.4]
  assign _T_173 = _T_172 | dmiProgramBufferAccessVec_7; // @[Debug.scala 1147:69:freechips.rocketchip.system.DefaultRV32Config.fir@109965.4]
  assign _T_174 = _T_173 | dmiProgramBufferAccessVec_8; // @[Debug.scala 1147:69:freechips.rocketchip.system.DefaultRV32Config.fir@109966.4]
  assign dmiProgramBufferWrEnMaybe_9 = _T_3659 & _T_2814; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@111410.4]
  assign dmiProgramBufferRdEn_9 = _T_3493 & _T_2812; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@111408.4]
  assign dmiProgramBufferAccessVec_9 = dmiProgramBufferWrEnMaybe_9 | dmiProgramBufferRdEn_9; // @[Debug.scala 1144:108:freechips.rocketchip.system.DefaultRV32Config.fir@109837.4]
  assign _T_175 = _T_174 | dmiProgramBufferAccessVec_9; // @[Debug.scala 1147:69:freechips.rocketchip.system.DefaultRV32Config.fir@109967.4]
  assign dmiProgramBufferWrEnMaybe_10 = _T_3659 & _T_2839; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@111440.4]
  assign dmiProgramBufferRdEn_10 = _T_3493 & _T_2837; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@111438.4]
  assign dmiProgramBufferAccessVec_10 = dmiProgramBufferWrEnMaybe_10 | dmiProgramBufferRdEn_10; // @[Debug.scala 1144:108:freechips.rocketchip.system.DefaultRV32Config.fir@109838.4]
  assign _T_176 = _T_175 | dmiProgramBufferAccessVec_10; // @[Debug.scala 1147:69:freechips.rocketchip.system.DefaultRV32Config.fir@109968.4]
  assign dmiProgramBufferWrEnMaybe_11 = _T_3659 & _T_2864; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@111470.4]
  assign dmiProgramBufferRdEn_11 = _T_3493 & _T_2862; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@111468.4]
  assign dmiProgramBufferAccessVec_11 = dmiProgramBufferWrEnMaybe_11 | dmiProgramBufferRdEn_11; // @[Debug.scala 1144:108:freechips.rocketchip.system.DefaultRV32Config.fir@109839.4]
  assign _T_177 = _T_176 | dmiProgramBufferAccessVec_11; // @[Debug.scala 1147:69:freechips.rocketchip.system.DefaultRV32Config.fir@109969.4]
  assign _T_178 = _T_177 | dmiProgramBufferAccessVec_12; // @[Debug.scala 1147:69:freechips.rocketchip.system.DefaultRV32Config.fir@109970.4]
  assign dmiProgramBufferWrEnMaybe_13 = _T_3664 & _T_2814; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@112501.4]
  assign dmiProgramBufferRdEn_13 = _T_3498 & _T_2812; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@112499.4]
  assign dmiProgramBufferAccessVec_13 = dmiProgramBufferWrEnMaybe_13 | dmiProgramBufferRdEn_13; // @[Debug.scala 1144:108:freechips.rocketchip.system.DefaultRV32Config.fir@109841.4]
  assign _T_179 = _T_178 | dmiProgramBufferAccessVec_13; // @[Debug.scala 1147:69:freechips.rocketchip.system.DefaultRV32Config.fir@109971.4]
  assign dmiProgramBufferWrEnMaybe_14 = _T_3664 & _T_2839; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@112531.4]
  assign dmiProgramBufferRdEn_14 = _T_3498 & _T_2837; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@112529.4]
  assign dmiProgramBufferAccessVec_14 = dmiProgramBufferWrEnMaybe_14 | dmiProgramBufferRdEn_14; // @[Debug.scala 1144:108:freechips.rocketchip.system.DefaultRV32Config.fir@109842.4]
  assign _T_180 = _T_179 | dmiProgramBufferAccessVec_14; // @[Debug.scala 1147:69:freechips.rocketchip.system.DefaultRV32Config.fir@109972.4]
  assign dmiProgramBufferWrEnMaybe_15 = _T_3664 & _T_2864; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@112561.4]
  assign dmiProgramBufferRdEn_15 = _T_3498 & _T_2862; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@112559.4]
  assign dmiProgramBufferAccessVec_15 = dmiProgramBufferWrEnMaybe_15 | dmiProgramBufferRdEn_15; // @[Debug.scala 1144:108:freechips.rocketchip.system.DefaultRV32Config.fir@109843.4]
  assign _T_181 = _T_180 | dmiProgramBufferAccessVec_15; // @[Debug.scala 1147:69:freechips.rocketchip.system.DefaultRV32Config.fir@109973.4]
  assign _T_182 = _T_181 | dmiProgramBufferAccessVec_16; // @[Debug.scala 1147:69:freechips.rocketchip.system.DefaultRV32Config.fir@109974.4]
  assign dmiProgramBufferWrEnMaybe_17 = _T_3669 & _T_2814; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@112996.4]
  assign dmiProgramBufferRdEn_17 = _T_3503 & _T_2812; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@112994.4]
  assign dmiProgramBufferAccessVec_17 = dmiProgramBufferWrEnMaybe_17 | dmiProgramBufferRdEn_17; // @[Debug.scala 1144:108:freechips.rocketchip.system.DefaultRV32Config.fir@109845.4]
  assign _T_183 = _T_182 | dmiProgramBufferAccessVec_17; // @[Debug.scala 1147:69:freechips.rocketchip.system.DefaultRV32Config.fir@109975.4]
  assign dmiProgramBufferWrEnMaybe_18 = _T_3669 & _T_2839; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@113026.4]
  assign dmiProgramBufferRdEn_18 = _T_3503 & _T_2837; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@113024.4]
  assign dmiProgramBufferAccessVec_18 = dmiProgramBufferWrEnMaybe_18 | dmiProgramBufferRdEn_18; // @[Debug.scala 1144:108:freechips.rocketchip.system.DefaultRV32Config.fir@109846.4]
  assign _T_184 = _T_183 | dmiProgramBufferAccessVec_18; // @[Debug.scala 1147:69:freechips.rocketchip.system.DefaultRV32Config.fir@109976.4]
  assign dmiProgramBufferWrEnMaybe_19 = _T_3669 & _T_2864; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@113056.4]
  assign dmiProgramBufferRdEn_19 = _T_3503 & _T_2862; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@113054.4]
  assign dmiProgramBufferAccessVec_19 = dmiProgramBufferWrEnMaybe_19 | dmiProgramBufferRdEn_19; // @[Debug.scala 1144:108:freechips.rocketchip.system.DefaultRV32Config.fir@109847.4]
  assign _T_185 = _T_184 | dmiProgramBufferAccessVec_19; // @[Debug.scala 1147:69:freechips.rocketchip.system.DefaultRV32Config.fir@109977.4]
  assign _T_186 = _T_185 | dmiProgramBufferAccessVec_20; // @[Debug.scala 1147:69:freechips.rocketchip.system.DefaultRV32Config.fir@109978.4]
  assign dmiProgramBufferWrEnMaybe_21 = _T_3674 & _T_2814; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@110702.4]
  assign dmiProgramBufferRdEn_21 = _T_3508 & _T_2812; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@110700.4]
  assign dmiProgramBufferAccessVec_21 = dmiProgramBufferWrEnMaybe_21 | dmiProgramBufferRdEn_21; // @[Debug.scala 1144:108:freechips.rocketchip.system.DefaultRV32Config.fir@109849.4]
  assign _T_187 = _T_186 | dmiProgramBufferAccessVec_21; // @[Debug.scala 1147:69:freechips.rocketchip.system.DefaultRV32Config.fir@109979.4]
  assign dmiProgramBufferWrEnMaybe_22 = _T_3674 & _T_2839; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@110732.4]
  assign dmiProgramBufferRdEn_22 = _T_3508 & _T_2837; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@110730.4]
  assign dmiProgramBufferAccessVec_22 = dmiProgramBufferWrEnMaybe_22 | dmiProgramBufferRdEn_22; // @[Debug.scala 1144:108:freechips.rocketchip.system.DefaultRV32Config.fir@109850.4]
  assign _T_188 = _T_187 | dmiProgramBufferAccessVec_22; // @[Debug.scala 1147:69:freechips.rocketchip.system.DefaultRV32Config.fir@109980.4]
  assign dmiProgramBufferWrEnMaybe_23 = _T_3674 & _T_2864; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@110762.4]
  assign dmiProgramBufferRdEn_23 = _T_3508 & _T_2862; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@110760.4]
  assign dmiProgramBufferAccessVec_23 = dmiProgramBufferWrEnMaybe_23 | dmiProgramBufferRdEn_23; // @[Debug.scala 1144:108:freechips.rocketchip.system.DefaultRV32Config.fir@109851.4]
  assign _T_189 = _T_188 | dmiProgramBufferAccessVec_23; // @[Debug.scala 1147:69:freechips.rocketchip.system.DefaultRV32Config.fir@109981.4]
  assign _T_190 = _T_189 | dmiProgramBufferAccessVec_24; // @[Debug.scala 1147:69:freechips.rocketchip.system.DefaultRV32Config.fir@109982.4]
  assign dmiProgramBufferWrEnMaybe_25 = _T_3679 & _T_2814; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@110938.4]
  assign dmiProgramBufferRdEn_25 = _T_3513 & _T_2812; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@110936.4]
  assign dmiProgramBufferAccessVec_25 = dmiProgramBufferWrEnMaybe_25 | dmiProgramBufferRdEn_25; // @[Debug.scala 1144:108:freechips.rocketchip.system.DefaultRV32Config.fir@109853.4]
  assign _T_191 = _T_190 | dmiProgramBufferAccessVec_25; // @[Debug.scala 1147:69:freechips.rocketchip.system.DefaultRV32Config.fir@109983.4]
  assign dmiProgramBufferWrEnMaybe_26 = _T_3679 & _T_2839; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@110968.4]
  assign dmiProgramBufferRdEn_26 = _T_3513 & _T_2837; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@110966.4]
  assign dmiProgramBufferAccessVec_26 = dmiProgramBufferWrEnMaybe_26 | dmiProgramBufferRdEn_26; // @[Debug.scala 1144:108:freechips.rocketchip.system.DefaultRV32Config.fir@109854.4]
  assign _T_192 = _T_191 | dmiProgramBufferAccessVec_26; // @[Debug.scala 1147:69:freechips.rocketchip.system.DefaultRV32Config.fir@109984.4]
  assign dmiProgramBufferWrEnMaybe_27 = _T_3679 & _T_2864; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@110998.4]
  assign dmiProgramBufferRdEn_27 = _T_3513 & _T_2862; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@110996.4]
  assign dmiProgramBufferAccessVec_27 = dmiProgramBufferWrEnMaybe_27 | dmiProgramBufferRdEn_27; // @[Debug.scala 1144:108:freechips.rocketchip.system.DefaultRV32Config.fir@109855.4]
  assign _T_193 = _T_192 | dmiProgramBufferAccessVec_27; // @[Debug.scala 1147:69:freechips.rocketchip.system.DefaultRV32Config.fir@109985.4]
  assign _T_194 = _T_193 | dmiProgramBufferAccessVec_28; // @[Debug.scala 1147:69:freechips.rocketchip.system.DefaultRV32Config.fir@109986.4]
  assign dmiProgramBufferWrEnMaybe_29 = _T_3684 & _T_2814; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@112383.4]
  assign dmiProgramBufferRdEn_29 = _T_3518 & _T_2812; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@112381.4]
  assign dmiProgramBufferAccessVec_29 = dmiProgramBufferWrEnMaybe_29 | dmiProgramBufferRdEn_29; // @[Debug.scala 1144:108:freechips.rocketchip.system.DefaultRV32Config.fir@109857.4]
  assign _T_195 = _T_194 | dmiProgramBufferAccessVec_29; // @[Debug.scala 1147:69:freechips.rocketchip.system.DefaultRV32Config.fir@109987.4]
  assign dmiProgramBufferWrEnMaybe_30 = _T_3684 & _T_2839; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@112413.4]
  assign dmiProgramBufferRdEn_30 = _T_3518 & _T_2837; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@112411.4]
  assign dmiProgramBufferAccessVec_30 = dmiProgramBufferWrEnMaybe_30 | dmiProgramBufferRdEn_30; // @[Debug.scala 1144:108:freechips.rocketchip.system.DefaultRV32Config.fir@109858.4]
  assign _T_196 = _T_195 | dmiProgramBufferAccessVec_30; // @[Debug.scala 1147:69:freechips.rocketchip.system.DefaultRV32Config.fir@109988.4]
  assign dmiProgramBufferWrEnMaybe_31 = _T_3684 & _T_2864; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@112443.4]
  assign dmiProgramBufferRdEn_31 = _T_3518 & _T_2862; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@112441.4]
  assign dmiProgramBufferAccessVec_31 = dmiProgramBufferWrEnMaybe_31 | dmiProgramBufferRdEn_31; // @[Debug.scala 1144:108:freechips.rocketchip.system.DefaultRV32Config.fir@109859.4]
  assign _T_197 = _T_196 | dmiProgramBufferAccessVec_31; // @[Debug.scala 1147:69:freechips.rocketchip.system.DefaultRV32Config.fir@109989.4]
  assign _T_198 = _T_197 | dmiProgramBufferAccessVec_32; // @[Debug.scala 1147:69:freechips.rocketchip.system.DefaultRV32Config.fir@109990.4]
  assign dmiProgramBufferWrEnMaybe_33 = _T_3689 & _T_2814; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@112850.4]
  assign dmiProgramBufferRdEn_33 = _T_3523 & _T_2812; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@112848.4]
  assign dmiProgramBufferAccessVec_33 = dmiProgramBufferWrEnMaybe_33 | dmiProgramBufferRdEn_33; // @[Debug.scala 1144:108:freechips.rocketchip.system.DefaultRV32Config.fir@109861.4]
  assign _T_199 = _T_198 | dmiProgramBufferAccessVec_33; // @[Debug.scala 1147:69:freechips.rocketchip.system.DefaultRV32Config.fir@109991.4]
  assign dmiProgramBufferWrEnMaybe_34 = _T_3689 & _T_2839; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@112880.4]
  assign dmiProgramBufferRdEn_34 = _T_3523 & _T_2837; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@112878.4]
  assign dmiProgramBufferAccessVec_34 = dmiProgramBufferWrEnMaybe_34 | dmiProgramBufferRdEn_34; // @[Debug.scala 1144:108:freechips.rocketchip.system.DefaultRV32Config.fir@109862.4]
  assign _T_200 = _T_199 | dmiProgramBufferAccessVec_34; // @[Debug.scala 1147:69:freechips.rocketchip.system.DefaultRV32Config.fir@109992.4]
  assign dmiProgramBufferWrEnMaybe_35 = _T_3689 & _T_2864; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@112910.4]
  assign dmiProgramBufferRdEn_35 = _T_3523 & _T_2862; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@112908.4]
  assign dmiProgramBufferAccessVec_35 = dmiProgramBufferWrEnMaybe_35 | dmiProgramBufferRdEn_35; // @[Debug.scala 1144:108:freechips.rocketchip.system.DefaultRV32Config.fir@109863.4]
  assign _T_201 = _T_200 | dmiProgramBufferAccessVec_35; // @[Debug.scala 1147:69:freechips.rocketchip.system.DefaultRV32Config.fir@109993.4]
  assign _T_202 = _T_201 | dmiProgramBufferAccessVec_36; // @[Debug.scala 1147:69:freechips.rocketchip.system.DefaultRV32Config.fir@109994.4]
  assign dmiProgramBufferWrEnMaybe_37 = _T_3694 & _T_2814; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@111174.4]
  assign dmiProgramBufferRdEn_37 = _T_3528 & _T_2812; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@111172.4]
  assign dmiProgramBufferAccessVec_37 = dmiProgramBufferWrEnMaybe_37 | dmiProgramBufferRdEn_37; // @[Debug.scala 1144:108:freechips.rocketchip.system.DefaultRV32Config.fir@109865.4]
  assign _T_203 = _T_202 | dmiProgramBufferAccessVec_37; // @[Debug.scala 1147:69:freechips.rocketchip.system.DefaultRV32Config.fir@109995.4]
  assign dmiProgramBufferWrEnMaybe_38 = _T_3694 & _T_2839; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@111204.4]
  assign dmiProgramBufferRdEn_38 = _T_3528 & _T_2837; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@111202.4]
  assign dmiProgramBufferAccessVec_38 = dmiProgramBufferWrEnMaybe_38 | dmiProgramBufferRdEn_38; // @[Debug.scala 1144:108:freechips.rocketchip.system.DefaultRV32Config.fir@109866.4]
  assign _T_204 = _T_203 | dmiProgramBufferAccessVec_38; // @[Debug.scala 1147:69:freechips.rocketchip.system.DefaultRV32Config.fir@109996.4]
  assign dmiProgramBufferWrEnMaybe_39 = _T_3694 & _T_2864; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@111234.4]
  assign dmiProgramBufferRdEn_39 = _T_3528 & _T_2862; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@111232.4]
  assign dmiProgramBufferAccessVec_39 = dmiProgramBufferWrEnMaybe_39 | dmiProgramBufferRdEn_39; // @[Debug.scala 1144:108:freechips.rocketchip.system.DefaultRV32Config.fir@109867.4]
  assign _T_205 = _T_204 | dmiProgramBufferAccessVec_39; // @[Debug.scala 1147:69:freechips.rocketchip.system.DefaultRV32Config.fir@109997.4]
  assign _T_206 = _T_205 | dmiProgramBufferAccessVec_40; // @[Debug.scala 1147:69:freechips.rocketchip.system.DefaultRV32Config.fir@109998.4]
  assign dmiProgramBufferWrEnMaybe_41 = _T_3699 & _T_2814; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@110509.4]
  assign dmiProgramBufferRdEn_41 = _T_3533 & _T_2812; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@110507.4]
  assign dmiProgramBufferAccessVec_41 = dmiProgramBufferWrEnMaybe_41 | dmiProgramBufferRdEn_41; // @[Debug.scala 1144:108:freechips.rocketchip.system.DefaultRV32Config.fir@109869.4]
  assign _T_207 = _T_206 | dmiProgramBufferAccessVec_41; // @[Debug.scala 1147:69:freechips.rocketchip.system.DefaultRV32Config.fir@109999.4]
  assign dmiProgramBufferWrEnMaybe_42 = _T_3699 & _T_2839; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@110539.4]
  assign dmiProgramBufferRdEn_42 = _T_3533 & _T_2837; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@110537.4]
  assign dmiProgramBufferAccessVec_42 = dmiProgramBufferWrEnMaybe_42 | dmiProgramBufferRdEn_42; // @[Debug.scala 1144:108:freechips.rocketchip.system.DefaultRV32Config.fir@109870.4]
  assign _T_208 = _T_207 | dmiProgramBufferAccessVec_42; // @[Debug.scala 1147:69:freechips.rocketchip.system.DefaultRV32Config.fir@110000.4]
  assign dmiProgramBufferWrEnMaybe_43 = _T_3699 & _T_2864; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@110569.4]
  assign dmiProgramBufferRdEn_43 = _T_3533 & _T_2862; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@110567.4]
  assign dmiProgramBufferAccessVec_43 = dmiProgramBufferWrEnMaybe_43 | dmiProgramBufferRdEn_43; // @[Debug.scala 1144:108:freechips.rocketchip.system.DefaultRV32Config.fir@109871.4]
  assign _T_209 = _T_208 | dmiProgramBufferAccessVec_43; // @[Debug.scala 1147:69:freechips.rocketchip.system.DefaultRV32Config.fir@110001.4]
  assign _T_210 = _T_209 | dmiProgramBufferAccessVec_44; // @[Debug.scala 1147:69:freechips.rocketchip.system.DefaultRV32Config.fir@110002.4]
  assign dmiProgramBufferWrEnMaybe_45 = _T_3704 & _T_2814; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@112732.4]
  assign dmiProgramBufferRdEn_45 = _T_3538 & _T_2812; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@112730.4]
  assign dmiProgramBufferAccessVec_45 = dmiProgramBufferWrEnMaybe_45 | dmiProgramBufferRdEn_45; // @[Debug.scala 1144:108:freechips.rocketchip.system.DefaultRV32Config.fir@109873.4]
  assign _T_211 = _T_210 | dmiProgramBufferAccessVec_45; // @[Debug.scala 1147:69:freechips.rocketchip.system.DefaultRV32Config.fir@110003.4]
  assign dmiProgramBufferWrEnMaybe_46 = _T_3704 & _T_2839; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@112762.4]
  assign dmiProgramBufferRdEn_46 = _T_3538 & _T_2837; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@112760.4]
  assign dmiProgramBufferAccessVec_46 = dmiProgramBufferWrEnMaybe_46 | dmiProgramBufferRdEn_46; // @[Debug.scala 1144:108:freechips.rocketchip.system.DefaultRV32Config.fir@109874.4]
  assign _T_212 = _T_211 | dmiProgramBufferAccessVec_46; // @[Debug.scala 1147:69:freechips.rocketchip.system.DefaultRV32Config.fir@110004.4]
  assign dmiProgramBufferWrEnMaybe_47 = _T_3704 & _T_2864; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@112792.4]
  assign dmiProgramBufferRdEn_47 = _T_3538 & _T_2862; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@112790.4]
  assign dmiProgramBufferAccessVec_47 = dmiProgramBufferWrEnMaybe_47 | dmiProgramBufferRdEn_47; // @[Debug.scala 1144:108:freechips.rocketchip.system.DefaultRV32Config.fir@109875.4]
  assign _T_213 = _T_212 | dmiProgramBufferAccessVec_47; // @[Debug.scala 1147:69:freechips.rocketchip.system.DefaultRV32Config.fir@110005.4]
  assign _T_214 = _T_213 | dmiProgramBufferAccessVec_48; // @[Debug.scala 1147:69:freechips.rocketchip.system.DefaultRV32Config.fir@110006.4]
  assign dmiProgramBufferWrEnMaybe_49 = _T_3709 & _T_2814; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@112265.4]
  assign dmiProgramBufferRdEn_49 = _T_3543 & _T_2812; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@112263.4]
  assign dmiProgramBufferAccessVec_49 = dmiProgramBufferWrEnMaybe_49 | dmiProgramBufferRdEn_49; // @[Debug.scala 1144:108:freechips.rocketchip.system.DefaultRV32Config.fir@109877.4]
  assign _T_215 = _T_214 | dmiProgramBufferAccessVec_49; // @[Debug.scala 1147:69:freechips.rocketchip.system.DefaultRV32Config.fir@110007.4]
  assign dmiProgramBufferWrEnMaybe_50 = _T_3709 & _T_2839; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@112295.4]
  assign dmiProgramBufferRdEn_50 = _T_3543 & _T_2837; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@112293.4]
  assign dmiProgramBufferAccessVec_50 = dmiProgramBufferWrEnMaybe_50 | dmiProgramBufferRdEn_50; // @[Debug.scala 1144:108:freechips.rocketchip.system.DefaultRV32Config.fir@109878.4]
  assign _T_216 = _T_215 | dmiProgramBufferAccessVec_50; // @[Debug.scala 1147:69:freechips.rocketchip.system.DefaultRV32Config.fir@110008.4]
  assign dmiProgramBufferWrEnMaybe_51 = _T_3709 & _T_2864; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@112325.4]
  assign dmiProgramBufferRdEn_51 = _T_3543 & _T_2862; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@112323.4]
  assign dmiProgramBufferAccessVec_51 = dmiProgramBufferWrEnMaybe_51 | dmiProgramBufferRdEn_51; // @[Debug.scala 1144:108:freechips.rocketchip.system.DefaultRV32Config.fir@109879.4]
  assign _T_217 = _T_216 | dmiProgramBufferAccessVec_51; // @[Debug.scala 1147:69:freechips.rocketchip.system.DefaultRV32Config.fir@110009.4]
  assign _T_218 = _T_217 | dmiProgramBufferAccessVec_52; // @[Debug.scala 1147:69:freechips.rocketchip.system.DefaultRV32Config.fir@110010.4]
  assign dmiProgramBufferWrEnMaybe_53 = _T_3714 & _T_2814; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@111528.4]
  assign dmiProgramBufferRdEn_53 = _T_3548 & _T_2812; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@111526.4]
  assign dmiProgramBufferAccessVec_53 = dmiProgramBufferWrEnMaybe_53 | dmiProgramBufferRdEn_53; // @[Debug.scala 1144:108:freechips.rocketchip.system.DefaultRV32Config.fir@109881.4]
  assign _T_219 = _T_218 | dmiProgramBufferAccessVec_53; // @[Debug.scala 1147:69:freechips.rocketchip.system.DefaultRV32Config.fir@110011.4]
  assign dmiProgramBufferWrEnMaybe_54 = _T_3714 & _T_2839; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@111558.4]
  assign dmiProgramBufferRdEn_54 = _T_3548 & _T_2837; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@111556.4]
  assign dmiProgramBufferAccessVec_54 = dmiProgramBufferWrEnMaybe_54 | dmiProgramBufferRdEn_54; // @[Debug.scala 1144:108:freechips.rocketchip.system.DefaultRV32Config.fir@109882.4]
  assign _T_220 = _T_219 | dmiProgramBufferAccessVec_54; // @[Debug.scala 1147:69:freechips.rocketchip.system.DefaultRV32Config.fir@110012.4]
  assign dmiProgramBufferWrEnMaybe_55 = _T_3714 & _T_2864; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@111588.4]
  assign dmiProgramBufferRdEn_55 = _T_3548 & _T_2862; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@111586.4]
  assign dmiProgramBufferAccessVec_55 = dmiProgramBufferWrEnMaybe_55 | dmiProgramBufferRdEn_55; // @[Debug.scala 1144:108:freechips.rocketchip.system.DefaultRV32Config.fir@109883.4]
  assign _T_221 = _T_220 | dmiProgramBufferAccessVec_55; // @[Debug.scala 1147:69:freechips.rocketchip.system.DefaultRV32Config.fir@110013.4]
  assign _T_222 = _T_221 | dmiProgramBufferAccessVec_56; // @[Debug.scala 1147:69:freechips.rocketchip.system.DefaultRV32Config.fir@110014.4]
  assign dmiProgramBufferWrEnMaybe_57 = _T_3719 & _T_2814; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@110820.4]
  assign dmiProgramBufferRdEn_57 = _T_3553 & _T_2812; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@110818.4]
  assign dmiProgramBufferAccessVec_57 = dmiProgramBufferWrEnMaybe_57 | dmiProgramBufferRdEn_57; // @[Debug.scala 1144:108:freechips.rocketchip.system.DefaultRV32Config.fir@109885.4]
  assign _T_223 = _T_222 | dmiProgramBufferAccessVec_57; // @[Debug.scala 1147:69:freechips.rocketchip.system.DefaultRV32Config.fir@110015.4]
  assign dmiProgramBufferWrEnMaybe_58 = _T_3719 & _T_2839; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@110850.4]
  assign dmiProgramBufferRdEn_58 = _T_3553 & _T_2837; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@110848.4]
  assign dmiProgramBufferAccessVec_58 = dmiProgramBufferWrEnMaybe_58 | dmiProgramBufferRdEn_58; // @[Debug.scala 1144:108:freechips.rocketchip.system.DefaultRV32Config.fir@109886.4]
  assign _T_224 = _T_223 | dmiProgramBufferAccessVec_58; // @[Debug.scala 1147:69:freechips.rocketchip.system.DefaultRV32Config.fir@110016.4]
  assign dmiProgramBufferWrEnMaybe_59 = _T_3719 & _T_2864; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@110880.4]
  assign dmiProgramBufferRdEn_59 = _T_3553 & _T_2862; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@110878.4]
  assign dmiProgramBufferAccessVec_59 = dmiProgramBufferWrEnMaybe_59 | dmiProgramBufferRdEn_59; // @[Debug.scala 1144:108:freechips.rocketchip.system.DefaultRV32Config.fir@109887.4]
  assign _T_225 = _T_224 | dmiProgramBufferAccessVec_59; // @[Debug.scala 1147:69:freechips.rocketchip.system.DefaultRV32Config.fir@110017.4]
  assign _T_226 = _T_225 | dmiProgramBufferAccessVec_60; // @[Debug.scala 1147:69:freechips.rocketchip.system.DefaultRV32Config.fir@110018.4]
  assign dmiProgramBufferWrEnMaybe_61 = _T_3724 & _T_2814; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@113253.4]
  assign dmiProgramBufferRdEn_61 = _T_3558 & _T_2812; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@113251.4]
  assign dmiProgramBufferAccessVec_61 = dmiProgramBufferWrEnMaybe_61 | dmiProgramBufferRdEn_61; // @[Debug.scala 1144:108:freechips.rocketchip.system.DefaultRV32Config.fir@109889.4]
  assign _T_227 = _T_226 | dmiProgramBufferAccessVec_61; // @[Debug.scala 1147:69:freechips.rocketchip.system.DefaultRV32Config.fir@110019.4]
  assign dmiProgramBufferWrEnMaybe_62 = _T_3724 & _T_2839; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@113283.4]
  assign dmiProgramBufferRdEn_62 = _T_3558 & _T_2837; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@113281.4]
  assign dmiProgramBufferAccessVec_62 = dmiProgramBufferWrEnMaybe_62 | dmiProgramBufferRdEn_62; // @[Debug.scala 1144:108:freechips.rocketchip.system.DefaultRV32Config.fir@109890.4]
  assign _T_228 = _T_227 | dmiProgramBufferAccessVec_62; // @[Debug.scala 1147:69:freechips.rocketchip.system.DefaultRV32Config.fir@110020.4]
  assign dmiProgramBufferWrEnMaybe_63 = _T_3724 & _T_2864; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@113313.4]
  assign dmiProgramBufferRdEn_63 = _T_3558 & _T_2862; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@113311.4]
  assign dmiProgramBufferAccessVec_63 = dmiProgramBufferWrEnMaybe_63 | dmiProgramBufferRdEn_63; // @[Debug.scala 1144:108:freechips.rocketchip.system.DefaultRV32Config.fir@109891.4]
  assign dmiProgramBufferAccess = _T_228 | dmiProgramBufferAccessVec_63; // @[Debug.scala 1147:69:freechips.rocketchip.system.DefaultRV32Config.fir@110021.4]
  assign _T_44800 = dmiProgramBufferAccess & _T_44785; // @[Debug.scala 1580:42:freechips.rocketchip.system.DefaultRV32Config.fir@168687.4]
  assign errorBusy = _T_44798 | _T_44800; // @[Debug.scala 1579:74:freechips.rocketchip.system.DefaultRV32Config.fir@168688.4]
  assign _T_91 = autoexecprogbufWrEnMaybe & ABSTRACTCSWrEnLegal; // @[Debug.scala 1132:38:freechips.rocketchip.system.DefaultRV32Config.fir@109669.6]
  assign ABSTRACTAUTOWrData_autoexecprogbuf = auto_dmi_in_a_bits_data[31:16]; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@110648.4]
  assign _T_93 = autoexecdataWrEnMaybe & ABSTRACTCSWrEnLegal; // @[Debug.scala 1135:35:freechips.rocketchip.system.DefaultRV32Config.fir@109674.6]
  assign ABSTRACTAUTOWrData_autoexecdata = {{11'd0}, auto_dmi_in_a_bits_data[0]}; // @[:freechips.rocketchip.system.DefaultRV32Config.fir@109644.4 :freechips.rocketchip.system.DefaultRV32Config.fir@109645.4 Debug.scala 278:12:freechips.rocketchip.system.DefaultRV32Config.fir@110602.4]
  assign _T_94 = ABSTRACTAUTOWrData_autoexecdata & 12'h1; // @[Debug.scala 1136:73:freechips.rocketchip.system.DefaultRV32Config.fir@109676.8]
  assign COMMANDWrData_control = COMMANDWrDataVal[23:0]; // @[Debug.scala 1163:65:freechips.rocketchip.system.DefaultRV32Config.fir@110150.4]
  assign _T_42528 = _T_42196 & _T_33985[66]; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@162780.4]
  assign _T_42529 = _T_42528 & _T_6089; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@162781.4]
  assign hartResumingWrEn = _T_42529 & _T_25711; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@134493.4]
  assign _GEN_68 = hartResumingWrEn ? 1'h0 : haltedBitRegs_0; // @[Debug.scala 1208:39:freechips.rocketchip.system.DefaultRV32Config.fir@110269.10]
  assign _T_42518 = _T_42196 & _T_33985[64]; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@162764.4]
  assign _T_42519 = _T_42518 & _T_6089; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@162765.4]
  assign hartHaltedWrEn = _T_42519 & _T_25711; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@130810.4]
  assign _GEN_69 = hartHaltedWrEn | _GEN_68; // @[Debug.scala 1204:37:freechips.rocketchip.system.DefaultRV32Config.fir@110262.8]
  assign _GEN_71 = hartIsInResetSync_0 ? 1'h0 : resumeReqRegs_0; // @[Debug.scala 1201:45:freechips.rocketchip.system.DefaultRV32Config.fir@110257.6]
  assign _GEN_73 = hartResumingWrEn ? 1'h0 : _GEN_71; // @[Debug.scala 1218:33:freechips.rocketchip.system.DefaultRV32Config.fir@110275.6]
  assign _GEN_74 = _T_307 | _GEN_73; // @[Debug.scala 1223:52:freechips.rocketchip.system.DefaultRV32Config.fir@110282.6]
  assign _T_564 = {programBufferMem_43,programBufferMem_42,programBufferMem_41,programBufferMem_40}; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@110585.4]
  assign _T_610 = {1'h0,ABSTRACTAUTOReg_autoexecdata[0]}; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@110633.4]
  assign _T_611 = {{14'd0}, _T_610}; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@110634.4]
  assign _T_635 = {ABSTRACTAUTOReg_autoexecprogbuf,_T_611}; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@110660.4]
  assign _T_733 = {programBufferMem_23,programBufferMem_22,programBufferMem_21,programBufferMem_20}; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@110778.4]
  assign _T_831 = {programBufferMem_59,programBufferMem_58,programBufferMem_57,programBufferMem_56}; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@110896.4]
  assign _T_929 = {programBufferMem_27,programBufferMem_26,programBufferMem_25,programBufferMem_24}; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@111014.4]
  assign _T_1027 = {programBufferMem_7,programBufferMem_6,programBufferMem_5,programBufferMem_4}; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@111132.4]
  assign _T_1125 = {programBufferMem_39,programBufferMem_38,programBufferMem_37,programBufferMem_36}; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@111250.4]
  assign _T_1223 = {programBufferMem_3,programBufferMem_2,programBufferMem_1,programBufferMem_0}; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@111368.4]
  assign _T_1321 = {programBufferMem_11,programBufferMem_10,programBufferMem_9,programBufferMem_8}; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@111486.4]
  assign _T_1419 = {programBufferMem_55,programBufferMem_54,programBufferMem_53,programBufferMem_52}; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@111604.4]
  assign _T_1760 = {resumeAcks_0,1'h0,1'h0,1'h0,1'h0,_T_23,_T_23,haltedBitRegs_0,haltedBitRegs_0,8'ha2}; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@111945.4]
  assign _T_1852 = {1'h0,haveResetBitRegs_0,haveResetBitRegs_0,resumeAcks_0,_T_1760}; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@112037.4]
  assign _T_1853 = {{1'd0}, _T_1852}; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@112038.4]
  assign _T_1875 = {1'h0,_T_1853}; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@112060.4]
  assign abstractCommandBusy = ctrlStateReg != 2'h0; // @[Debug.scala 1567:42:freechips.rocketchip.system.DefaultRV32Config.fir@168660.4]
  assign _T_2013 = {1'h0,abstractCommandBusy,1'h0,ABSTRACTCSReg_cmderr,8'h1}; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@112200.4]
  assign _T_2014 = {{10'd0}, _T_2013}; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@112201.4]
  assign _T_2036 = {5'h10,_T_2014}; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@112223.4]
  assign _T_2134 = {programBufferMem_51,programBufferMem_50,programBufferMem_49,programBufferMem_48}; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@112341.4]
  assign _T_2232 = {programBufferMem_31,programBufferMem_30,programBufferMem_29,programBufferMem_28}; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@112459.4]
  assign _T_2330 = {programBufferMem_15,programBufferMem_14,programBufferMem_13,programBufferMem_12}; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@112577.4]
  assign _T_2541 = {programBufferMem_47,programBufferMem_46,programBufferMem_45,programBufferMem_44}; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@112808.4]
  assign _T_2639 = {programBufferMem_35,programBufferMem_34,programBufferMem_33,programBufferMem_32}; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@112926.4]
  assign _T_2760 = {programBufferMem_19,programBufferMem_18,programBufferMem_17,programBufferMem_16}; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@113072.4]
  assign _T_2879 = {abstractDataMem_3,abstractDataMem_2,abstractDataMem_1,abstractDataMem_0}; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@113211.4]
  assign _T_2977 = {programBufferMem_63,programBufferMem_62,programBufferMem_61,programBufferMem_60}; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@113329.4]
  assign _GEN_275 = 5'h1 == _T_2990 ? _T_389 : _T_407; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@114936.4]
  assign _GEN_276 = 5'h2 == _T_2990 ? _T_389 : _GEN_275; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@114936.4]
  assign _GEN_277 = 5'h3 == _T_2990 ? _T_389 : _GEN_276; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@114936.4]
  assign _GEN_278 = 5'h4 == _T_2990 ? _T_433 : _GEN_277; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@114936.4]
  assign _GEN_3664 = 5'h5 == _T_2990; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@114936.4]
  assign _GEN_279 = _GEN_3664 | _GEN_278; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@114936.4]
  assign _GEN_280 = 5'h6 == _T_2990 ? _T_389 : _GEN_279; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@114936.4]
  assign _GEN_281 = 5'h7 == _T_2990 ? _T_389 : _GEN_280; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@114936.4]
  assign _GEN_282 = 5'h8 == _T_2990 ? _T_389 : _GEN_281; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@114936.4]
  assign _GEN_3665 = 5'h9 == _T_2990; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@114936.4]
  assign _GEN_283 = _GEN_3665 | _GEN_282; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@114936.4]
  assign _GEN_3666 = 5'ha == _T_2990; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@114936.4]
  assign _GEN_284 = _GEN_3666 | _GEN_283; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@114936.4]
  assign _GEN_3667 = 5'hb == _T_2990; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@114936.4]
  assign _GEN_285 = _GEN_3667 | _GEN_284; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@114936.4]
  assign _GEN_3668 = 5'hc == _T_2990; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@114936.4]
  assign _GEN_286 = _GEN_3668 | _GEN_285; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@114936.4]
  assign _GEN_3669 = 5'hd == _T_2990; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@114936.4]
  assign _GEN_287 = _GEN_3669 | _GEN_286; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@114936.4]
  assign _GEN_3670 = 5'he == _T_2990; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@114936.4]
  assign _GEN_288 = _GEN_3670 | _GEN_287; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@114936.4]
  assign _GEN_3671 = 5'hf == _T_2990; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@114936.4]
  assign _GEN_289 = _GEN_3671 | _GEN_288; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@114936.4]
  assign _GEN_290 = 5'h10 == _T_2990 ? _T_433 : _GEN_289; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@114936.4]
  assign _GEN_291 = 5'h11 == _T_2990 ? _T_433 : _GEN_290; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@114936.4]
  assign _GEN_292 = 5'h12 == _T_2990 ? _T_433 : _GEN_291; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@114936.4]
  assign _GEN_293 = 5'h13 == _T_2990 ? _T_433 : _GEN_292; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@114936.4]
  assign _GEN_294 = 5'h14 == _T_2990 ? _T_433 : _GEN_293; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@114936.4]
  assign _GEN_295 = 5'h15 == _T_2990 ? _T_433 : _GEN_294; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@114936.4]
  assign _GEN_296 = 5'h16 == _T_2990 ? _T_433 : _GEN_295; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@114936.4]
  assign _GEN_297 = 5'h17 == _T_2990 ? _T_433 : _GEN_296; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@114936.4]
  assign _GEN_298 = 5'h18 == _T_2990 ? _T_433 : _GEN_297; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@114936.4]
  assign _GEN_299 = 5'h19 == _T_2990 ? _T_433 : _GEN_298; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@114936.4]
  assign _GEN_300 = 5'h1a == _T_2990 ? _T_433 : _GEN_299; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@114936.4]
  assign _GEN_301 = 5'h1b == _T_2990 ? _T_433 : _GEN_300; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@114936.4]
  assign _GEN_302 = 5'h1c == _T_2990 ? _T_433 : _GEN_301; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@114936.4]
  assign _GEN_303 = 5'h1d == _T_2990 ? _T_433 : _GEN_302; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@114936.4]
  assign _GEN_304 = 5'h1e == _T_2990 ? _T_433 : _GEN_303; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@114936.4]
  assign _GEN_305 = 5'h1f == _T_2990 ? _T_433 : _GEN_304; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@114936.4]
  assign _T_3740_1 = {{9'd0}, _T_1875}; // @[MuxLiteral.scala 48:48:freechips.rocketchip.system.DefaultRV32Config.fir@114938.4 MuxLiteral.scala 48:48:freechips.rocketchip.system.DefaultRV32Config.fir@114941.4]
  assign _GEN_307 = 5'h1 == _T_2990 ? _T_3740_1 : haltedStatus_0; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@114972.4]
  assign _GEN_308 = 5'h2 == _T_2990 ? 32'h111380 : _GEN_307; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@114972.4]
  assign _GEN_309 = 5'h3 == _T_2990 ? HALTSUM1RdData_haltsum1 : _GEN_308; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@114972.4]
  assign _GEN_310 = 5'h4 == _T_2990 ? _T_2879 : _GEN_309; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@114972.4]
  assign _GEN_311 = 5'h5 == _T_2990 ? 32'h0 : _GEN_310; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@114972.4]
  assign _T_3740_6 = {{3'd0}, _T_2036}; // @[MuxLiteral.scala 48:48:freechips.rocketchip.system.DefaultRV32Config.fir@114938.4 MuxLiteral.scala 48:48:freechips.rocketchip.system.DefaultRV32Config.fir@114946.4]
  assign _GEN_312 = 5'h6 == _T_2990 ? _T_3740_6 : _GEN_311; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@114972.4]
  assign _GEN_313 = 5'h7 == _T_2990 ? _T_3960 : _GEN_312; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@114972.4]
  assign _GEN_314 = 5'h8 == _T_2990 ? _T_635 : _GEN_313; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@114972.4]
  assign _GEN_315 = 5'h9 == _T_2990 ? 32'h0 : _GEN_314; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@114972.4]
  assign _GEN_316 = 5'ha == _T_2990 ? 32'h0 : _GEN_315; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@114972.4]
  assign _GEN_317 = 5'hb == _T_2990 ? 32'h0 : _GEN_316; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@114972.4]
  assign _GEN_318 = 5'hc == _T_2990 ? 32'h0 : _GEN_317; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@114972.4]
  assign _GEN_319 = 5'hd == _T_2990 ? 32'h0 : _GEN_318; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@114972.4]
  assign _GEN_320 = 5'he == _T_2990 ? 32'h0 : _GEN_319; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@114972.4]
  assign _GEN_321 = 5'hf == _T_2990 ? 32'h0 : _GEN_320; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@114972.4]
  assign _GEN_322 = 5'h10 == _T_2990 ? _T_1223 : _GEN_321; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@114972.4]
  assign _GEN_323 = 5'h11 == _T_2990 ? _T_1027 : _GEN_322; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@114972.4]
  assign _GEN_324 = 5'h12 == _T_2990 ? _T_1321 : _GEN_323; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@114972.4]
  assign _GEN_325 = 5'h13 == _T_2990 ? _T_2330 : _GEN_324; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@114972.4]
  assign _GEN_326 = 5'h14 == _T_2990 ? _T_2760 : _GEN_325; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@114972.4]
  assign _GEN_327 = 5'h15 == _T_2990 ? _T_733 : _GEN_326; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@114972.4]
  assign _GEN_328 = 5'h16 == _T_2990 ? _T_929 : _GEN_327; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@114972.4]
  assign _GEN_329 = 5'h17 == _T_2990 ? _T_2232 : _GEN_328; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@114972.4]
  assign _GEN_330 = 5'h18 == _T_2990 ? _T_2639 : _GEN_329; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@114972.4]
  assign _GEN_331 = 5'h19 == _T_2990 ? _T_1125 : _GEN_330; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@114972.4]
  assign _GEN_332 = 5'h1a == _T_2990 ? _T_564 : _GEN_331; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@114972.4]
  assign _GEN_333 = 5'h1b == _T_2990 ? _T_2541 : _GEN_332; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@114972.4]
  assign _GEN_334 = 5'h1c == _T_2990 ? _T_2134 : _GEN_333; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@114972.4]
  assign _GEN_335 = 5'h1d == _T_2990 ? _T_1419 : _GEN_334; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@114972.4]
  assign _GEN_336 = 5'h1e == _T_2990 ? _T_831 : _GEN_335; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@114972.4]
  assign _GEN_337 = 5'h1f == _T_2990 ? _T_2977 : _GEN_336; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@114972.4]
  assign _T_3749 = dmiAbstractDataWrEnMaybe_0 & ABSTRACTCSWrEnLegal; // @[Debug.scala 1346:60:freechips.rocketchip.system.DefaultRV32Config.fir@115004.4]
  assign _T_3751 = dmiAbstractDataWrEnMaybe_1 & ABSTRACTCSWrEnLegal; // @[Debug.scala 1346:60:freechips.rocketchip.system.DefaultRV32Config.fir@115009.4]
  assign _T_3753 = dmiAbstractDataWrEnMaybe_2 & ABSTRACTCSWrEnLegal; // @[Debug.scala 1346:60:freechips.rocketchip.system.DefaultRV32Config.fir@115014.4]
  assign _T_3755 = dmiAbstractDataWrEnMaybe_3 & ABSTRACTCSWrEnLegal; // @[Debug.scala 1346:60:freechips.rocketchip.system.DefaultRV32Config.fir@115019.4]
  assign _T_3757 = dmiProgramBufferWrEnMaybe_0 & ABSTRACTCSWrEnLegal; // @[Debug.scala 1368:61:freechips.rocketchip.system.DefaultRV32Config.fir@115024.4]
  assign _T_3759 = dmiProgramBufferWrEnMaybe_1 & ABSTRACTCSWrEnLegal; // @[Debug.scala 1368:61:freechips.rocketchip.system.DefaultRV32Config.fir@115029.4]
  assign _T_3761 = dmiProgramBufferWrEnMaybe_2 & ABSTRACTCSWrEnLegal; // @[Debug.scala 1368:61:freechips.rocketchip.system.DefaultRV32Config.fir@115034.4]
  assign _T_3763 = dmiProgramBufferWrEnMaybe_3 & ABSTRACTCSWrEnLegal; // @[Debug.scala 1368:61:freechips.rocketchip.system.DefaultRV32Config.fir@115039.4]
  assign _T_3765 = dmiProgramBufferWrEnMaybe_4 & ABSTRACTCSWrEnLegal; // @[Debug.scala 1368:61:freechips.rocketchip.system.DefaultRV32Config.fir@115044.4]
  assign _T_3767 = dmiProgramBufferWrEnMaybe_5 & ABSTRACTCSWrEnLegal; // @[Debug.scala 1368:61:freechips.rocketchip.system.DefaultRV32Config.fir@115049.4]
  assign _T_3769 = dmiProgramBufferWrEnMaybe_6 & ABSTRACTCSWrEnLegal; // @[Debug.scala 1368:61:freechips.rocketchip.system.DefaultRV32Config.fir@115054.4]
  assign _T_3771 = dmiProgramBufferWrEnMaybe_7 & ABSTRACTCSWrEnLegal; // @[Debug.scala 1368:61:freechips.rocketchip.system.DefaultRV32Config.fir@115059.4]
  assign _T_3773 = dmiProgramBufferWrEnMaybe_8 & ABSTRACTCSWrEnLegal; // @[Debug.scala 1368:61:freechips.rocketchip.system.DefaultRV32Config.fir@115064.4]
  assign _T_3775 = dmiProgramBufferWrEnMaybe_9 & ABSTRACTCSWrEnLegal; // @[Debug.scala 1368:61:freechips.rocketchip.system.DefaultRV32Config.fir@115069.4]
  assign _T_3777 = dmiProgramBufferWrEnMaybe_10 & ABSTRACTCSWrEnLegal; // @[Debug.scala 1368:61:freechips.rocketchip.system.DefaultRV32Config.fir@115074.4]
  assign _T_3779 = dmiProgramBufferWrEnMaybe_11 & ABSTRACTCSWrEnLegal; // @[Debug.scala 1368:61:freechips.rocketchip.system.DefaultRV32Config.fir@115079.4]
  assign _T_3781 = dmiProgramBufferWrEnMaybe_12 & ABSTRACTCSWrEnLegal; // @[Debug.scala 1368:61:freechips.rocketchip.system.DefaultRV32Config.fir@115084.4]
  assign _T_3783 = dmiProgramBufferWrEnMaybe_13 & ABSTRACTCSWrEnLegal; // @[Debug.scala 1368:61:freechips.rocketchip.system.DefaultRV32Config.fir@115089.4]
  assign _T_3785 = dmiProgramBufferWrEnMaybe_14 & ABSTRACTCSWrEnLegal; // @[Debug.scala 1368:61:freechips.rocketchip.system.DefaultRV32Config.fir@115094.4]
  assign _T_3787 = dmiProgramBufferWrEnMaybe_15 & ABSTRACTCSWrEnLegal; // @[Debug.scala 1368:61:freechips.rocketchip.system.DefaultRV32Config.fir@115099.4]
  assign _T_3789 = dmiProgramBufferWrEnMaybe_16 & ABSTRACTCSWrEnLegal; // @[Debug.scala 1368:61:freechips.rocketchip.system.DefaultRV32Config.fir@115104.4]
  assign _T_3791 = dmiProgramBufferWrEnMaybe_17 & ABSTRACTCSWrEnLegal; // @[Debug.scala 1368:61:freechips.rocketchip.system.DefaultRV32Config.fir@115109.4]
  assign _T_3793 = dmiProgramBufferWrEnMaybe_18 & ABSTRACTCSWrEnLegal; // @[Debug.scala 1368:61:freechips.rocketchip.system.DefaultRV32Config.fir@115114.4]
  assign _T_3795 = dmiProgramBufferWrEnMaybe_19 & ABSTRACTCSWrEnLegal; // @[Debug.scala 1368:61:freechips.rocketchip.system.DefaultRV32Config.fir@115119.4]
  assign _T_3797 = dmiProgramBufferWrEnMaybe_20 & ABSTRACTCSWrEnLegal; // @[Debug.scala 1368:61:freechips.rocketchip.system.DefaultRV32Config.fir@115124.4]
  assign _T_3799 = dmiProgramBufferWrEnMaybe_21 & ABSTRACTCSWrEnLegal; // @[Debug.scala 1368:61:freechips.rocketchip.system.DefaultRV32Config.fir@115129.4]
  assign _T_3801 = dmiProgramBufferWrEnMaybe_22 & ABSTRACTCSWrEnLegal; // @[Debug.scala 1368:61:freechips.rocketchip.system.DefaultRV32Config.fir@115134.4]
  assign _T_3803 = dmiProgramBufferWrEnMaybe_23 & ABSTRACTCSWrEnLegal; // @[Debug.scala 1368:61:freechips.rocketchip.system.DefaultRV32Config.fir@115139.4]
  assign _T_3805 = dmiProgramBufferWrEnMaybe_24 & ABSTRACTCSWrEnLegal; // @[Debug.scala 1368:61:freechips.rocketchip.system.DefaultRV32Config.fir@115144.4]
  assign _T_3807 = dmiProgramBufferWrEnMaybe_25 & ABSTRACTCSWrEnLegal; // @[Debug.scala 1368:61:freechips.rocketchip.system.DefaultRV32Config.fir@115149.4]
  assign _T_3809 = dmiProgramBufferWrEnMaybe_26 & ABSTRACTCSWrEnLegal; // @[Debug.scala 1368:61:freechips.rocketchip.system.DefaultRV32Config.fir@115154.4]
  assign _T_3811 = dmiProgramBufferWrEnMaybe_27 & ABSTRACTCSWrEnLegal; // @[Debug.scala 1368:61:freechips.rocketchip.system.DefaultRV32Config.fir@115159.4]
  assign _T_3813 = dmiProgramBufferWrEnMaybe_28 & ABSTRACTCSWrEnLegal; // @[Debug.scala 1368:61:freechips.rocketchip.system.DefaultRV32Config.fir@115164.4]
  assign _T_3815 = dmiProgramBufferWrEnMaybe_29 & ABSTRACTCSWrEnLegal; // @[Debug.scala 1368:61:freechips.rocketchip.system.DefaultRV32Config.fir@115169.4]
  assign _T_3817 = dmiProgramBufferWrEnMaybe_30 & ABSTRACTCSWrEnLegal; // @[Debug.scala 1368:61:freechips.rocketchip.system.DefaultRV32Config.fir@115174.4]
  assign _T_3819 = dmiProgramBufferWrEnMaybe_31 & ABSTRACTCSWrEnLegal; // @[Debug.scala 1368:61:freechips.rocketchip.system.DefaultRV32Config.fir@115179.4]
  assign _T_3821 = dmiProgramBufferWrEnMaybe_32 & ABSTRACTCSWrEnLegal; // @[Debug.scala 1368:61:freechips.rocketchip.system.DefaultRV32Config.fir@115184.4]
  assign _T_3823 = dmiProgramBufferWrEnMaybe_33 & ABSTRACTCSWrEnLegal; // @[Debug.scala 1368:61:freechips.rocketchip.system.DefaultRV32Config.fir@115189.4]
  assign _T_3825 = dmiProgramBufferWrEnMaybe_34 & ABSTRACTCSWrEnLegal; // @[Debug.scala 1368:61:freechips.rocketchip.system.DefaultRV32Config.fir@115194.4]
  assign _T_3827 = dmiProgramBufferWrEnMaybe_35 & ABSTRACTCSWrEnLegal; // @[Debug.scala 1368:61:freechips.rocketchip.system.DefaultRV32Config.fir@115199.4]
  assign _T_3829 = dmiProgramBufferWrEnMaybe_36 & ABSTRACTCSWrEnLegal; // @[Debug.scala 1368:61:freechips.rocketchip.system.DefaultRV32Config.fir@115204.4]
  assign _T_3831 = dmiProgramBufferWrEnMaybe_37 & ABSTRACTCSWrEnLegal; // @[Debug.scala 1368:61:freechips.rocketchip.system.DefaultRV32Config.fir@115209.4]
  assign _T_3833 = dmiProgramBufferWrEnMaybe_38 & ABSTRACTCSWrEnLegal; // @[Debug.scala 1368:61:freechips.rocketchip.system.DefaultRV32Config.fir@115214.4]
  assign _T_3835 = dmiProgramBufferWrEnMaybe_39 & ABSTRACTCSWrEnLegal; // @[Debug.scala 1368:61:freechips.rocketchip.system.DefaultRV32Config.fir@115219.4]
  assign _T_3837 = dmiProgramBufferWrEnMaybe_40 & ABSTRACTCSWrEnLegal; // @[Debug.scala 1368:61:freechips.rocketchip.system.DefaultRV32Config.fir@115224.4]
  assign _T_3839 = dmiProgramBufferWrEnMaybe_41 & ABSTRACTCSWrEnLegal; // @[Debug.scala 1368:61:freechips.rocketchip.system.DefaultRV32Config.fir@115229.4]
  assign _T_3841 = dmiProgramBufferWrEnMaybe_42 & ABSTRACTCSWrEnLegal; // @[Debug.scala 1368:61:freechips.rocketchip.system.DefaultRV32Config.fir@115234.4]
  assign _T_3843 = dmiProgramBufferWrEnMaybe_43 & ABSTRACTCSWrEnLegal; // @[Debug.scala 1368:61:freechips.rocketchip.system.DefaultRV32Config.fir@115239.4]
  assign _T_3845 = dmiProgramBufferWrEnMaybe_44 & ABSTRACTCSWrEnLegal; // @[Debug.scala 1368:61:freechips.rocketchip.system.DefaultRV32Config.fir@115244.4]
  assign _T_3847 = dmiProgramBufferWrEnMaybe_45 & ABSTRACTCSWrEnLegal; // @[Debug.scala 1368:61:freechips.rocketchip.system.DefaultRV32Config.fir@115249.4]
  assign _T_3849 = dmiProgramBufferWrEnMaybe_46 & ABSTRACTCSWrEnLegal; // @[Debug.scala 1368:61:freechips.rocketchip.system.DefaultRV32Config.fir@115254.4]
  assign _T_3851 = dmiProgramBufferWrEnMaybe_47 & ABSTRACTCSWrEnLegal; // @[Debug.scala 1368:61:freechips.rocketchip.system.DefaultRV32Config.fir@115259.4]
  assign _T_3853 = dmiProgramBufferWrEnMaybe_48 & ABSTRACTCSWrEnLegal; // @[Debug.scala 1368:61:freechips.rocketchip.system.DefaultRV32Config.fir@115264.4]
  assign _T_3855 = dmiProgramBufferWrEnMaybe_49 & ABSTRACTCSWrEnLegal; // @[Debug.scala 1368:61:freechips.rocketchip.system.DefaultRV32Config.fir@115269.4]
  assign _T_3857 = dmiProgramBufferWrEnMaybe_50 & ABSTRACTCSWrEnLegal; // @[Debug.scala 1368:61:freechips.rocketchip.system.DefaultRV32Config.fir@115274.4]
  assign _T_3859 = dmiProgramBufferWrEnMaybe_51 & ABSTRACTCSWrEnLegal; // @[Debug.scala 1368:61:freechips.rocketchip.system.DefaultRV32Config.fir@115279.4]
  assign _T_3861 = dmiProgramBufferWrEnMaybe_52 & ABSTRACTCSWrEnLegal; // @[Debug.scala 1368:61:freechips.rocketchip.system.DefaultRV32Config.fir@115284.4]
  assign _T_3863 = dmiProgramBufferWrEnMaybe_53 & ABSTRACTCSWrEnLegal; // @[Debug.scala 1368:61:freechips.rocketchip.system.DefaultRV32Config.fir@115289.4]
  assign _T_3865 = dmiProgramBufferWrEnMaybe_54 & ABSTRACTCSWrEnLegal; // @[Debug.scala 1368:61:freechips.rocketchip.system.DefaultRV32Config.fir@115294.4]
  assign _T_3867 = dmiProgramBufferWrEnMaybe_55 & ABSTRACTCSWrEnLegal; // @[Debug.scala 1368:61:freechips.rocketchip.system.DefaultRV32Config.fir@115299.4]
  assign _T_3869 = dmiProgramBufferWrEnMaybe_56 & ABSTRACTCSWrEnLegal; // @[Debug.scala 1368:61:freechips.rocketchip.system.DefaultRV32Config.fir@115304.4]
  assign _T_3871 = dmiProgramBufferWrEnMaybe_57 & ABSTRACTCSWrEnLegal; // @[Debug.scala 1368:61:freechips.rocketchip.system.DefaultRV32Config.fir@115309.4]
  assign _T_3873 = dmiProgramBufferWrEnMaybe_58 & ABSTRACTCSWrEnLegal; // @[Debug.scala 1368:61:freechips.rocketchip.system.DefaultRV32Config.fir@115314.4]
  assign _T_3875 = dmiProgramBufferWrEnMaybe_59 & ABSTRACTCSWrEnLegal; // @[Debug.scala 1368:61:freechips.rocketchip.system.DefaultRV32Config.fir@115319.4]
  assign _T_3877 = dmiProgramBufferWrEnMaybe_60 & ABSTRACTCSWrEnLegal; // @[Debug.scala 1368:61:freechips.rocketchip.system.DefaultRV32Config.fir@115324.4]
  assign _T_3879 = dmiProgramBufferWrEnMaybe_61 & ABSTRACTCSWrEnLegal; // @[Debug.scala 1368:61:freechips.rocketchip.system.DefaultRV32Config.fir@115329.4]
  assign _T_3881 = dmiProgramBufferWrEnMaybe_62 & ABSTRACTCSWrEnLegal; // @[Debug.scala 1368:61:freechips.rocketchip.system.DefaultRV32Config.fir@115334.4]
  assign _T_3883 = dmiProgramBufferWrEnMaybe_63 & ABSTRACTCSWrEnLegal; // @[Debug.scala 1368:61:freechips.rocketchip.system.DefaultRV32Config.fir@115339.4]
  assign hartGoingId = auto_tl_in_a_bits_data[9:0]; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@126788.4]
  assign _T_3935 = hartGoingId == 10'h0; // @[Debug.scala 1389:28:freechips.rocketchip.system.DefaultRV32Config.fir@115468.10]
  assign _T_3937 = _T_3935 | reset; // @[Debug.scala 1389:15:freechips.rocketchip.system.DefaultRV32Config.fir@115470.10]
  assign _T_3938 = ~_T_3937; // @[Debug.scala 1389:15:freechips.rocketchip.system.DefaultRV32Config.fir@115471.10]
  assign _T_42523 = _T_42196 & _T_33985[65]; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@162772.4]
  assign _T_42524 = _T_42523 & _T_6089; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@162773.4]
  assign hartGoingWrEn = _T_42524 & _T_25711; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@126787.4]
  assign _GEN_406 = hartGoingWrEn ? 1'h0 : goReg; // @[Debug.scala 1388:33:freechips.rocketchip.system.DefaultRV32Config.fir@115467.8]
  assign _GEN_3637 = commandRegBadHaltResume ? 1'h0 : 1'h1; // @[Debug.scala 1633:43:freechips.rocketchip.system.DefaultRV32Config.fir@168747.10]
  assign _GEN_3641 = commandRegIsUnsupported ? 1'h0 : _GEN_3637; // @[Debug.scala 1630:38:freechips.rocketchip.system.DefaultRV32Config.fir@168742.8]
  assign _GEN_3654 = _T_44818 & _GEN_3641; // @[Debug.scala 1623:59:freechips.rocketchip.system.DefaultRV32Config.fir@168741.6]
  assign goAbstract = ABSTRACTCSWrEnLegal ? 1'h0 : _GEN_3654; // @[Debug.scala 1615:47:freechips.rocketchip.system.DefaultRV32Config.fir@168724.4]
  assign _GEN_407 = goAbstract | _GEN_406; // @[Debug.scala 1386:25:freechips.rocketchip.system.DefaultRV32Config.fir@115463.6]
  assign accessRegisterCommandReg_postexec = _T_3960[18]; // @[Debug.scala 1415:73:freechips.rocketchip.system.DefaultRV32Config.fir@115554.4]
  assign accessRegisterCommandReg_size = _T_3960[22:20]; // @[Debug.scala 1415:73:freechips.rocketchip.system.DefaultRV32Config.fir@115558.4]
  assign _T_3972 = accessRegisterCommandReg_regno & 16'h1f; // @[Debug.scala 1464:66:freechips.rocketchip.system.DefaultRV32Config.fir@115584.4]
  assign abstractGeneratedI_rd = _T_3972[4:0]; // @[Debug.scala 1459:34:freechips.rocketchip.system.DefaultRV32Config.fir@115574.4 Debug.scala 1464:31:freechips.rocketchip.system.DefaultRV32Config.fir@115585.4]
  assign _T_3979 = {17'h7000,accessRegisterCommandReg_size,abstractGeneratedI_rd,7'h3}; // @[Debug.scala 1485:36:freechips.rocketchip.system.DefaultRV32Config.fir@115621.6]
  assign _T_3984 = {7'h1c,abstractGeneratedI_rd,5'h0,accessRegisterCommandReg_size,5'h0,7'h23}; // @[Debug.scala 1487:36:freechips.rocketchip.system.DefaultRV32Config.fir@115626.6]
  assign _T_6696 = &_T_6692[7:0]; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@118357.4]
  assign _T_6717 = &_T_6692[15:8]; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@118378.4]
  assign _T_6740 = &_T_6692[23:16]; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@118401.4]
  assign _T_6757 = {6'h0,resumeReqRegs_0,goReg,6'h0,resumeReqRegs_0,goReg,6'h0,resumeReqRegs_0,goReg}; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@118418.4]
  assign _T_6763 = &_T_6692[31:24]; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@118424.4]
  assign _T_6780 = {6'h0,resumeReqRegs_0,goReg,_T_6757}; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@118441.4]
  assign _T_38152 = _T_42196 & _T_33985[217]; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@153307.4]
  assign _T_38153 = _T_38152 & _T_6089; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@153308.4]
  assign _T_7603 = _T_38153 & _T_6696; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@119264.4]
  assign _T_7626 = _T_38153 & _T_6717; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@119290.4]
  assign _T_7651 = _T_38153 & _T_6740; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@119318.4]
  assign _T_7676 = _T_38153 & _T_6763; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@119346.4]
  assign _T_38147 = _T_42196 & _T_33985[216]; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@153296.4]
  assign _T_38148 = _T_38147 & _T_6089; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@153297.4]
  assign _T_10671 = _T_38148 & _T_6696; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@122344.4]
  assign _T_10694 = _T_38148 & _T_6717; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@122370.4]
  assign _T_10719 = _T_38148 & _T_6740; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@122398.4]
  assign _T_10744 = _T_38148 & _T_6763; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@122426.4]
  assign _T_38122 = _T_42196 & _T_33985[211]; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@153241.4]
  assign _T_38123 = _T_38122 & _T_6089; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@153242.4]
  assign _T_11219 = _T_38123 & _T_6696; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@122904.4]
  assign _T_11242 = _T_38123 & _T_6717; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@122930.4]
  assign _T_11267 = _T_38123 & _T_6740; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@122958.4]
  assign _T_11292 = _T_38123 & _T_6763; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@122986.4]
  assign _T_38172 = _T_42196 & _T_33985[221]; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@153351.4]
  assign _T_38173 = _T_38172 & _T_6089; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@153352.4]
  assign _T_11947 = _T_38173 & _T_6696; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@123644.4]
  assign _T_11970 = _T_38173 & _T_6717; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@123670.4]
  assign _T_11995 = _T_38173 & _T_6740; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@123698.4]
  assign _T_12020 = _T_38173 & _T_6763; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@123726.4]
  assign _T_38167 = _T_42196 & _T_33985[220]; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@153340.4]
  assign _T_38168 = _T_38167 & _T_6089; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@153341.4]
  assign _T_13686 = _T_38168 & _T_6696; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@125395.4]
  assign _T_13709 = _T_38168 & _T_6717; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@125421.4]
  assign _T_13734 = _T_38168 & _T_6740; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@125449.4]
  assign _T_13759 = _T_38168 & _T_6763; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@125477.4]
  assign _T_38187 = _T_42196 & _T_33985[224]; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@153384.4]
  assign _T_38188 = _T_38187 & _T_6089; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@153385.4]
  assign _T_15806 = _T_38188 & _T_6696; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@127529.4]
  assign _T_15829 = _T_38188 & _T_6717; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@127555.4]
  assign _T_15854 = _T_38188 & _T_6740; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@127583.4]
  assign _T_15879 = _T_38188 & _T_6763; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@127611.4]
  assign _T_38127 = _T_42196 & _T_33985[212]; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@153252.4]
  assign _T_38128 = _T_38127 & _T_6089; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@153253.4]
  assign _T_17254 = _T_38128 & _T_6696; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@128989.4]
  assign _T_17277 = _T_38128 & _T_6717; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@129015.4]
  assign _T_17302 = _T_38128 & _T_6740; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@129043.4]
  assign _T_17327 = _T_38128 & _T_6763; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@129071.4]
  assign _T_38162 = _T_42196 & _T_33985[219]; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@153329.4]
  assign _T_38163 = _T_38162 & _T_6089; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@153330.4]
  assign _T_20793 = _T_38163 & _T_6696; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@132542.4]
  assign _T_20816 = _T_38163 & _T_6717; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@132568.4]
  assign _T_20841 = _T_38163 & _T_6740; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@132596.4]
  assign _T_20866 = _T_38163 & _T_6763; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@132624.4]
  assign _T_38107 = _T_42196 & _T_33985[208]; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@153208.4]
  assign _T_38108 = _T_38107 & _T_6089; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@153209.4]
  assign _T_21791 = _T_38108 & _T_6696; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@133552.4]
  assign _T_21814 = _T_38108 & _T_6717; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@133578.4]
  assign _T_21839 = _T_38108 & _T_6740; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@133606.4]
  assign _T_21864 = _T_38108 & _T_6763; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@133634.4]
  assign _T_38132 = _T_42196 & _T_33985[213]; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@153263.4]
  assign _T_38133 = _T_38132 & _T_6089; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@153264.4]
  assign _T_22429 = _T_38133 & _T_6696; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@134202.4]
  assign _T_22452 = _T_38133 & _T_6717; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@134228.4]
  assign _T_22477 = _T_38133 & _T_6740; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@134256.4]
  assign _T_22502 = _T_38133 & _T_6763; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@134284.4]
  assign _T_38182 = _T_42196 & _T_33985[223]; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@153373.4]
  assign _T_38183 = _T_38182 & _T_6089; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@153374.4]
  assign _T_23268 = _T_38183 & _T_6696; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@135055.4]
  assign _T_23291 = _T_38183 & _T_6717; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@135081.4]
  assign _T_23316 = _T_38183 & _T_6740; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@135109.4]
  assign _T_23341 = _T_38183 & _T_6763; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@135137.4]
  assign _T_38112 = _T_42196 & _T_33985[209]; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@153219.4]
  assign _T_38113 = _T_38112 & _T_6089; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@153220.4]
  assign _T_24446 = _T_38113 & _T_6696; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@136245.4]
  assign _T_24469 = _T_38113 & _T_6717; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@136271.4]
  assign _T_24494 = _T_38113 & _T_6740; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@136299.4]
  assign _T_24519 = _T_38113 & _T_6763; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@136327.4]
  assign _T_38157 = _T_42196 & _T_33985[218]; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@153318.4]
  assign _T_38158 = _T_38157 & _T_6089; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@153319.4]
  assign _T_27445 = _T_38158 & _T_6696; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@139258.4]
  assign _T_27468 = _T_38158 & _T_6717; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@139284.4]
  assign _T_27493 = _T_38158 & _T_6740; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@139312.4]
  assign _T_27518 = _T_38158 & _T_6763; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@139340.4]
  assign _T_38137 = _T_42196 & _T_33985[214]; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@153274.4]
  assign _T_38138 = _T_38137 & _T_6089; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@153275.4]
  assign _T_29094 = _T_38138 & _T_6696; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@140919.4]
  assign _T_29117 = _T_38138 & _T_6717; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@140945.4]
  assign _T_29142 = _T_38138 & _T_6740; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@140973.4]
  assign _T_29167 = _T_38138 & _T_6763; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@141001.4]
  assign _T_38117 = _T_42196 & _T_33985[210]; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@153230.4]
  assign _T_38118 = _T_38117 & _T_6089; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@153231.4]
  assign _T_30272 = _T_38118 & _T_6696; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@142109.4]
  assign _T_30295 = _T_38118 & _T_6717; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@142135.4]
  assign _T_30320 = _T_38118 & _T_6740; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@142163.4]
  assign _T_30345 = _T_38118 & _T_6763; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@142191.4]
  assign _T_38142 = _T_42196 & _T_33985[215]; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@153285.4]
  assign _T_38143 = _T_38142 & _T_6089; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@153286.4]
  assign _T_32890 = _T_38143 & _T_6696; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@144739.4]
  assign _T_32913 = _T_38143 & _T_6717; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@144765.4]
  assign _T_32938 = _T_38143 & _T_6740; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@144793.4]
  assign _T_32963 = _T_38143 & _T_6763; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@144821.4]
  assign _T_38177 = _T_42196 & _T_33985[222]; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@153362.4]
  assign _T_38178 = _T_38177 & _T_6089; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@153363.4]
  assign _T_33078 = _T_38178 & _T_6696; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@144939.4]
  assign _T_33101 = _T_38178 & _T_6717; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@144965.4]
  assign _T_33126 = _T_38178 & _T_6740; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@144993.4]
  assign _T_33151 = _T_38178 & _T_6763; // @[RegisterRouter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@145021.4]
  assign _GEN_2532 = 9'h1 == _T_33453 ? _T_6609 : _T_6609; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_2533 = 9'h2 == _T_33453 ? _T_6609 : _GEN_2532; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_2534 = 9'h3 == _T_33453 ? _T_6609 : _GEN_2533; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_2535 = 9'h4 == _T_33453 ? _T_6609 : _GEN_2534; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_2536 = 9'h5 == _T_33453 ? _T_6609 : _GEN_2535; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_2537 = 9'h6 == _T_33453 ? _T_6609 : _GEN_2536; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_2538 = 9'h7 == _T_33453 ? _T_6609 : _GEN_2537; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_2539 = 9'h8 == _T_33453 ? _T_6609 : _GEN_2538; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_2540 = 9'h9 == _T_33453 ? _T_6609 : _GEN_2539; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_2541 = 9'ha == _T_33453 ? _T_6609 : _GEN_2540; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_2542 = 9'hb == _T_33453 ? _T_6609 : _GEN_2541; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_2543 = 9'hc == _T_33453 ? _T_6609 : _GEN_2542; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_2544 = 9'hd == _T_33453 ? _T_6609 : _GEN_2543; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_2545 = 9'he == _T_33453 ? _T_6609 : _GEN_2544; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_2546 = 9'hf == _T_33453 ? _T_6609 : _GEN_2545; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_2547 = 9'h10 == _T_33453 ? _T_6609 : _GEN_2546; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_2548 = 9'h11 == _T_33453 ? _T_6609 : _GEN_2547; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_2549 = 9'h12 == _T_33453 ? _T_6609 : _GEN_2548; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_2550 = 9'h13 == _T_33453 ? _T_6609 : _GEN_2549; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_2551 = 9'h14 == _T_33453 ? _T_6609 : _GEN_2550; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_3672 = 9'h15 == _T_33453; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_2552 = _GEN_3672 | _GEN_2551; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_3673 = 9'h16 == _T_33453; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_2553 = _GEN_3673 | _GEN_2552; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_3674 = 9'h17 == _T_33453; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_2554 = _GEN_3674 | _GEN_2553; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_3675 = 9'h18 == _T_33453; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_2555 = _GEN_3675 | _GEN_2554; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_3676 = 9'h19 == _T_33453; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_2556 = _GEN_3676 | _GEN_2555; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_3677 = 9'h1a == _T_33453; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_2557 = _GEN_3677 | _GEN_2556; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_3678 = 9'h1b == _T_33453; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_2558 = _GEN_3678 | _GEN_2557; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_3679 = 9'h1c == _T_33453; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_2559 = _GEN_3679 | _GEN_2558; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_3680 = 9'h1d == _T_33453; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_2560 = _GEN_3680 | _GEN_2559; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_3681 = 9'h1e == _T_33453; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_2561 = _GEN_3681 | _GEN_2560; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_3682 = 9'h1f == _T_33453; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_2562 = _GEN_3682 | _GEN_2561; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_3683 = 9'h20 == _T_33453; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_2563 = _GEN_3683 | _GEN_2562; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_3684 = 9'h21 == _T_33453; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_2564 = _GEN_3684 | _GEN_2563; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_3685 = 9'h22 == _T_33453; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_2565 = _GEN_3685 | _GEN_2564; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_3686 = 9'h23 == _T_33453; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_2566 = _GEN_3686 | _GEN_2565; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_3687 = 9'h24 == _T_33453; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_2567 = _GEN_3687 | _GEN_2566; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_3688 = 9'h25 == _T_33453; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_2568 = _GEN_3688 | _GEN_2567; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_3689 = 9'h26 == _T_33453; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_2569 = _GEN_3689 | _GEN_2568; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_3690 = 9'h27 == _T_33453; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_2570 = _GEN_3690 | _GEN_2569; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_3691 = 9'h28 == _T_33453; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_2571 = _GEN_3691 | _GEN_2570; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_3692 = 9'h29 == _T_33453; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_2572 = _GEN_3692 | _GEN_2571; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_3693 = 9'h2a == _T_33453; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_2573 = _GEN_3693 | _GEN_2572; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_3694 = 9'h2b == _T_33453; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_2574 = _GEN_3694 | _GEN_2573; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_3695 = 9'h2c == _T_33453; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_2575 = _GEN_3695 | _GEN_2574; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_3696 = 9'h2d == _T_33453; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_2576 = _GEN_3696 | _GEN_2575; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_3697 = 9'h2e == _T_33453; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_2577 = _GEN_3697 | _GEN_2576; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_3698 = 9'h2f == _T_33453; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_2578 = _GEN_3698 | _GEN_2577; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_3699 = 9'h30 == _T_33453; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_2579 = _GEN_3699 | _GEN_2578; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_3700 = 9'h31 == _T_33453; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_2580 = _GEN_3700 | _GEN_2579; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_3701 = 9'h32 == _T_33453; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_2581 = _GEN_3701 | _GEN_2580; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_3702 = 9'h33 == _T_33453; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_2582 = _GEN_3702 | _GEN_2581; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_3703 = 9'h34 == _T_33453; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_2583 = _GEN_3703 | _GEN_2582; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_3704 = 9'h35 == _T_33453; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_2584 = _GEN_3704 | _GEN_2583; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_3705 = 9'h36 == _T_33453; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_2585 = _GEN_3705 | _GEN_2584; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_3706 = 9'h37 == _T_33453; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_2586 = _GEN_3706 | _GEN_2585; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_3707 = 9'h38 == _T_33453; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_2587 = _GEN_3707 | _GEN_2586; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_3708 = 9'h39 == _T_33453; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_2588 = _GEN_3708 | _GEN_2587; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_3709 = 9'h3a == _T_33453; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_2589 = _GEN_3709 | _GEN_2588; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_3710 = 9'h3b == _T_33453; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_2590 = _GEN_3710 | _GEN_2589; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_3711 = 9'h3c == _T_33453; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_2591 = _GEN_3711 | _GEN_2590; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_3712 = 9'h3d == _T_33453; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_2592 = _GEN_3712 | _GEN_2591; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_3713 = 9'h3e == _T_33453; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_2593 = _GEN_3713 | _GEN_2592; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_3714 = 9'h3f == _T_33453; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_2594 = _GEN_3714 | _GEN_2593; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_2595 = 9'h40 == _T_33453 ? _T_6089 : _GEN_2594; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_2596 = 9'h41 == _T_33453 ? _T_6089 : _GEN_2595; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_2597 = 9'h42 == _T_33453 ? _T_6089 : _GEN_2596; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_2598 = 9'h43 == _T_33453 ? _T_6089 : _GEN_2597; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_3715 = 9'h44 == _T_33453; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_2599 = _GEN_3715 | _GEN_2598; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_3716 = 9'h45 == _T_33453; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_2600 = _GEN_3716 | _GEN_2599; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_3717 = 9'h46 == _T_33453; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_2601 = _GEN_3717 | _GEN_2600; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_3718 = 9'h47 == _T_33453; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_2602 = _GEN_3718 | _GEN_2601; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_3719 = 9'h48 == _T_33453; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_2603 = _GEN_3719 | _GEN_2602; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_3720 = 9'h49 == _T_33453; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_2604 = _GEN_3720 | _GEN_2603; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_3721 = 9'h4a == _T_33453; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_2605 = _GEN_3721 | _GEN_2604; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_3722 = 9'h4b == _T_33453; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_2606 = _GEN_3722 | _GEN_2605; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_3723 = 9'h4c == _T_33453; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_2607 = _GEN_3723 | _GEN_2606; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_3724 = 9'h4d == _T_33453; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_2608 = _GEN_3724 | _GEN_2607; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_3725 = 9'h4e == _T_33453; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_2609 = _GEN_3725 | _GEN_2608; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_3726 = 9'h4f == _T_33453; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_2610 = _GEN_3726 | _GEN_2609; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_3727 = 9'h50 == _T_33453; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_2611 = _GEN_3727 | _GEN_2610; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_3728 = 9'h51 == _T_33453; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_2612 = _GEN_3728 | _GEN_2611; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_3729 = 9'h52 == _T_33453; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_2613 = _GEN_3729 | _GEN_2612; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_3730 = 9'h53 == _T_33453; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_2614 = _GEN_3730 | _GEN_2613; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_3731 = 9'h54 == _T_33453; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_2615 = _GEN_3731 | _GEN_2614; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_3732 = 9'h55 == _T_33453; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_2616 = _GEN_3732 | _GEN_2615; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_3733 = 9'h56 == _T_33453; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_2617 = _GEN_3733 | _GEN_2616; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_3734 = 9'h57 == _T_33453; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_2618 = _GEN_3734 | _GEN_2617; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_3735 = 9'h58 == _T_33453; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_2619 = _GEN_3735 | _GEN_2618; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_3736 = 9'h59 == _T_33453; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_2620 = _GEN_3736 | _GEN_2619; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_3737 = 9'h5a == _T_33453; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_2621 = _GEN_3737 | _GEN_2620; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_3738 = 9'h5b == _T_33453; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_2622 = _GEN_3738 | _GEN_2621; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_3739 = 9'h5c == _T_33453; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_2623 = _GEN_3739 | _GEN_2622; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_3740 = 9'h5d == _T_33453; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_2624 = _GEN_3740 | _GEN_2623; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_3741 = 9'h5e == _T_33453; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_2625 = _GEN_3741 | _GEN_2624; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_3742 = 9'h5f == _T_33453; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_2626 = _GEN_3742 | _GEN_2625; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_3743 = 9'h60 == _T_33453; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_2627 = _GEN_3743 | _GEN_2626; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_3744 = 9'h61 == _T_33453; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_2628 = _GEN_3744 | _GEN_2627; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_3745 = 9'h62 == _T_33453; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_2629 = _GEN_3745 | _GEN_2628; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_3746 = 9'h63 == _T_33453; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_2630 = _GEN_3746 | _GEN_2629; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_3747 = 9'h64 == _T_33453; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_2631 = _GEN_3747 | _GEN_2630; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_3748 = 9'h65 == _T_33453; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_2632 = _GEN_3748 | _GEN_2631; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_3749 = 9'h66 == _T_33453; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_2633 = _GEN_3749 | _GEN_2632; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_3750 = 9'h67 == _T_33453; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_2634 = _GEN_3750 | _GEN_2633; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_3751 = 9'h68 == _T_33453; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_2635 = _GEN_3751 | _GEN_2634; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_3752 = 9'h69 == _T_33453; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_2636 = _GEN_3752 | _GEN_2635; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_3753 = 9'h6a == _T_33453; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_2637 = _GEN_3753 | _GEN_2636; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_3754 = 9'h6b == _T_33453; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_2638 = _GEN_3754 | _GEN_2637; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_3755 = 9'h6c == _T_33453; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_2639 = _GEN_3755 | _GEN_2638; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_3756 = 9'h6d == _T_33453; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_2640 = _GEN_3756 | _GEN_2639; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_3757 = 9'h6e == _T_33453; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_2641 = _GEN_3757 | _GEN_2640; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_3758 = 9'h6f == _T_33453; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_2642 = _GEN_3758 | _GEN_2641; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_3759 = 9'h70 == _T_33453; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_2643 = _GEN_3759 | _GEN_2642; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_3760 = 9'h71 == _T_33453; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_2644 = _GEN_3760 | _GEN_2643; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_3761 = 9'h72 == _T_33453; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_2645 = _GEN_3761 | _GEN_2644; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_3762 = 9'h73 == _T_33453; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_2646 = _GEN_3762 | _GEN_2645; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_3763 = 9'h74 == _T_33453; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_2647 = _GEN_3763 | _GEN_2646; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_3764 = 9'h75 == _T_33453; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_2648 = _GEN_3764 | _GEN_2647; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_3765 = 9'h76 == _T_33453; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_2649 = _GEN_3765 | _GEN_2648; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_3766 = 9'h77 == _T_33453; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_2650 = _GEN_3766 | _GEN_2649; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_3767 = 9'h78 == _T_33453; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_2651 = _GEN_3767 | _GEN_2650; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_3768 = 9'h79 == _T_33453; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_2652 = _GEN_3768 | _GEN_2651; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_3769 = 9'h7a == _T_33453; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_2653 = _GEN_3769 | _GEN_2652; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_3770 = 9'h7b == _T_33453; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_2654 = _GEN_3770 | _GEN_2653; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_3771 = 9'h7c == _T_33453; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_2655 = _GEN_3771 | _GEN_2654; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_3772 = 9'h7d == _T_33453; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_2656 = _GEN_3772 | _GEN_2655; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_3773 = 9'h7e == _T_33453; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_2657 = _GEN_3773 | _GEN_2656; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_3774 = 9'h7f == _T_33453; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_2658 = _GEN_3774 | _GEN_2657; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_3775 = 9'h80 == _T_33453; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_2659 = _GEN_3775 | _GEN_2658; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_3776 = 9'h81 == _T_33453; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_2660 = _GEN_3776 | _GEN_2659; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_3777 = 9'h82 == _T_33453; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_2661 = _GEN_3777 | _GEN_2660; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_3778 = 9'h83 == _T_33453; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_2662 = _GEN_3778 | _GEN_2661; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_3779 = 9'h84 == _T_33453; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_2663 = _GEN_3779 | _GEN_2662; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_3780 = 9'h85 == _T_33453; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_2664 = _GEN_3780 | _GEN_2663; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_3781 = 9'h86 == _T_33453; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_2665 = _GEN_3781 | _GEN_2664; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_3782 = 9'h87 == _T_33453; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_2666 = _GEN_3782 | _GEN_2665; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_3783 = 9'h88 == _T_33453; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_2667 = _GEN_3783 | _GEN_2666; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_3784 = 9'h89 == _T_33453; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_2668 = _GEN_3784 | _GEN_2667; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_3785 = 9'h8a == _T_33453; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_2669 = _GEN_3785 | _GEN_2668; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_3786 = 9'h8b == _T_33453; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_2670 = _GEN_3786 | _GEN_2669; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_3787 = 9'h8c == _T_33453; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_2671 = _GEN_3787 | _GEN_2670; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_3788 = 9'h8d == _T_33453; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_2672 = _GEN_3788 | _GEN_2671; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_3789 = 9'h8e == _T_33453; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_2673 = _GEN_3789 | _GEN_2672; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_3790 = 9'h8f == _T_33453; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_2674 = _GEN_3790 | _GEN_2673; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_3791 = 9'h90 == _T_33453; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_2675 = _GEN_3791 | _GEN_2674; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_3792 = 9'h91 == _T_33453; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_2676 = _GEN_3792 | _GEN_2675; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_3793 = 9'h92 == _T_33453; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_2677 = _GEN_3793 | _GEN_2676; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_3794 = 9'h93 == _T_33453; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_2678 = _GEN_3794 | _GEN_2677; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_3795 = 9'h94 == _T_33453; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_2679 = _GEN_3795 | _GEN_2678; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_3796 = 9'h95 == _T_33453; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_2680 = _GEN_3796 | _GEN_2679; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_3797 = 9'h96 == _T_33453; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_2681 = _GEN_3797 | _GEN_2680; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_3798 = 9'h97 == _T_33453; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_2682 = _GEN_3798 | _GEN_2681; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_3799 = 9'h98 == _T_33453; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_2683 = _GEN_3799 | _GEN_2682; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_3800 = 9'h99 == _T_33453; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_2684 = _GEN_3800 | _GEN_2683; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_3801 = 9'h9a == _T_33453; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_2685 = _GEN_3801 | _GEN_2684; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_3802 = 9'h9b == _T_33453; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_2686 = _GEN_3802 | _GEN_2685; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_3803 = 9'h9c == _T_33453; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_2687 = _GEN_3803 | _GEN_2686; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_3804 = 9'h9d == _T_33453; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_2688 = _GEN_3804 | _GEN_2687; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_3805 = 9'h9e == _T_33453; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_2689 = _GEN_3805 | _GEN_2688; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_3806 = 9'h9f == _T_33453; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_2690 = _GEN_3806 | _GEN_2689; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_3807 = 9'ha0 == _T_33453; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_2691 = _GEN_3807 | _GEN_2690; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_3808 = 9'ha1 == _T_33453; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_2692 = _GEN_3808 | _GEN_2691; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_3809 = 9'ha2 == _T_33453; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_2693 = _GEN_3809 | _GEN_2692; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_3810 = 9'ha3 == _T_33453; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_2694 = _GEN_3810 | _GEN_2693; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_3811 = 9'ha4 == _T_33453; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_2695 = _GEN_3811 | _GEN_2694; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_3812 = 9'ha5 == _T_33453; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_2696 = _GEN_3812 | _GEN_2695; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_3813 = 9'ha6 == _T_33453; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_2697 = _GEN_3813 | _GEN_2696; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_3814 = 9'ha7 == _T_33453; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_2698 = _GEN_3814 | _GEN_2697; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_3815 = 9'ha8 == _T_33453; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_2699 = _GEN_3815 | _GEN_2698; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_3816 = 9'ha9 == _T_33453; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_2700 = _GEN_3816 | _GEN_2699; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_3817 = 9'haa == _T_33453; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_2701 = _GEN_3817 | _GEN_2700; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_3818 = 9'hab == _T_33453; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_2702 = _GEN_3818 | _GEN_2701; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_3819 = 9'hac == _T_33453; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_2703 = _GEN_3819 | _GEN_2702; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_3820 = 9'had == _T_33453; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_2704 = _GEN_3820 | _GEN_2703; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_3821 = 9'hae == _T_33453; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_2705 = _GEN_3821 | _GEN_2704; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_3822 = 9'haf == _T_33453; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_2706 = _GEN_3822 | _GEN_2705; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_3823 = 9'hb0 == _T_33453; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_2707 = _GEN_3823 | _GEN_2706; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_3824 = 9'hb1 == _T_33453; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_2708 = _GEN_3824 | _GEN_2707; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_3825 = 9'hb2 == _T_33453; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_2709 = _GEN_3825 | _GEN_2708; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_3826 = 9'hb3 == _T_33453; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_2710 = _GEN_3826 | _GEN_2709; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_3827 = 9'hb4 == _T_33453; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_2711 = _GEN_3827 | _GEN_2710; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_3828 = 9'hb5 == _T_33453; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_2712 = _GEN_3828 | _GEN_2711; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_3829 = 9'hb6 == _T_33453; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_2713 = _GEN_3829 | _GEN_2712; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_3830 = 9'hb7 == _T_33453; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_2714 = _GEN_3830 | _GEN_2713; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_3831 = 9'hb8 == _T_33453; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_2715 = _GEN_3831 | _GEN_2714; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_3832 = 9'hb9 == _T_33453; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_2716 = _GEN_3832 | _GEN_2715; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_3833 = 9'hba == _T_33453; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_2717 = _GEN_3833 | _GEN_2716; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_3834 = 9'hbb == _T_33453; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_2718 = _GEN_3834 | _GEN_2717; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_3835 = 9'hbc == _T_33453; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_2719 = _GEN_3835 | _GEN_2718; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_3836 = 9'hbd == _T_33453; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_2720 = _GEN_3836 | _GEN_2719; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_3837 = 9'hbe == _T_33453; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_2721 = _GEN_3837 | _GEN_2720; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_3838 = 9'hbf == _T_33453; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_2722 = _GEN_3838 | _GEN_2721; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_2723 = 9'hc0 == _T_33453 ? _T_6089 : _GEN_2722; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_3839 = 9'hc1 == _T_33453; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_2724 = _GEN_3839 | _GEN_2723; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_3840 = 9'hc2 == _T_33453; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_2725 = _GEN_3840 | _GEN_2724; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_3841 = 9'hc3 == _T_33453; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_2726 = _GEN_3841 | _GEN_2725; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_3842 = 9'hc4 == _T_33453; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_2727 = _GEN_3842 | _GEN_2726; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_3843 = 9'hc5 == _T_33453; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_2728 = _GEN_3843 | _GEN_2727; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_3844 = 9'hc6 == _T_33453; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_2729 = _GEN_3844 | _GEN_2728; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_3845 = 9'hc7 == _T_33453; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_2730 = _GEN_3845 | _GEN_2729; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_3846 = 9'hc8 == _T_33453; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_2731 = _GEN_3846 | _GEN_2730; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_3847 = 9'hc9 == _T_33453; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_2732 = _GEN_3847 | _GEN_2731; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_3848 = 9'hca == _T_33453; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_2733 = _GEN_3848 | _GEN_2732; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_3849 = 9'hcb == _T_33453; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_2734 = _GEN_3849 | _GEN_2733; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_3850 = 9'hcc == _T_33453; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_2735 = _GEN_3850 | _GEN_2734; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_3851 = 9'hcd == _T_33453; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_2736 = _GEN_3851 | _GEN_2735; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_2737 = 9'hce == _T_33453 ? _T_6089 : _GEN_2736; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_2738 = 9'hcf == _T_33453 ? _T_6089 : _GEN_2737; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_2739 = 9'hd0 == _T_33453 ? _T_6089 : _GEN_2738; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_2740 = 9'hd1 == _T_33453 ? _T_6089 : _GEN_2739; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_2741 = 9'hd2 == _T_33453 ? _T_6089 : _GEN_2740; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_2742 = 9'hd3 == _T_33453 ? _T_6089 : _GEN_2741; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_2743 = 9'hd4 == _T_33453 ? _T_6089 : _GEN_2742; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_2744 = 9'hd5 == _T_33453 ? _T_6089 : _GEN_2743; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_2745 = 9'hd6 == _T_33453 ? _T_6089 : _GEN_2744; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_2746 = 9'hd7 == _T_33453 ? _T_6089 : _GEN_2745; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_2747 = 9'hd8 == _T_33453 ? _T_6089 : _GEN_2746; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_2748 = 9'hd9 == _T_33453 ? _T_6089 : _GEN_2747; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_2749 = 9'hda == _T_33453 ? _T_6089 : _GEN_2748; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_2750 = 9'hdb == _T_33453 ? _T_6089 : _GEN_2749; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_2751 = 9'hdc == _T_33453 ? _T_6089 : _GEN_2750; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_2752 = 9'hdd == _T_33453 ? _T_6089 : _GEN_2751; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_2753 = 9'hde == _T_33453 ? _T_6089 : _GEN_2752; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_2754 = 9'hdf == _T_33453 ? _T_6089 : _GEN_2753; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_2755 = 9'he0 == _T_33453 ? _T_6089 : _GEN_2754; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_3852 = 9'he1 == _T_33453; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_2756 = _GEN_3852 | _GEN_2755; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_3853 = 9'he2 == _T_33453; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_2757 = _GEN_3853 | _GEN_2756; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_3854 = 9'he3 == _T_33453; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_2758 = _GEN_3854 | _GEN_2757; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_3855 = 9'he4 == _T_33453; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_2759 = _GEN_3855 | _GEN_2758; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_3856 = 9'he5 == _T_33453; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_2760 = _GEN_3856 | _GEN_2759; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_3857 = 9'he6 == _T_33453; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_2761 = _GEN_3857 | _GEN_2760; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_3858 = 9'he7 == _T_33453; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_2762 = _GEN_3858 | _GEN_2761; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_3859 = 9'he8 == _T_33453; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_2763 = _GEN_3859 | _GEN_2762; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_3860 = 9'he9 == _T_33453; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_2764 = _GEN_3860 | _GEN_2763; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_3861 = 9'hea == _T_33453; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_2765 = _GEN_3861 | _GEN_2764; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_3862 = 9'heb == _T_33453; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_2766 = _GEN_3862 | _GEN_2765; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_3863 = 9'hec == _T_33453; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_2767 = _GEN_3863 | _GEN_2766; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_3864 = 9'hed == _T_33453; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_2768 = _GEN_3864 | _GEN_2767; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_3865 = 9'hee == _T_33453; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_2769 = _GEN_3865 | _GEN_2768; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_3866 = 9'hef == _T_33453; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_2770 = _GEN_3866 | _GEN_2769; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_3867 = 9'hf0 == _T_33453; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_2771 = _GEN_3867 | _GEN_2770; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_3868 = 9'hf1 == _T_33453; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_2772 = _GEN_3868 | _GEN_2771; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_3869 = 9'hf2 == _T_33453; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_2773 = _GEN_3869 | _GEN_2772; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_3870 = 9'hf3 == _T_33453; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_2774 = _GEN_3870 | _GEN_2773; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_3871 = 9'hf4 == _T_33453; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_2775 = _GEN_3871 | _GEN_2774; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_3872 = 9'hf5 == _T_33453; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_2776 = _GEN_3872 | _GEN_2775; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_3873 = 9'hf6 == _T_33453; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_2777 = _GEN_3873 | _GEN_2776; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_3874 = 9'hf7 == _T_33453; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_2778 = _GEN_3874 | _GEN_2777; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_3875 = 9'hf8 == _T_33453; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_2779 = _GEN_3875 | _GEN_2778; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_3876 = 9'hf9 == _T_33453; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_2780 = _GEN_3876 | _GEN_2779; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_3877 = 9'hfa == _T_33453; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_2781 = _GEN_3877 | _GEN_2780; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_3878 = 9'hfb == _T_33453; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_2782 = _GEN_3878 | _GEN_2781; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_3879 = 9'hfc == _T_33453; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_2783 = _GEN_3879 | _GEN_2782; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_3880 = 9'hfd == _T_33453; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_2784 = _GEN_3880 | _GEN_2783; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_3881 = 9'hfe == _T_33453; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_2785 = _GEN_3881 | _GEN_2784; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_3882 = 9'hff == _T_33453; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_2786 = _GEN_3882 | _GEN_2785; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_2787 = 9'h100 == _T_33453 ? _T_6089 : _GEN_2786; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_2788 = 9'h101 == _T_33453 ? _T_6089 : _GEN_2787; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_2789 = 9'h102 == _T_33453 ? _T_6089 : _GEN_2788; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_2790 = 9'h103 == _T_33453 ? _T_6089 : _GEN_2789; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_2791 = 9'h104 == _T_33453 ? _T_6089 : _GEN_2790; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_2792 = 9'h105 == _T_33453 ? _T_6089 : _GEN_2791; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_2793 = 9'h106 == _T_33453 ? _T_6089 : _GEN_2792; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_2794 = 9'h107 == _T_33453 ? _T_6089 : _GEN_2793; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_2795 = 9'h108 == _T_33453 ? _T_6089 : _GEN_2794; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_2796 = 9'h109 == _T_33453 ? _T_6089 : _GEN_2795; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_2797 = 9'h10a == _T_33453 ? _T_6089 : _GEN_2796; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_2798 = 9'h10b == _T_33453 ? _T_6089 : _GEN_2797; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_2799 = 9'h10c == _T_33453 ? _T_6089 : _GEN_2798; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_2800 = 9'h10d == _T_33453 ? _T_6089 : _GEN_2799; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_2801 = 9'h10e == _T_33453 ? _T_6089 : _GEN_2800; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_2802 = 9'h10f == _T_33453 ? _T_6089 : _GEN_2801; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_2803 = 9'h110 == _T_33453 ? _T_6089 : _GEN_2802; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_2804 = 9'h111 == _T_33453 ? _T_6089 : _GEN_2803; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_2805 = 9'h112 == _T_33453 ? _T_6089 : _GEN_2804; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_2806 = 9'h113 == _T_33453 ? _T_6089 : _GEN_2805; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_2807 = 9'h114 == _T_33453 ? _T_6089 : _GEN_2806; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_2808 = 9'h115 == _T_33453 ? _T_6089 : _GEN_2807; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_2809 = 9'h116 == _T_33453 ? _T_6089 : _GEN_2808; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_2810 = 9'h117 == _T_33453 ? _T_6089 : _GEN_2809; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_2811 = 9'h118 == _T_33453 ? _T_6089 : _GEN_2810; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_2812 = 9'h119 == _T_33453 ? _T_6089 : _GEN_2811; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_2813 = 9'h11a == _T_33453 ? _T_6089 : _GEN_2812; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_2814 = 9'h11b == _T_33453 ? _T_6089 : _GEN_2813; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_2815 = 9'h11c == _T_33453 ? _T_6089 : _GEN_2814; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_2816 = 9'h11d == _T_33453 ? _T_6089 : _GEN_2815; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_2817 = 9'h11e == _T_33453 ? _T_6089 : _GEN_2816; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_2818 = 9'h11f == _T_33453 ? _T_6089 : _GEN_2817; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_2819 = 9'h120 == _T_33453 ? _T_6089 : _GEN_2818; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_2820 = 9'h121 == _T_33453 ? _T_6089 : _GEN_2819; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_2821 = 9'h122 == _T_33453 ? _T_6089 : _GEN_2820; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_2822 = 9'h123 == _T_33453 ? _T_6089 : _GEN_2821; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_2823 = 9'h124 == _T_33453 ? _T_6089 : _GEN_2822; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_2824 = 9'h125 == _T_33453 ? _T_6089 : _GEN_2823; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_2825 = 9'h126 == _T_33453 ? _T_6089 : _GEN_2824; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_2826 = 9'h127 == _T_33453 ? _T_6089 : _GEN_2825; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_2827 = 9'h128 == _T_33453 ? _T_6089 : _GEN_2826; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_2828 = 9'h129 == _T_33453 ? _T_6089 : _GEN_2827; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_2829 = 9'h12a == _T_33453 ? _T_6089 : _GEN_2828; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_2830 = 9'h12b == _T_33453 ? _T_6089 : _GEN_2829; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_2831 = 9'h12c == _T_33453 ? _T_6089 : _GEN_2830; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_2832 = 9'h12d == _T_33453 ? _T_6089 : _GEN_2831; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_2833 = 9'h12e == _T_33453 ? _T_6089 : _GEN_2832; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_2834 = 9'h12f == _T_33453 ? _T_6089 : _GEN_2833; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_2835 = 9'h130 == _T_33453 ? _T_6089 : _GEN_2834; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_2836 = 9'h131 == _T_33453 ? _T_6089 : _GEN_2835; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_2837 = 9'h132 == _T_33453 ? _T_6089 : _GEN_2836; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_2838 = 9'h133 == _T_33453 ? _T_6089 : _GEN_2837; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_2839 = 9'h134 == _T_33453 ? _T_6089 : _GEN_2838; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_2840 = 9'h135 == _T_33453 ? _T_6089 : _GEN_2839; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_2841 = 9'h136 == _T_33453 ? _T_6089 : _GEN_2840; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_2842 = 9'h137 == _T_33453 ? _T_6089 : _GEN_2841; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_2843 = 9'h138 == _T_33453 ? _T_6089 : _GEN_2842; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_2844 = 9'h139 == _T_33453 ? _T_6089 : _GEN_2843; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_2845 = 9'h13a == _T_33453 ? _T_6089 : _GEN_2844; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_2846 = 9'h13b == _T_33453 ? _T_6089 : _GEN_2845; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_2847 = 9'h13c == _T_33453 ? _T_6089 : _GEN_2846; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_2848 = 9'h13d == _T_33453 ? _T_6089 : _GEN_2847; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_2849 = 9'h13e == _T_33453 ? _T_6089 : _GEN_2848; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_2850 = 9'h13f == _T_33453 ? _T_6089 : _GEN_2849; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_2851 = 9'h140 == _T_33453 ? _T_6089 : _GEN_2850; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_2852 = 9'h141 == _T_33453 ? _T_6089 : _GEN_2851; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_2853 = 9'h142 == _T_33453 ? _T_6089 : _GEN_2852; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_2854 = 9'h143 == _T_33453 ? _T_6089 : _GEN_2853; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_2855 = 9'h144 == _T_33453 ? _T_6089 : _GEN_2854; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_2856 = 9'h145 == _T_33453 ? _T_6089 : _GEN_2855; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_2857 = 9'h146 == _T_33453 ? _T_6089 : _GEN_2856; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_2858 = 9'h147 == _T_33453 ? _T_6089 : _GEN_2857; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_2859 = 9'h148 == _T_33453 ? _T_6089 : _GEN_2858; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_2860 = 9'h149 == _T_33453 ? _T_6089 : _GEN_2859; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_2861 = 9'h14a == _T_33453 ? _T_6089 : _GEN_2860; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_2862 = 9'h14b == _T_33453 ? _T_6089 : _GEN_2861; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_2863 = 9'h14c == _T_33453 ? _T_6089 : _GEN_2862; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_2864 = 9'h14d == _T_33453 ? _T_6089 : _GEN_2863; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_2865 = 9'h14e == _T_33453 ? _T_6089 : _GEN_2864; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_2866 = 9'h14f == _T_33453 ? _T_6089 : _GEN_2865; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_2867 = 9'h150 == _T_33453 ? _T_6089 : _GEN_2866; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_2868 = 9'h151 == _T_33453 ? _T_6089 : _GEN_2867; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_2869 = 9'h152 == _T_33453 ? _T_6089 : _GEN_2868; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_2870 = 9'h153 == _T_33453 ? _T_6089 : _GEN_2869; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_2871 = 9'h154 == _T_33453 ? _T_6089 : _GEN_2870; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_2872 = 9'h155 == _T_33453 ? _T_6089 : _GEN_2871; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_2873 = 9'h156 == _T_33453 ? _T_6089 : _GEN_2872; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_2874 = 9'h157 == _T_33453 ? _T_6089 : _GEN_2873; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_2875 = 9'h158 == _T_33453 ? _T_6089 : _GEN_2874; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_2876 = 9'h159 == _T_33453 ? _T_6089 : _GEN_2875; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_2877 = 9'h15a == _T_33453 ? _T_6089 : _GEN_2876; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_2878 = 9'h15b == _T_33453 ? _T_6089 : _GEN_2877; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_2879 = 9'h15c == _T_33453 ? _T_6089 : _GEN_2878; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_2880 = 9'h15d == _T_33453 ? _T_6089 : _GEN_2879; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_2881 = 9'h15e == _T_33453 ? _T_6089 : _GEN_2880; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_2882 = 9'h15f == _T_33453 ? _T_6089 : _GEN_2881; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_2883 = 9'h160 == _T_33453 ? _T_6089 : _GEN_2882; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_2884 = 9'h161 == _T_33453 ? _T_6089 : _GEN_2883; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_2885 = 9'h162 == _T_33453 ? _T_6089 : _GEN_2884; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_2886 = 9'h163 == _T_33453 ? _T_6089 : _GEN_2885; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_2887 = 9'h164 == _T_33453 ? _T_6089 : _GEN_2886; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_2888 = 9'h165 == _T_33453 ? _T_6089 : _GEN_2887; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_2889 = 9'h166 == _T_33453 ? _T_6089 : _GEN_2888; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_2890 = 9'h167 == _T_33453 ? _T_6089 : _GEN_2889; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_2891 = 9'h168 == _T_33453 ? _T_6089 : _GEN_2890; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_2892 = 9'h169 == _T_33453 ? _T_6089 : _GEN_2891; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_2893 = 9'h16a == _T_33453 ? _T_6089 : _GEN_2892; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_2894 = 9'h16b == _T_33453 ? _T_6089 : _GEN_2893; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_2895 = 9'h16c == _T_33453 ? _T_6089 : _GEN_2894; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_2896 = 9'h16d == _T_33453 ? _T_6089 : _GEN_2895; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_2897 = 9'h16e == _T_33453 ? _T_6089 : _GEN_2896; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_2898 = 9'h16f == _T_33453 ? _T_6089 : _GEN_2897; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_2899 = 9'h170 == _T_33453 ? _T_6089 : _GEN_2898; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_2900 = 9'h171 == _T_33453 ? _T_6089 : _GEN_2899; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_2901 = 9'h172 == _T_33453 ? _T_6089 : _GEN_2900; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_2902 = 9'h173 == _T_33453 ? _T_6089 : _GEN_2901; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_2903 = 9'h174 == _T_33453 ? _T_6089 : _GEN_2902; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_2904 = 9'h175 == _T_33453 ? _T_6089 : _GEN_2903; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_2905 = 9'h176 == _T_33453 ? _T_6089 : _GEN_2904; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_2906 = 9'h177 == _T_33453 ? _T_6089 : _GEN_2905; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_2907 = 9'h178 == _T_33453 ? _T_6089 : _GEN_2906; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_2908 = 9'h179 == _T_33453 ? _T_6089 : _GEN_2907; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_2909 = 9'h17a == _T_33453 ? _T_6089 : _GEN_2908; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_2910 = 9'h17b == _T_33453 ? _T_6089 : _GEN_2909; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_2911 = 9'h17c == _T_33453 ? _T_6089 : _GEN_2910; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_2912 = 9'h17d == _T_33453 ? _T_6089 : _GEN_2911; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_2913 = 9'h17e == _T_33453 ? _T_6089 : _GEN_2912; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_2914 = 9'h17f == _T_33453 ? _T_6089 : _GEN_2913; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_2915 = 9'h180 == _T_33453 ? _T_6089 : _GEN_2914; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_2916 = 9'h181 == _T_33453 ? _T_6089 : _GEN_2915; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_2917 = 9'h182 == _T_33453 ? _T_6089 : _GEN_2916; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_2918 = 9'h183 == _T_33453 ? _T_6089 : _GEN_2917; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_2919 = 9'h184 == _T_33453 ? _T_6089 : _GEN_2918; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_2920 = 9'h185 == _T_33453 ? _T_6089 : _GEN_2919; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_2921 = 9'h186 == _T_33453 ? _T_6089 : _GEN_2920; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_2922 = 9'h187 == _T_33453 ? _T_6089 : _GEN_2921; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_2923 = 9'h188 == _T_33453 ? _T_6089 : _GEN_2922; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_2924 = 9'h189 == _T_33453 ? _T_6089 : _GEN_2923; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_2925 = 9'h18a == _T_33453 ? _T_6089 : _GEN_2924; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_2926 = 9'h18b == _T_33453 ? _T_6089 : _GEN_2925; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_2927 = 9'h18c == _T_33453 ? _T_6089 : _GEN_2926; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_2928 = 9'h18d == _T_33453 ? _T_6089 : _GEN_2927; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_2929 = 9'h18e == _T_33453 ? _T_6089 : _GEN_2928; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_2930 = 9'h18f == _T_33453 ? _T_6089 : _GEN_2929; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_2931 = 9'h190 == _T_33453 ? _T_6089 : _GEN_2930; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_2932 = 9'h191 == _T_33453 ? _T_6089 : _GEN_2931; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_2933 = 9'h192 == _T_33453 ? _T_6089 : _GEN_2932; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_2934 = 9'h193 == _T_33453 ? _T_6089 : _GEN_2933; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_2935 = 9'h194 == _T_33453 ? _T_6089 : _GEN_2934; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_2936 = 9'h195 == _T_33453 ? _T_6089 : _GEN_2935; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_2937 = 9'h196 == _T_33453 ? _T_6089 : _GEN_2936; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_2938 = 9'h197 == _T_33453 ? _T_6089 : _GEN_2937; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_2939 = 9'h198 == _T_33453 ? _T_6089 : _GEN_2938; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_2940 = 9'h199 == _T_33453 ? _T_6089 : _GEN_2939; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_2941 = 9'h19a == _T_33453 ? _T_6089 : _GEN_2940; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_2942 = 9'h19b == _T_33453 ? _T_6089 : _GEN_2941; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_2943 = 9'h19c == _T_33453 ? _T_6089 : _GEN_2942; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_2944 = 9'h19d == _T_33453 ? _T_6089 : _GEN_2943; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_2945 = 9'h19e == _T_33453 ? _T_6089 : _GEN_2944; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_2946 = 9'h19f == _T_33453 ? _T_6089 : _GEN_2945; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_2947 = 9'h1a0 == _T_33453 ? _T_6089 : _GEN_2946; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_2948 = 9'h1a1 == _T_33453 ? _T_6089 : _GEN_2947; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_2949 = 9'h1a2 == _T_33453 ? _T_6089 : _GEN_2948; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_2950 = 9'h1a3 == _T_33453 ? _T_6089 : _GEN_2949; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_2951 = 9'h1a4 == _T_33453 ? _T_6089 : _GEN_2950; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_2952 = 9'h1a5 == _T_33453 ? _T_6089 : _GEN_2951; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_2953 = 9'h1a6 == _T_33453 ? _T_6089 : _GEN_2952; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_2954 = 9'h1a7 == _T_33453 ? _T_6089 : _GEN_2953; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_2955 = 9'h1a8 == _T_33453 ? _T_6089 : _GEN_2954; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_2956 = 9'h1a9 == _T_33453 ? _T_6089 : _GEN_2955; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_2957 = 9'h1aa == _T_33453 ? _T_6089 : _GEN_2956; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_2958 = 9'h1ab == _T_33453 ? _T_6089 : _GEN_2957; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_2959 = 9'h1ac == _T_33453 ? _T_6089 : _GEN_2958; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_2960 = 9'h1ad == _T_33453 ? _T_6089 : _GEN_2959; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_2961 = 9'h1ae == _T_33453 ? _T_6089 : _GEN_2960; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_2962 = 9'h1af == _T_33453 ? _T_6089 : _GEN_2961; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_2963 = 9'h1b0 == _T_33453 ? _T_6089 : _GEN_2962; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_2964 = 9'h1b1 == _T_33453 ? _T_6089 : _GEN_2963; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_2965 = 9'h1b2 == _T_33453 ? _T_6089 : _GEN_2964; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_2966 = 9'h1b3 == _T_33453 ? _T_6089 : _GEN_2965; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_2967 = 9'h1b4 == _T_33453 ? _T_6089 : _GEN_2966; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_2968 = 9'h1b5 == _T_33453 ? _T_6089 : _GEN_2967; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_2969 = 9'h1b6 == _T_33453 ? _T_6089 : _GEN_2968; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_2970 = 9'h1b7 == _T_33453 ? _T_6089 : _GEN_2969; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_2971 = 9'h1b8 == _T_33453 ? _T_6089 : _GEN_2970; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_2972 = 9'h1b9 == _T_33453 ? _T_6089 : _GEN_2971; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_2973 = 9'h1ba == _T_33453 ? _T_6089 : _GEN_2972; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_2974 = 9'h1bb == _T_33453 ? _T_6089 : _GEN_2973; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_2975 = 9'h1bc == _T_33453 ? _T_6089 : _GEN_2974; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_2976 = 9'h1bd == _T_33453 ? _T_6089 : _GEN_2975; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_2977 = 9'h1be == _T_33453 ? _T_6089 : _GEN_2976; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_2978 = 9'h1bf == _T_33453 ? _T_6089 : _GEN_2977; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_2979 = 9'h1c0 == _T_33453 ? _T_6089 : _GEN_2978; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_2980 = 9'h1c1 == _T_33453 ? _T_6089 : _GEN_2979; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_2981 = 9'h1c2 == _T_33453 ? _T_6089 : _GEN_2980; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_2982 = 9'h1c3 == _T_33453 ? _T_6089 : _GEN_2981; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_2983 = 9'h1c4 == _T_33453 ? _T_6089 : _GEN_2982; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_2984 = 9'h1c5 == _T_33453 ? _T_6089 : _GEN_2983; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_2985 = 9'h1c6 == _T_33453 ? _T_6089 : _GEN_2984; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_2986 = 9'h1c7 == _T_33453 ? _T_6089 : _GEN_2985; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_2987 = 9'h1c8 == _T_33453 ? _T_6089 : _GEN_2986; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_2988 = 9'h1c9 == _T_33453 ? _T_6089 : _GEN_2987; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_2989 = 9'h1ca == _T_33453 ? _T_6089 : _GEN_2988; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_2990 = 9'h1cb == _T_33453 ? _T_6089 : _GEN_2989; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_2991 = 9'h1cc == _T_33453 ? _T_6089 : _GEN_2990; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_2992 = 9'h1cd == _T_33453 ? _T_6089 : _GEN_2991; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_2993 = 9'h1ce == _T_33453 ? _T_6089 : _GEN_2992; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_2994 = 9'h1cf == _T_33453 ? _T_6089 : _GEN_2993; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_2995 = 9'h1d0 == _T_33453 ? _T_6089 : _GEN_2994; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_2996 = 9'h1d1 == _T_33453 ? _T_6089 : _GEN_2995; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_2997 = 9'h1d2 == _T_33453 ? _T_6089 : _GEN_2996; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_2998 = 9'h1d3 == _T_33453 ? _T_6089 : _GEN_2997; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_2999 = 9'h1d4 == _T_33453 ? _T_6089 : _GEN_2998; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_3000 = 9'h1d5 == _T_33453 ? _T_6089 : _GEN_2999; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_3001 = 9'h1d6 == _T_33453 ? _T_6089 : _GEN_3000; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_3002 = 9'h1d7 == _T_33453 ? _T_6089 : _GEN_3001; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_3003 = 9'h1d8 == _T_33453 ? _T_6089 : _GEN_3002; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_3004 = 9'h1d9 == _T_33453 ? _T_6089 : _GEN_3003; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_3005 = 9'h1da == _T_33453 ? _T_6089 : _GEN_3004; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_3006 = 9'h1db == _T_33453 ? _T_6089 : _GEN_3005; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_3007 = 9'h1dc == _T_33453 ? _T_6089 : _GEN_3006; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_3008 = 9'h1dd == _T_33453 ? _T_6089 : _GEN_3007; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_3009 = 9'h1de == _T_33453 ? _T_6089 : _GEN_3008; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_3010 = 9'h1df == _T_33453 ? _T_6089 : _GEN_3009; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_3011 = 9'h1e0 == _T_33453 ? _T_6089 : _GEN_3010; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_3012 = 9'h1e1 == _T_33453 ? _T_6089 : _GEN_3011; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_3013 = 9'h1e2 == _T_33453 ? _T_6089 : _GEN_3012; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_3014 = 9'h1e3 == _T_33453 ? _T_6089 : _GEN_3013; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_3015 = 9'h1e4 == _T_33453 ? _T_6089 : _GEN_3014; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_3016 = 9'h1e5 == _T_33453 ? _T_6089 : _GEN_3015; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_3017 = 9'h1e6 == _T_33453 ? _T_6089 : _GEN_3016; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_3018 = 9'h1e7 == _T_33453 ? _T_6089 : _GEN_3017; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_3019 = 9'h1e8 == _T_33453 ? _T_6089 : _GEN_3018; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_3020 = 9'h1e9 == _T_33453 ? _T_6089 : _GEN_3019; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_3021 = 9'h1ea == _T_33453 ? _T_6089 : _GEN_3020; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_3022 = 9'h1eb == _T_33453 ? _T_6089 : _GEN_3021; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_3023 = 9'h1ec == _T_33453 ? _T_6089 : _GEN_3022; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_3024 = 9'h1ed == _T_33453 ? _T_6089 : _GEN_3023; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_3025 = 9'h1ee == _T_33453 ? _T_6089 : _GEN_3024; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_3026 = 9'h1ef == _T_33453 ? _T_6089 : _GEN_3025; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_3027 = 9'h1f0 == _T_33453 ? _T_6089 : _GEN_3026; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_3028 = 9'h1f1 == _T_33453 ? _T_6089 : _GEN_3027; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_3029 = 9'h1f2 == _T_33453 ? _T_6089 : _GEN_3028; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_3030 = 9'h1f3 == _T_33453 ? _T_6089 : _GEN_3029; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_3031 = 9'h1f4 == _T_33453 ? _T_6089 : _GEN_3030; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_3032 = 9'h1f5 == _T_33453 ? _T_6089 : _GEN_3031; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_3033 = 9'h1f6 == _T_33453 ? _T_6089 : _GEN_3032; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_3034 = 9'h1f7 == _T_33453 ? _T_6089 : _GEN_3033; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_3035 = 9'h1f8 == _T_33453 ? _T_6089 : _GEN_3034; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_3036 = 9'h1f9 == _T_33453 ? _T_6089 : _GEN_3035; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_3037 = 9'h1fa == _T_33453 ? _T_6089 : _GEN_3036; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_3038 = 9'h1fb == _T_33453 ? _T_6089 : _GEN_3037; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_3039 = 9'h1fc == _T_33453 ? _T_6089 : _GEN_3038; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_3040 = 9'h1fd == _T_33453 ? _T_6089 : _GEN_3039; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_3041 = 9'h1fe == _T_33453 ? _T_6089 : _GEN_3040; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_3042 = 9'h1ff == _T_33453 ? _T_6089 : _GEN_3041; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168039.4]
  assign _GEN_3044 = 9'h1 == _T_33453 ? 32'h380006f : 32'hc0006f; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  assign _GEN_3045 = 9'h2 == _T_33453 ? 32'h440006f : _GEN_3044; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  assign _GEN_3046 = 9'h3 == _T_33453 ? 32'hff0000f : _GEN_3045; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  assign _GEN_3047 = 9'h4 == _T_33453 ? 32'h7b241073 : _GEN_3046; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  assign _GEN_3048 = 9'h5 == _T_33453 ? 32'hf1402473 : _GEN_3047; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  assign _GEN_3049 = 9'h6 == _T_33453 ? 32'h10802023 : _GEN_3048; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  assign _GEN_3050 = 9'h7 == _T_33453 ? 32'h40044403 : _GEN_3049; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  assign _GEN_3051 = 9'h8 == _T_33453 ? 32'h347413 : _GEN_3050; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  assign _GEN_3052 = 9'h9 == _T_33453 ? 32'hfe0408e3 : _GEN_3051; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  assign _GEN_3053 = 9'ha == _T_33453 ? 32'h147413 : _GEN_3052; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  assign _GEN_3054 = 9'hb == _T_33453 ? 32'h40863 : _GEN_3053; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  assign _GEN_3055 = 9'hc == _T_33453 ? 32'h7b202473 : _GEN_3054; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  assign _GEN_3056 = 9'hd == _T_33453 ? 32'h10002223 : _GEN_3055; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  assign _GEN_3057 = 9'he == _T_33453 ? 32'h30000067 : _GEN_3056; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  assign _GEN_3058 = 9'hf == _T_33453 ? 32'hf1402473 : _GEN_3057; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  assign _GEN_3059 = 9'h10 == _T_33453 ? 32'h10802423 : _GEN_3058; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  assign _GEN_3060 = 9'h11 == _T_33453 ? 32'h7b202473 : _GEN_3059; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  assign _GEN_3061 = 9'h12 == _T_33453 ? 32'h7b200073 : _GEN_3060; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  assign _GEN_3062 = 9'h13 == _T_33453 ? 32'h10002623 : _GEN_3061; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  assign _GEN_3063 = 9'h14 == _T_33453 ? 32'h100073 : _GEN_3062; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  assign _GEN_3064 = 9'h15 == _T_33453 ? 32'h0 : _GEN_3063; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  assign _GEN_3065 = 9'h16 == _T_33453 ? 32'h0 : _GEN_3064; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  assign _GEN_3066 = 9'h17 == _T_33453 ? 32'h0 : _GEN_3065; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  assign _GEN_3067 = 9'h18 == _T_33453 ? 32'h0 : _GEN_3066; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  assign _GEN_3068 = 9'h19 == _T_33453 ? 32'h0 : _GEN_3067; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  assign _GEN_3069 = 9'h1a == _T_33453 ? 32'h0 : _GEN_3068; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  assign _GEN_3070 = 9'h1b == _T_33453 ? 32'h0 : _GEN_3069; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  assign _GEN_3071 = 9'h1c == _T_33453 ? 32'h0 : _GEN_3070; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  assign _GEN_3072 = 9'h1d == _T_33453 ? 32'h0 : _GEN_3071; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  assign _GEN_3073 = 9'h1e == _T_33453 ? 32'h0 : _GEN_3072; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  assign _GEN_3074 = 9'h1f == _T_33453 ? 32'h0 : _GEN_3073; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  assign _GEN_3075 = 9'h20 == _T_33453 ? 32'h0 : _GEN_3074; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  assign _GEN_3076 = 9'h21 == _T_33453 ? 32'h0 : _GEN_3075; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  assign _GEN_3077 = 9'h22 == _T_33453 ? 32'h0 : _GEN_3076; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  assign _GEN_3078 = 9'h23 == _T_33453 ? 32'h0 : _GEN_3077; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  assign _GEN_3079 = 9'h24 == _T_33453 ? 32'h0 : _GEN_3078; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  assign _GEN_3080 = 9'h25 == _T_33453 ? 32'h0 : _GEN_3079; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  assign _GEN_3081 = 9'h26 == _T_33453 ? 32'h0 : _GEN_3080; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  assign _GEN_3082 = 9'h27 == _T_33453 ? 32'h0 : _GEN_3081; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  assign _GEN_3083 = 9'h28 == _T_33453 ? 32'h0 : _GEN_3082; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  assign _GEN_3084 = 9'h29 == _T_33453 ? 32'h0 : _GEN_3083; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  assign _GEN_3085 = 9'h2a == _T_33453 ? 32'h0 : _GEN_3084; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  assign _GEN_3086 = 9'h2b == _T_33453 ? 32'h0 : _GEN_3085; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  assign _GEN_3087 = 9'h2c == _T_33453 ? 32'h0 : _GEN_3086; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  assign _GEN_3088 = 9'h2d == _T_33453 ? 32'h0 : _GEN_3087; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  assign _GEN_3089 = 9'h2e == _T_33453 ? 32'h0 : _GEN_3088; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  assign _GEN_3090 = 9'h2f == _T_33453 ? 32'h0 : _GEN_3089; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  assign _GEN_3091 = 9'h30 == _T_33453 ? 32'h0 : _GEN_3090; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  assign _GEN_3092 = 9'h31 == _T_33453 ? 32'h0 : _GEN_3091; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  assign _GEN_3093 = 9'h32 == _T_33453 ? 32'h0 : _GEN_3092; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  assign _GEN_3094 = 9'h33 == _T_33453 ? 32'h0 : _GEN_3093; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  assign _GEN_3095 = 9'h34 == _T_33453 ? 32'h0 : _GEN_3094; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  assign _GEN_3096 = 9'h35 == _T_33453 ? 32'h0 : _GEN_3095; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  assign _GEN_3097 = 9'h36 == _T_33453 ? 32'h0 : _GEN_3096; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  assign _GEN_3098 = 9'h37 == _T_33453 ? 32'h0 : _GEN_3097; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  assign _GEN_3099 = 9'h38 == _T_33453 ? 32'h0 : _GEN_3098; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  assign _GEN_3100 = 9'h39 == _T_33453 ? 32'h0 : _GEN_3099; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  assign _GEN_3101 = 9'h3a == _T_33453 ? 32'h0 : _GEN_3100; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  assign _GEN_3102 = 9'h3b == _T_33453 ? 32'h0 : _GEN_3101; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  assign _GEN_3103 = 9'h3c == _T_33453 ? 32'h0 : _GEN_3102; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  assign _GEN_3104 = 9'h3d == _T_33453 ? 32'h0 : _GEN_3103; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  assign _GEN_3105 = 9'h3e == _T_33453 ? 32'h0 : _GEN_3104; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  assign _GEN_3106 = 9'h3f == _T_33453 ? 32'h0 : _GEN_3105; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  assign _GEN_3107 = 9'h40 == _T_33453 ? 32'h0 : _GEN_3106; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  assign _GEN_3108 = 9'h41 == _T_33453 ? 32'h0 : _GEN_3107; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  assign _GEN_3109 = 9'h42 == _T_33453 ? 32'h0 : _GEN_3108; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  assign _GEN_3110 = 9'h43 == _T_33453 ? 32'h0 : _GEN_3109; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  assign _GEN_3111 = 9'h44 == _T_33453 ? 32'h0 : _GEN_3110; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  assign _GEN_3112 = 9'h45 == _T_33453 ? 32'h0 : _GEN_3111; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  assign _GEN_3113 = 9'h46 == _T_33453 ? 32'h0 : _GEN_3112; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  assign _GEN_3114 = 9'h47 == _T_33453 ? 32'h0 : _GEN_3113; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  assign _GEN_3115 = 9'h48 == _T_33453 ? 32'h0 : _GEN_3114; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  assign _GEN_3116 = 9'h49 == _T_33453 ? 32'h0 : _GEN_3115; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  assign _GEN_3117 = 9'h4a == _T_33453 ? 32'h0 : _GEN_3116; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  assign _GEN_3118 = 9'h4b == _T_33453 ? 32'h0 : _GEN_3117; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  assign _GEN_3119 = 9'h4c == _T_33453 ? 32'h0 : _GEN_3118; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  assign _GEN_3120 = 9'h4d == _T_33453 ? 32'h0 : _GEN_3119; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  assign _GEN_3121 = 9'h4e == _T_33453 ? 32'h0 : _GEN_3120; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  assign _GEN_3122 = 9'h4f == _T_33453 ? 32'h0 : _GEN_3121; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  assign _GEN_3123 = 9'h50 == _T_33453 ? 32'h0 : _GEN_3122; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  assign _GEN_3124 = 9'h51 == _T_33453 ? 32'h0 : _GEN_3123; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  assign _GEN_3125 = 9'h52 == _T_33453 ? 32'h0 : _GEN_3124; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  assign _GEN_3126 = 9'h53 == _T_33453 ? 32'h0 : _GEN_3125; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  assign _GEN_3127 = 9'h54 == _T_33453 ? 32'h0 : _GEN_3126; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  assign _GEN_3128 = 9'h55 == _T_33453 ? 32'h0 : _GEN_3127; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  assign _GEN_3129 = 9'h56 == _T_33453 ? 32'h0 : _GEN_3128; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  assign _GEN_3130 = 9'h57 == _T_33453 ? 32'h0 : _GEN_3129; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  assign _GEN_3131 = 9'h58 == _T_33453 ? 32'h0 : _GEN_3130; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  assign _GEN_3132 = 9'h59 == _T_33453 ? 32'h0 : _GEN_3131; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  assign _GEN_3133 = 9'h5a == _T_33453 ? 32'h0 : _GEN_3132; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  assign _GEN_3134 = 9'h5b == _T_33453 ? 32'h0 : _GEN_3133; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  assign _GEN_3135 = 9'h5c == _T_33453 ? 32'h0 : _GEN_3134; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  assign _GEN_3136 = 9'h5d == _T_33453 ? 32'h0 : _GEN_3135; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  assign _GEN_3137 = 9'h5e == _T_33453 ? 32'h0 : _GEN_3136; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  assign _GEN_3138 = 9'h5f == _T_33453 ? 32'h0 : _GEN_3137; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  assign _GEN_3139 = 9'h60 == _T_33453 ? 32'h0 : _GEN_3138; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  assign _GEN_3140 = 9'h61 == _T_33453 ? 32'h0 : _GEN_3139; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  assign _GEN_3141 = 9'h62 == _T_33453 ? 32'h0 : _GEN_3140; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  assign _GEN_3142 = 9'h63 == _T_33453 ? 32'h0 : _GEN_3141; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  assign _GEN_3143 = 9'h64 == _T_33453 ? 32'h0 : _GEN_3142; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  assign _GEN_3144 = 9'h65 == _T_33453 ? 32'h0 : _GEN_3143; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  assign _GEN_3145 = 9'h66 == _T_33453 ? 32'h0 : _GEN_3144; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  assign _GEN_3146 = 9'h67 == _T_33453 ? 32'h0 : _GEN_3145; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  assign _GEN_3147 = 9'h68 == _T_33453 ? 32'h0 : _GEN_3146; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  assign _GEN_3148 = 9'h69 == _T_33453 ? 32'h0 : _GEN_3147; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  assign _GEN_3149 = 9'h6a == _T_33453 ? 32'h0 : _GEN_3148; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  assign _GEN_3150 = 9'h6b == _T_33453 ? 32'h0 : _GEN_3149; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  assign _GEN_3151 = 9'h6c == _T_33453 ? 32'h0 : _GEN_3150; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  assign _GEN_3152 = 9'h6d == _T_33453 ? 32'h0 : _GEN_3151; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  assign _GEN_3153 = 9'h6e == _T_33453 ? 32'h0 : _GEN_3152; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  assign _GEN_3154 = 9'h6f == _T_33453 ? 32'h0 : _GEN_3153; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  assign _GEN_3155 = 9'h70 == _T_33453 ? 32'h0 : _GEN_3154; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  assign _GEN_3156 = 9'h71 == _T_33453 ? 32'h0 : _GEN_3155; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  assign _GEN_3157 = 9'h72 == _T_33453 ? 32'h0 : _GEN_3156; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  assign _GEN_3158 = 9'h73 == _T_33453 ? 32'h0 : _GEN_3157; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  assign _GEN_3159 = 9'h74 == _T_33453 ? 32'h0 : _GEN_3158; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  assign _GEN_3160 = 9'h75 == _T_33453 ? 32'h0 : _GEN_3159; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  assign _GEN_3161 = 9'h76 == _T_33453 ? 32'h0 : _GEN_3160; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  assign _GEN_3162 = 9'h77 == _T_33453 ? 32'h0 : _GEN_3161; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  assign _GEN_3163 = 9'h78 == _T_33453 ? 32'h0 : _GEN_3162; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  assign _GEN_3164 = 9'h79 == _T_33453 ? 32'h0 : _GEN_3163; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  assign _GEN_3165 = 9'h7a == _T_33453 ? 32'h0 : _GEN_3164; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  assign _GEN_3166 = 9'h7b == _T_33453 ? 32'h0 : _GEN_3165; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  assign _GEN_3167 = 9'h7c == _T_33453 ? 32'h0 : _GEN_3166; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  assign _GEN_3168 = 9'h7d == _T_33453 ? 32'h0 : _GEN_3167; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  assign _GEN_3169 = 9'h7e == _T_33453 ? 32'h0 : _GEN_3168; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  assign _GEN_3170 = 9'h7f == _T_33453 ? 32'h0 : _GEN_3169; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  assign _GEN_3171 = 9'h80 == _T_33453 ? 32'h0 : _GEN_3170; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  assign _GEN_3172 = 9'h81 == _T_33453 ? 32'h0 : _GEN_3171; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  assign _GEN_3173 = 9'h82 == _T_33453 ? 32'h0 : _GEN_3172; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  assign _GEN_3174 = 9'h83 == _T_33453 ? 32'h0 : _GEN_3173; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  assign _GEN_3175 = 9'h84 == _T_33453 ? 32'h0 : _GEN_3174; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  assign _GEN_3176 = 9'h85 == _T_33453 ? 32'h0 : _GEN_3175; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  assign _GEN_3177 = 9'h86 == _T_33453 ? 32'h0 : _GEN_3176; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  assign _GEN_3178 = 9'h87 == _T_33453 ? 32'h0 : _GEN_3177; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  assign _GEN_3179 = 9'h88 == _T_33453 ? 32'h0 : _GEN_3178; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  assign _GEN_3180 = 9'h89 == _T_33453 ? 32'h0 : _GEN_3179; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  assign _GEN_3181 = 9'h8a == _T_33453 ? 32'h0 : _GEN_3180; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  assign _GEN_3182 = 9'h8b == _T_33453 ? 32'h0 : _GEN_3181; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  assign _GEN_3183 = 9'h8c == _T_33453 ? 32'h0 : _GEN_3182; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  assign _GEN_3184 = 9'h8d == _T_33453 ? 32'h0 : _GEN_3183; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  assign _GEN_3185 = 9'h8e == _T_33453 ? 32'h0 : _GEN_3184; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  assign _GEN_3186 = 9'h8f == _T_33453 ? 32'h0 : _GEN_3185; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  assign _GEN_3187 = 9'h90 == _T_33453 ? 32'h0 : _GEN_3186; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  assign _GEN_3188 = 9'h91 == _T_33453 ? 32'h0 : _GEN_3187; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  assign _GEN_3189 = 9'h92 == _T_33453 ? 32'h0 : _GEN_3188; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  assign _GEN_3190 = 9'h93 == _T_33453 ? 32'h0 : _GEN_3189; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  assign _GEN_3191 = 9'h94 == _T_33453 ? 32'h0 : _GEN_3190; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  assign _GEN_3192 = 9'h95 == _T_33453 ? 32'h0 : _GEN_3191; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  assign _GEN_3193 = 9'h96 == _T_33453 ? 32'h0 : _GEN_3192; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  assign _GEN_3194 = 9'h97 == _T_33453 ? 32'h0 : _GEN_3193; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  assign _GEN_3195 = 9'h98 == _T_33453 ? 32'h0 : _GEN_3194; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  assign _GEN_3196 = 9'h99 == _T_33453 ? 32'h0 : _GEN_3195; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  assign _GEN_3197 = 9'h9a == _T_33453 ? 32'h0 : _GEN_3196; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  assign _GEN_3198 = 9'h9b == _T_33453 ? 32'h0 : _GEN_3197; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  assign _GEN_3199 = 9'h9c == _T_33453 ? 32'h0 : _GEN_3198; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  assign _GEN_3200 = 9'h9d == _T_33453 ? 32'h0 : _GEN_3199; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  assign _GEN_3201 = 9'h9e == _T_33453 ? 32'h0 : _GEN_3200; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  assign _GEN_3202 = 9'h9f == _T_33453 ? 32'h0 : _GEN_3201; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  assign _GEN_3203 = 9'ha0 == _T_33453 ? 32'h0 : _GEN_3202; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  assign _GEN_3204 = 9'ha1 == _T_33453 ? 32'h0 : _GEN_3203; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  assign _GEN_3205 = 9'ha2 == _T_33453 ? 32'h0 : _GEN_3204; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  assign _GEN_3206 = 9'ha3 == _T_33453 ? 32'h0 : _GEN_3205; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  assign _GEN_3207 = 9'ha4 == _T_33453 ? 32'h0 : _GEN_3206; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  assign _GEN_3208 = 9'ha5 == _T_33453 ? 32'h0 : _GEN_3207; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  assign _GEN_3209 = 9'ha6 == _T_33453 ? 32'h0 : _GEN_3208; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  assign _GEN_3210 = 9'ha7 == _T_33453 ? 32'h0 : _GEN_3209; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  assign _GEN_3211 = 9'ha8 == _T_33453 ? 32'h0 : _GEN_3210; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  assign _GEN_3212 = 9'ha9 == _T_33453 ? 32'h0 : _GEN_3211; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  assign _GEN_3213 = 9'haa == _T_33453 ? 32'h0 : _GEN_3212; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  assign _GEN_3214 = 9'hab == _T_33453 ? 32'h0 : _GEN_3213; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  assign _GEN_3215 = 9'hac == _T_33453 ? 32'h0 : _GEN_3214; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  assign _GEN_3216 = 9'had == _T_33453 ? 32'h0 : _GEN_3215; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  assign _GEN_3217 = 9'hae == _T_33453 ? 32'h0 : _GEN_3216; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  assign _GEN_3218 = 9'haf == _T_33453 ? 32'h0 : _GEN_3217; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  assign _GEN_3219 = 9'hb0 == _T_33453 ? 32'h0 : _GEN_3218; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  assign _GEN_3220 = 9'hb1 == _T_33453 ? 32'h0 : _GEN_3219; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  assign _GEN_3221 = 9'hb2 == _T_33453 ? 32'h0 : _GEN_3220; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  assign _GEN_3222 = 9'hb3 == _T_33453 ? 32'h0 : _GEN_3221; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  assign _GEN_3223 = 9'hb4 == _T_33453 ? 32'h0 : _GEN_3222; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  assign _GEN_3224 = 9'hb5 == _T_33453 ? 32'h0 : _GEN_3223; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  assign _GEN_3225 = 9'hb6 == _T_33453 ? 32'h0 : _GEN_3224; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  assign _GEN_3226 = 9'hb7 == _T_33453 ? 32'h0 : _GEN_3225; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  assign _GEN_3227 = 9'hb8 == _T_33453 ? 32'h0 : _GEN_3226; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  assign _GEN_3228 = 9'hb9 == _T_33453 ? 32'h0 : _GEN_3227; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  assign _GEN_3229 = 9'hba == _T_33453 ? 32'h0 : _GEN_3228; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  assign _GEN_3230 = 9'hbb == _T_33453 ? 32'h0 : _GEN_3229; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  assign _GEN_3231 = 9'hbc == _T_33453 ? 32'h0 : _GEN_3230; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  assign _GEN_3232 = 9'hbd == _T_33453 ? 32'h0 : _GEN_3231; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  assign _GEN_3233 = 9'hbe == _T_33453 ? 32'h0 : _GEN_3232; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  assign _GEN_3234 = 9'hbf == _T_33453 ? 32'h0 : _GEN_3233; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  assign _GEN_3235 = 9'hc0 == _T_33453 ? 32'h380006f : _GEN_3234; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  assign _GEN_3236 = 9'hc1 == _T_33453 ? 32'h0 : _GEN_3235; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  assign _GEN_3237 = 9'hc2 == _T_33453 ? 32'h0 : _GEN_3236; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  assign _GEN_3238 = 9'hc3 == _T_33453 ? 32'h0 : _GEN_3237; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  assign _GEN_3239 = 9'hc4 == _T_33453 ? 32'h0 : _GEN_3238; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  assign _GEN_3240 = 9'hc5 == _T_33453 ? 32'h0 : _GEN_3239; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  assign _GEN_3241 = 9'hc6 == _T_33453 ? 32'h0 : _GEN_3240; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  assign _GEN_3242 = 9'hc7 == _T_33453 ? 32'h0 : _GEN_3241; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  assign _GEN_3243 = 9'hc8 == _T_33453 ? 32'h0 : _GEN_3242; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  assign _GEN_3244 = 9'hc9 == _T_33453 ? 32'h0 : _GEN_3243; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  assign _GEN_3245 = 9'hca == _T_33453 ? 32'h0 : _GEN_3244; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  assign _GEN_3246 = 9'hcb == _T_33453 ? 32'h0 : _GEN_3245; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  assign _GEN_3247 = 9'hcc == _T_33453 ? 32'h0 : _GEN_3246; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  assign _GEN_3248 = 9'hcd == _T_33453 ? 32'h0 : _GEN_3247; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  assign _GEN_3249 = 9'hce == _T_33453 ? abstractGeneratedMem_0 : _GEN_3248; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  assign _GEN_3250 = 9'hcf == _T_33453 ? abstractGeneratedMem_1 : _GEN_3249; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  assign _GEN_3251 = 9'hd0 == _T_33453 ? _T_1223 : _GEN_3250; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  assign _GEN_3252 = 9'hd1 == _T_33453 ? _T_1027 : _GEN_3251; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  assign _GEN_3253 = 9'hd2 == _T_33453 ? _T_1321 : _GEN_3252; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  assign _GEN_3254 = 9'hd3 == _T_33453 ? _T_2330 : _GEN_3253; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  assign _GEN_3255 = 9'hd4 == _T_33453 ? _T_2760 : _GEN_3254; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  assign _GEN_3256 = 9'hd5 == _T_33453 ? _T_733 : _GEN_3255; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  assign _GEN_3257 = 9'hd6 == _T_33453 ? _T_929 : _GEN_3256; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  assign _GEN_3258 = 9'hd7 == _T_33453 ? _T_2232 : _GEN_3257; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  assign _GEN_3259 = 9'hd8 == _T_33453 ? _T_2639 : _GEN_3258; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  assign _GEN_3260 = 9'hd9 == _T_33453 ? _T_1125 : _GEN_3259; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  assign _GEN_3261 = 9'hda == _T_33453 ? _T_564 : _GEN_3260; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  assign _GEN_3262 = 9'hdb == _T_33453 ? _T_2541 : _GEN_3261; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  assign _GEN_3263 = 9'hdc == _T_33453 ? _T_2134 : _GEN_3262; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  assign _GEN_3264 = 9'hdd == _T_33453 ? _T_1419 : _GEN_3263; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  assign _GEN_3265 = 9'hde == _T_33453 ? _T_831 : _GEN_3264; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  assign _GEN_3266 = 9'hdf == _T_33453 ? _T_2977 : _GEN_3265; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  assign _GEN_3267 = 9'he0 == _T_33453 ? _T_2879 : _GEN_3266; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  assign _GEN_3268 = 9'he1 == _T_33453 ? 32'h0 : _GEN_3267; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  assign _GEN_3269 = 9'he2 == _T_33453 ? 32'h0 : _GEN_3268; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  assign _GEN_3270 = 9'he3 == _T_33453 ? 32'h0 : _GEN_3269; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  assign _GEN_3271 = 9'he4 == _T_33453 ? 32'h0 : _GEN_3270; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  assign _GEN_3272 = 9'he5 == _T_33453 ? 32'h0 : _GEN_3271; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  assign _GEN_3273 = 9'he6 == _T_33453 ? 32'h0 : _GEN_3272; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  assign _GEN_3274 = 9'he7 == _T_33453 ? 32'h0 : _GEN_3273; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  assign _GEN_3275 = 9'he8 == _T_33453 ? 32'h0 : _GEN_3274; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  assign _GEN_3276 = 9'he9 == _T_33453 ? 32'h0 : _GEN_3275; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  assign _GEN_3277 = 9'hea == _T_33453 ? 32'h0 : _GEN_3276; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  assign _GEN_3278 = 9'heb == _T_33453 ? 32'h0 : _GEN_3277; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  assign _GEN_3279 = 9'hec == _T_33453 ? 32'h0 : _GEN_3278; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  assign _GEN_3280 = 9'hed == _T_33453 ? 32'h0 : _GEN_3279; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  assign _GEN_3281 = 9'hee == _T_33453 ? 32'h0 : _GEN_3280; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  assign _GEN_3282 = 9'hef == _T_33453 ? 32'h0 : _GEN_3281; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  assign _GEN_3283 = 9'hf0 == _T_33453 ? 32'h0 : _GEN_3282; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  assign _GEN_3284 = 9'hf1 == _T_33453 ? 32'h0 : _GEN_3283; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  assign _GEN_3285 = 9'hf2 == _T_33453 ? 32'h0 : _GEN_3284; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  assign _GEN_3286 = 9'hf3 == _T_33453 ? 32'h0 : _GEN_3285; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  assign _GEN_3287 = 9'hf4 == _T_33453 ? 32'h0 : _GEN_3286; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  assign _GEN_3288 = 9'hf5 == _T_33453 ? 32'h0 : _GEN_3287; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  assign _GEN_3289 = 9'hf6 == _T_33453 ? 32'h0 : _GEN_3288; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  assign _GEN_3290 = 9'hf7 == _T_33453 ? 32'h0 : _GEN_3289; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  assign _GEN_3291 = 9'hf8 == _T_33453 ? 32'h0 : _GEN_3290; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  assign _GEN_3292 = 9'hf9 == _T_33453 ? 32'h0 : _GEN_3291; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  assign _GEN_3293 = 9'hfa == _T_33453 ? 32'h0 : _GEN_3292; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  assign _GEN_3294 = 9'hfb == _T_33453 ? 32'h0 : _GEN_3293; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  assign _GEN_3295 = 9'hfc == _T_33453 ? 32'h0 : _GEN_3294; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  assign _GEN_3296 = 9'hfd == _T_33453 ? 32'h0 : _GEN_3295; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  assign _GEN_3297 = 9'hfe == _T_33453 ? 32'h0 : _GEN_3296; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  assign _GEN_3298 = 9'hff == _T_33453 ? 32'h0 : _GEN_3297; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  assign _GEN_3299 = 9'h100 == _T_33453 ? _T_6780 : _GEN_3298; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  assign _GEN_3300 = 9'h101 == _T_33453 ? _T_6780 : _GEN_3299; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  assign _GEN_3301 = 9'h102 == _T_33453 ? _T_6780 : _GEN_3300; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  assign _GEN_3302 = 9'h103 == _T_33453 ? _T_6780 : _GEN_3301; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  assign _GEN_3303 = 9'h104 == _T_33453 ? _T_6780 : _GEN_3302; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  assign _GEN_3304 = 9'h105 == _T_33453 ? _T_6780 : _GEN_3303; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  assign _GEN_3305 = 9'h106 == _T_33453 ? _T_6780 : _GEN_3304; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  assign _GEN_3306 = 9'h107 == _T_33453 ? _T_6780 : _GEN_3305; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  assign _GEN_3307 = 9'h108 == _T_33453 ? _T_6780 : _GEN_3306; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  assign _GEN_3308 = 9'h109 == _T_33453 ? _T_6780 : _GEN_3307; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  assign _GEN_3309 = 9'h10a == _T_33453 ? _T_6780 : _GEN_3308; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  assign _GEN_3310 = 9'h10b == _T_33453 ? _T_6780 : _GEN_3309; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  assign _GEN_3311 = 9'h10c == _T_33453 ? _T_6780 : _GEN_3310; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  assign _GEN_3312 = 9'h10d == _T_33453 ? _T_6780 : _GEN_3311; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  assign _GEN_3313 = 9'h10e == _T_33453 ? _T_6780 : _GEN_3312; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  assign _GEN_3314 = 9'h10f == _T_33453 ? _T_6780 : _GEN_3313; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  assign _GEN_3315 = 9'h110 == _T_33453 ? _T_6780 : _GEN_3314; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  assign _GEN_3316 = 9'h111 == _T_33453 ? _T_6780 : _GEN_3315; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  assign _GEN_3317 = 9'h112 == _T_33453 ? _T_6780 : _GEN_3316; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  assign _GEN_3318 = 9'h113 == _T_33453 ? _T_6780 : _GEN_3317; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  assign _GEN_3319 = 9'h114 == _T_33453 ? _T_6780 : _GEN_3318; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  assign _GEN_3320 = 9'h115 == _T_33453 ? _T_6780 : _GEN_3319; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  assign _GEN_3321 = 9'h116 == _T_33453 ? _T_6780 : _GEN_3320; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  assign _GEN_3322 = 9'h117 == _T_33453 ? _T_6780 : _GEN_3321; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  assign _GEN_3323 = 9'h118 == _T_33453 ? _T_6780 : _GEN_3322; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  assign _GEN_3324 = 9'h119 == _T_33453 ? _T_6780 : _GEN_3323; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  assign _GEN_3325 = 9'h11a == _T_33453 ? _T_6780 : _GEN_3324; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  assign _GEN_3326 = 9'h11b == _T_33453 ? _T_6780 : _GEN_3325; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  assign _GEN_3327 = 9'h11c == _T_33453 ? _T_6780 : _GEN_3326; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  assign _GEN_3328 = 9'h11d == _T_33453 ? _T_6780 : _GEN_3327; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  assign _GEN_3329 = 9'h11e == _T_33453 ? _T_6780 : _GEN_3328; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  assign _GEN_3330 = 9'h11f == _T_33453 ? _T_6780 : _GEN_3329; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  assign _GEN_3331 = 9'h120 == _T_33453 ? _T_6780 : _GEN_3330; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  assign _GEN_3332 = 9'h121 == _T_33453 ? _T_6780 : _GEN_3331; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  assign _GEN_3333 = 9'h122 == _T_33453 ? _T_6780 : _GEN_3332; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  assign _GEN_3334 = 9'h123 == _T_33453 ? _T_6780 : _GEN_3333; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  assign _GEN_3335 = 9'h124 == _T_33453 ? _T_6780 : _GEN_3334; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  assign _GEN_3336 = 9'h125 == _T_33453 ? _T_6780 : _GEN_3335; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  assign _GEN_3337 = 9'h126 == _T_33453 ? _T_6780 : _GEN_3336; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  assign _GEN_3338 = 9'h127 == _T_33453 ? _T_6780 : _GEN_3337; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  assign _GEN_3339 = 9'h128 == _T_33453 ? _T_6780 : _GEN_3338; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  assign _GEN_3340 = 9'h129 == _T_33453 ? _T_6780 : _GEN_3339; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  assign _GEN_3341 = 9'h12a == _T_33453 ? _T_6780 : _GEN_3340; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  assign _GEN_3342 = 9'h12b == _T_33453 ? _T_6780 : _GEN_3341; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  assign _GEN_3343 = 9'h12c == _T_33453 ? _T_6780 : _GEN_3342; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  assign _GEN_3344 = 9'h12d == _T_33453 ? _T_6780 : _GEN_3343; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  assign _GEN_3345 = 9'h12e == _T_33453 ? _T_6780 : _GEN_3344; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  assign _GEN_3346 = 9'h12f == _T_33453 ? _T_6780 : _GEN_3345; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  assign _GEN_3347 = 9'h130 == _T_33453 ? _T_6780 : _GEN_3346; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  assign _GEN_3348 = 9'h131 == _T_33453 ? _T_6780 : _GEN_3347; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  assign _GEN_3349 = 9'h132 == _T_33453 ? _T_6780 : _GEN_3348; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  assign _GEN_3350 = 9'h133 == _T_33453 ? _T_6780 : _GEN_3349; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  assign _GEN_3351 = 9'h134 == _T_33453 ? _T_6780 : _GEN_3350; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  assign _GEN_3352 = 9'h135 == _T_33453 ? _T_6780 : _GEN_3351; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  assign _GEN_3353 = 9'h136 == _T_33453 ? _T_6780 : _GEN_3352; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  assign _GEN_3354 = 9'h137 == _T_33453 ? _T_6780 : _GEN_3353; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  assign _GEN_3355 = 9'h138 == _T_33453 ? _T_6780 : _GEN_3354; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  assign _GEN_3356 = 9'h139 == _T_33453 ? _T_6780 : _GEN_3355; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  assign _GEN_3357 = 9'h13a == _T_33453 ? _T_6780 : _GEN_3356; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  assign _GEN_3358 = 9'h13b == _T_33453 ? _T_6780 : _GEN_3357; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  assign _GEN_3359 = 9'h13c == _T_33453 ? _T_6780 : _GEN_3358; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  assign _GEN_3360 = 9'h13d == _T_33453 ? _T_6780 : _GEN_3359; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  assign _GEN_3361 = 9'h13e == _T_33453 ? _T_6780 : _GEN_3360; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  assign _GEN_3362 = 9'h13f == _T_33453 ? _T_6780 : _GEN_3361; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  assign _GEN_3363 = 9'h140 == _T_33453 ? _T_6780 : _GEN_3362; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  assign _GEN_3364 = 9'h141 == _T_33453 ? _T_6780 : _GEN_3363; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  assign _GEN_3365 = 9'h142 == _T_33453 ? _T_6780 : _GEN_3364; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  assign _GEN_3366 = 9'h143 == _T_33453 ? _T_6780 : _GEN_3365; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  assign _GEN_3367 = 9'h144 == _T_33453 ? _T_6780 : _GEN_3366; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  assign _GEN_3368 = 9'h145 == _T_33453 ? _T_6780 : _GEN_3367; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  assign _GEN_3369 = 9'h146 == _T_33453 ? _T_6780 : _GEN_3368; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  assign _GEN_3370 = 9'h147 == _T_33453 ? _T_6780 : _GEN_3369; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  assign _GEN_3371 = 9'h148 == _T_33453 ? _T_6780 : _GEN_3370; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  assign _GEN_3372 = 9'h149 == _T_33453 ? _T_6780 : _GEN_3371; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  assign _GEN_3373 = 9'h14a == _T_33453 ? _T_6780 : _GEN_3372; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  assign _GEN_3374 = 9'h14b == _T_33453 ? _T_6780 : _GEN_3373; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  assign _GEN_3375 = 9'h14c == _T_33453 ? _T_6780 : _GEN_3374; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  assign _GEN_3376 = 9'h14d == _T_33453 ? _T_6780 : _GEN_3375; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  assign _GEN_3377 = 9'h14e == _T_33453 ? _T_6780 : _GEN_3376; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  assign _GEN_3378 = 9'h14f == _T_33453 ? _T_6780 : _GEN_3377; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  assign _GEN_3379 = 9'h150 == _T_33453 ? _T_6780 : _GEN_3378; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  assign _GEN_3380 = 9'h151 == _T_33453 ? _T_6780 : _GEN_3379; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  assign _GEN_3381 = 9'h152 == _T_33453 ? _T_6780 : _GEN_3380; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  assign _GEN_3382 = 9'h153 == _T_33453 ? _T_6780 : _GEN_3381; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  assign _GEN_3383 = 9'h154 == _T_33453 ? _T_6780 : _GEN_3382; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  assign _GEN_3384 = 9'h155 == _T_33453 ? _T_6780 : _GEN_3383; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  assign _GEN_3385 = 9'h156 == _T_33453 ? _T_6780 : _GEN_3384; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  assign _GEN_3386 = 9'h157 == _T_33453 ? _T_6780 : _GEN_3385; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  assign _GEN_3387 = 9'h158 == _T_33453 ? _T_6780 : _GEN_3386; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  assign _GEN_3388 = 9'h159 == _T_33453 ? _T_6780 : _GEN_3387; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  assign _GEN_3389 = 9'h15a == _T_33453 ? _T_6780 : _GEN_3388; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  assign _GEN_3390 = 9'h15b == _T_33453 ? _T_6780 : _GEN_3389; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  assign _GEN_3391 = 9'h15c == _T_33453 ? _T_6780 : _GEN_3390; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  assign _GEN_3392 = 9'h15d == _T_33453 ? _T_6780 : _GEN_3391; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  assign _GEN_3393 = 9'h15e == _T_33453 ? _T_6780 : _GEN_3392; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  assign _GEN_3394 = 9'h15f == _T_33453 ? _T_6780 : _GEN_3393; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  assign _GEN_3395 = 9'h160 == _T_33453 ? _T_6780 : _GEN_3394; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  assign _GEN_3396 = 9'h161 == _T_33453 ? _T_6780 : _GEN_3395; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  assign _GEN_3397 = 9'h162 == _T_33453 ? _T_6780 : _GEN_3396; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  assign _GEN_3398 = 9'h163 == _T_33453 ? _T_6780 : _GEN_3397; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  assign _GEN_3399 = 9'h164 == _T_33453 ? _T_6780 : _GEN_3398; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  assign _GEN_3400 = 9'h165 == _T_33453 ? _T_6780 : _GEN_3399; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  assign _GEN_3401 = 9'h166 == _T_33453 ? _T_6780 : _GEN_3400; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  assign _GEN_3402 = 9'h167 == _T_33453 ? _T_6780 : _GEN_3401; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  assign _GEN_3403 = 9'h168 == _T_33453 ? _T_6780 : _GEN_3402; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  assign _GEN_3404 = 9'h169 == _T_33453 ? _T_6780 : _GEN_3403; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  assign _GEN_3405 = 9'h16a == _T_33453 ? _T_6780 : _GEN_3404; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  assign _GEN_3406 = 9'h16b == _T_33453 ? _T_6780 : _GEN_3405; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  assign _GEN_3407 = 9'h16c == _T_33453 ? _T_6780 : _GEN_3406; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  assign _GEN_3408 = 9'h16d == _T_33453 ? _T_6780 : _GEN_3407; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  assign _GEN_3409 = 9'h16e == _T_33453 ? _T_6780 : _GEN_3408; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  assign _GEN_3410 = 9'h16f == _T_33453 ? _T_6780 : _GEN_3409; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  assign _GEN_3411 = 9'h170 == _T_33453 ? _T_6780 : _GEN_3410; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  assign _GEN_3412 = 9'h171 == _T_33453 ? _T_6780 : _GEN_3411; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  assign _GEN_3413 = 9'h172 == _T_33453 ? _T_6780 : _GEN_3412; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  assign _GEN_3414 = 9'h173 == _T_33453 ? _T_6780 : _GEN_3413; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  assign _GEN_3415 = 9'h174 == _T_33453 ? _T_6780 : _GEN_3414; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  assign _GEN_3416 = 9'h175 == _T_33453 ? _T_6780 : _GEN_3415; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  assign _GEN_3417 = 9'h176 == _T_33453 ? _T_6780 : _GEN_3416; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  assign _GEN_3418 = 9'h177 == _T_33453 ? _T_6780 : _GEN_3417; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  assign _GEN_3419 = 9'h178 == _T_33453 ? _T_6780 : _GEN_3418; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  assign _GEN_3420 = 9'h179 == _T_33453 ? _T_6780 : _GEN_3419; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  assign _GEN_3421 = 9'h17a == _T_33453 ? _T_6780 : _GEN_3420; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  assign _GEN_3422 = 9'h17b == _T_33453 ? _T_6780 : _GEN_3421; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  assign _GEN_3423 = 9'h17c == _T_33453 ? _T_6780 : _GEN_3422; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  assign _GEN_3424 = 9'h17d == _T_33453 ? _T_6780 : _GEN_3423; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  assign _GEN_3425 = 9'h17e == _T_33453 ? _T_6780 : _GEN_3424; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  assign _GEN_3426 = 9'h17f == _T_33453 ? _T_6780 : _GEN_3425; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  assign _GEN_3427 = 9'h180 == _T_33453 ? _T_6780 : _GEN_3426; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  assign _GEN_3428 = 9'h181 == _T_33453 ? _T_6780 : _GEN_3427; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  assign _GEN_3429 = 9'h182 == _T_33453 ? _T_6780 : _GEN_3428; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  assign _GEN_3430 = 9'h183 == _T_33453 ? _T_6780 : _GEN_3429; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  assign _GEN_3431 = 9'h184 == _T_33453 ? _T_6780 : _GEN_3430; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  assign _GEN_3432 = 9'h185 == _T_33453 ? _T_6780 : _GEN_3431; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  assign _GEN_3433 = 9'h186 == _T_33453 ? _T_6780 : _GEN_3432; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  assign _GEN_3434 = 9'h187 == _T_33453 ? _T_6780 : _GEN_3433; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  assign _GEN_3435 = 9'h188 == _T_33453 ? _T_6780 : _GEN_3434; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  assign _GEN_3436 = 9'h189 == _T_33453 ? _T_6780 : _GEN_3435; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  assign _GEN_3437 = 9'h18a == _T_33453 ? _T_6780 : _GEN_3436; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  assign _GEN_3438 = 9'h18b == _T_33453 ? _T_6780 : _GEN_3437; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  assign _GEN_3439 = 9'h18c == _T_33453 ? _T_6780 : _GEN_3438; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  assign _GEN_3440 = 9'h18d == _T_33453 ? _T_6780 : _GEN_3439; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  assign _GEN_3441 = 9'h18e == _T_33453 ? _T_6780 : _GEN_3440; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  assign _GEN_3442 = 9'h18f == _T_33453 ? _T_6780 : _GEN_3441; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  assign _GEN_3443 = 9'h190 == _T_33453 ? _T_6780 : _GEN_3442; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  assign _GEN_3444 = 9'h191 == _T_33453 ? _T_6780 : _GEN_3443; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  assign _GEN_3445 = 9'h192 == _T_33453 ? _T_6780 : _GEN_3444; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  assign _GEN_3446 = 9'h193 == _T_33453 ? _T_6780 : _GEN_3445; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  assign _GEN_3447 = 9'h194 == _T_33453 ? _T_6780 : _GEN_3446; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  assign _GEN_3448 = 9'h195 == _T_33453 ? _T_6780 : _GEN_3447; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  assign _GEN_3449 = 9'h196 == _T_33453 ? _T_6780 : _GEN_3448; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  assign _GEN_3450 = 9'h197 == _T_33453 ? _T_6780 : _GEN_3449; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  assign _GEN_3451 = 9'h198 == _T_33453 ? _T_6780 : _GEN_3450; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  assign _GEN_3452 = 9'h199 == _T_33453 ? _T_6780 : _GEN_3451; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  assign _GEN_3453 = 9'h19a == _T_33453 ? _T_6780 : _GEN_3452; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  assign _GEN_3454 = 9'h19b == _T_33453 ? _T_6780 : _GEN_3453; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  assign _GEN_3455 = 9'h19c == _T_33453 ? _T_6780 : _GEN_3454; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  assign _GEN_3456 = 9'h19d == _T_33453 ? _T_6780 : _GEN_3455; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  assign _GEN_3457 = 9'h19e == _T_33453 ? _T_6780 : _GEN_3456; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  assign _GEN_3458 = 9'h19f == _T_33453 ? _T_6780 : _GEN_3457; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  assign _GEN_3459 = 9'h1a0 == _T_33453 ? _T_6780 : _GEN_3458; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  assign _GEN_3460 = 9'h1a1 == _T_33453 ? _T_6780 : _GEN_3459; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  assign _GEN_3461 = 9'h1a2 == _T_33453 ? _T_6780 : _GEN_3460; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  assign _GEN_3462 = 9'h1a3 == _T_33453 ? _T_6780 : _GEN_3461; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  assign _GEN_3463 = 9'h1a4 == _T_33453 ? _T_6780 : _GEN_3462; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  assign _GEN_3464 = 9'h1a5 == _T_33453 ? _T_6780 : _GEN_3463; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  assign _GEN_3465 = 9'h1a6 == _T_33453 ? _T_6780 : _GEN_3464; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  assign _GEN_3466 = 9'h1a7 == _T_33453 ? _T_6780 : _GEN_3465; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  assign _GEN_3467 = 9'h1a8 == _T_33453 ? _T_6780 : _GEN_3466; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  assign _GEN_3468 = 9'h1a9 == _T_33453 ? _T_6780 : _GEN_3467; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  assign _GEN_3469 = 9'h1aa == _T_33453 ? _T_6780 : _GEN_3468; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  assign _GEN_3470 = 9'h1ab == _T_33453 ? _T_6780 : _GEN_3469; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  assign _GEN_3471 = 9'h1ac == _T_33453 ? _T_6780 : _GEN_3470; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  assign _GEN_3472 = 9'h1ad == _T_33453 ? _T_6780 : _GEN_3471; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  assign _GEN_3473 = 9'h1ae == _T_33453 ? _T_6780 : _GEN_3472; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  assign _GEN_3474 = 9'h1af == _T_33453 ? _T_6780 : _GEN_3473; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  assign _GEN_3475 = 9'h1b0 == _T_33453 ? _T_6780 : _GEN_3474; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  assign _GEN_3476 = 9'h1b1 == _T_33453 ? _T_6780 : _GEN_3475; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  assign _GEN_3477 = 9'h1b2 == _T_33453 ? _T_6780 : _GEN_3476; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  assign _GEN_3478 = 9'h1b3 == _T_33453 ? _T_6780 : _GEN_3477; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  assign _GEN_3479 = 9'h1b4 == _T_33453 ? _T_6780 : _GEN_3478; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  assign _GEN_3480 = 9'h1b5 == _T_33453 ? _T_6780 : _GEN_3479; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  assign _GEN_3481 = 9'h1b6 == _T_33453 ? _T_6780 : _GEN_3480; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  assign _GEN_3482 = 9'h1b7 == _T_33453 ? _T_6780 : _GEN_3481; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  assign _GEN_3483 = 9'h1b8 == _T_33453 ? _T_6780 : _GEN_3482; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  assign _GEN_3484 = 9'h1b9 == _T_33453 ? _T_6780 : _GEN_3483; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  assign _GEN_3485 = 9'h1ba == _T_33453 ? _T_6780 : _GEN_3484; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  assign _GEN_3486 = 9'h1bb == _T_33453 ? _T_6780 : _GEN_3485; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  assign _GEN_3487 = 9'h1bc == _T_33453 ? _T_6780 : _GEN_3486; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  assign _GEN_3488 = 9'h1bd == _T_33453 ? _T_6780 : _GEN_3487; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  assign _GEN_3489 = 9'h1be == _T_33453 ? _T_6780 : _GEN_3488; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  assign _GEN_3490 = 9'h1bf == _T_33453 ? _T_6780 : _GEN_3489; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  assign _GEN_3491 = 9'h1c0 == _T_33453 ? _T_6780 : _GEN_3490; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  assign _GEN_3492 = 9'h1c1 == _T_33453 ? _T_6780 : _GEN_3491; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  assign _GEN_3493 = 9'h1c2 == _T_33453 ? _T_6780 : _GEN_3492; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  assign _GEN_3494 = 9'h1c3 == _T_33453 ? _T_6780 : _GEN_3493; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  assign _GEN_3495 = 9'h1c4 == _T_33453 ? _T_6780 : _GEN_3494; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  assign _GEN_3496 = 9'h1c5 == _T_33453 ? _T_6780 : _GEN_3495; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  assign _GEN_3497 = 9'h1c6 == _T_33453 ? _T_6780 : _GEN_3496; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  assign _GEN_3498 = 9'h1c7 == _T_33453 ? _T_6780 : _GEN_3497; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  assign _GEN_3499 = 9'h1c8 == _T_33453 ? _T_6780 : _GEN_3498; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  assign _GEN_3500 = 9'h1c9 == _T_33453 ? _T_6780 : _GEN_3499; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  assign _GEN_3501 = 9'h1ca == _T_33453 ? _T_6780 : _GEN_3500; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  assign _GEN_3502 = 9'h1cb == _T_33453 ? _T_6780 : _GEN_3501; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  assign _GEN_3503 = 9'h1cc == _T_33453 ? _T_6780 : _GEN_3502; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  assign _GEN_3504 = 9'h1cd == _T_33453 ? _T_6780 : _GEN_3503; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  assign _GEN_3505 = 9'h1ce == _T_33453 ? _T_6780 : _GEN_3504; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  assign _GEN_3506 = 9'h1cf == _T_33453 ? _T_6780 : _GEN_3505; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  assign _GEN_3507 = 9'h1d0 == _T_33453 ? _T_6780 : _GEN_3506; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  assign _GEN_3508 = 9'h1d1 == _T_33453 ? _T_6780 : _GEN_3507; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  assign _GEN_3509 = 9'h1d2 == _T_33453 ? _T_6780 : _GEN_3508; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  assign _GEN_3510 = 9'h1d3 == _T_33453 ? _T_6780 : _GEN_3509; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  assign _GEN_3511 = 9'h1d4 == _T_33453 ? _T_6780 : _GEN_3510; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  assign _GEN_3512 = 9'h1d5 == _T_33453 ? _T_6780 : _GEN_3511; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  assign _GEN_3513 = 9'h1d6 == _T_33453 ? _T_6780 : _GEN_3512; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  assign _GEN_3514 = 9'h1d7 == _T_33453 ? _T_6780 : _GEN_3513; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  assign _GEN_3515 = 9'h1d8 == _T_33453 ? _T_6780 : _GEN_3514; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  assign _GEN_3516 = 9'h1d9 == _T_33453 ? _T_6780 : _GEN_3515; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  assign _GEN_3517 = 9'h1da == _T_33453 ? _T_6780 : _GEN_3516; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  assign _GEN_3518 = 9'h1db == _T_33453 ? _T_6780 : _GEN_3517; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  assign _GEN_3519 = 9'h1dc == _T_33453 ? _T_6780 : _GEN_3518; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  assign _GEN_3520 = 9'h1dd == _T_33453 ? _T_6780 : _GEN_3519; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  assign _GEN_3521 = 9'h1de == _T_33453 ? _T_6780 : _GEN_3520; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  assign _GEN_3522 = 9'h1df == _T_33453 ? _T_6780 : _GEN_3521; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  assign _GEN_3523 = 9'h1e0 == _T_33453 ? _T_6780 : _GEN_3522; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  assign _GEN_3524 = 9'h1e1 == _T_33453 ? _T_6780 : _GEN_3523; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  assign _GEN_3525 = 9'h1e2 == _T_33453 ? _T_6780 : _GEN_3524; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  assign _GEN_3526 = 9'h1e3 == _T_33453 ? _T_6780 : _GEN_3525; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  assign _GEN_3527 = 9'h1e4 == _T_33453 ? _T_6780 : _GEN_3526; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  assign _GEN_3528 = 9'h1e5 == _T_33453 ? _T_6780 : _GEN_3527; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  assign _GEN_3529 = 9'h1e6 == _T_33453 ? _T_6780 : _GEN_3528; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  assign _GEN_3530 = 9'h1e7 == _T_33453 ? _T_6780 : _GEN_3529; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  assign _GEN_3531 = 9'h1e8 == _T_33453 ? _T_6780 : _GEN_3530; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  assign _GEN_3532 = 9'h1e9 == _T_33453 ? _T_6780 : _GEN_3531; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  assign _GEN_3533 = 9'h1ea == _T_33453 ? _T_6780 : _GEN_3532; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  assign _GEN_3534 = 9'h1eb == _T_33453 ? _T_6780 : _GEN_3533; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  assign _GEN_3535 = 9'h1ec == _T_33453 ? _T_6780 : _GEN_3534; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  assign _GEN_3536 = 9'h1ed == _T_33453 ? _T_6780 : _GEN_3535; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  assign _GEN_3537 = 9'h1ee == _T_33453 ? _T_6780 : _GEN_3536; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  assign _GEN_3538 = 9'h1ef == _T_33453 ? _T_6780 : _GEN_3537; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  assign _GEN_3539 = 9'h1f0 == _T_33453 ? _T_6780 : _GEN_3538; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  assign _GEN_3540 = 9'h1f1 == _T_33453 ? _T_6780 : _GEN_3539; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  assign _GEN_3541 = 9'h1f2 == _T_33453 ? _T_6780 : _GEN_3540; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  assign _GEN_3542 = 9'h1f3 == _T_33453 ? _T_6780 : _GEN_3541; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  assign _GEN_3543 = 9'h1f4 == _T_33453 ? _T_6780 : _GEN_3542; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  assign _GEN_3544 = 9'h1f5 == _T_33453 ? _T_6780 : _GEN_3543; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  assign _GEN_3545 = 9'h1f6 == _T_33453 ? _T_6780 : _GEN_3544; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  assign _GEN_3546 = 9'h1f7 == _T_33453 ? _T_6780 : _GEN_3545; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  assign _GEN_3547 = 9'h1f8 == _T_33453 ? _T_6780 : _GEN_3546; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  assign _GEN_3548 = 9'h1f9 == _T_33453 ? _T_6780 : _GEN_3547; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  assign _GEN_3549 = 9'h1fa == _T_33453 ? _T_6780 : _GEN_3548; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  assign _GEN_3550 = 9'h1fb == _T_33453 ? _T_6780 : _GEN_3549; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  assign _GEN_3551 = 9'h1fc == _T_33453 ? _T_6780 : _GEN_3550; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  assign _GEN_3552 = 9'h1fd == _T_33453 ? _T_6780 : _GEN_3551; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  assign _GEN_3553 = 9'h1fe == _T_33453 ? _T_6780 : _GEN_3552; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  assign _GEN_3554 = 9'h1ff == _T_33453 ? _T_6780 : _GEN_3553; // @[MuxLiteral.scala 48:10:freechips.rocketchip.system.DefaultRV32Config.fir@168555.4]
  assign _T_44820 = ~goReg; // @[Debug.scala 1649:18:freechips.rocketchip.system.DefaultRV32Config.fir@168764.10]
  assign _T_44821 = _T_44820 & hartHaltedWrEn; // @[Debug.scala 1649:30:freechips.rocketchip.system.DefaultRV32Config.fir@168765.10]
  assign _T_44828 = ctrlStateReg == 2'h3; // @[Debug.scala 1657:30:freechips.rocketchip.system.DefaultRV32Config.fir@168785.10]
  assign _T_44831 = ~reset; // @[Debug.scala 1658:13:freechips.rocketchip.system.DefaultRV32Config.fir@168789.12]
  assign _T_44837 = ~hartExceptionWrEn; // @[Debug.scala 1671:30:freechips.rocketchip.system.DefaultRV32Config.fir@168810.4]
  assign _T_44838 = _T_13 | _T_44837; // @[Debug.scala 1671:27:freechips.rocketchip.system.DefaultRV32Config.fir@168811.4]
  assign _T_44840 = _T_44838 | _T_44819; // @[Debug.scala 1671:49:freechips.rocketchip.system.DefaultRV32Config.fir@168813.4]
  assign _T_44842 = _T_44840 | reset; // @[Debug.scala 1671:12:freechips.rocketchip.system.DefaultRV32Config.fir@168815.4]
  assign _T_44843 = ~_T_44842; // @[Debug.scala 1671:12:freechips.rocketchip.system.DefaultRV32Config.fir@168816.4]
  assign auto_tl_in_a_ready = auto_tl_in_d_ready; // @[LazyModule.scala 303:16:freechips.rocketchip.system.DefaultRV32Config.fir@108970.4]
  assign auto_tl_in_d_valid = auto_tl_in_a_valid; // @[LazyModule.scala 303:16:freechips.rocketchip.system.DefaultRV32Config.fir@108970.4]
  assign auto_tl_in_d_bits_opcode = {{2'd0}, _T_6050}; // @[LazyModule.scala 303:16:freechips.rocketchip.system.DefaultRV32Config.fir@108970.4]
  assign auto_tl_in_d_bits_size = auto_tl_in_a_bits_size; // @[LazyModule.scala 303:16:freechips.rocketchip.system.DefaultRV32Config.fir@108970.4]
  assign auto_tl_in_d_bits_source = auto_tl_in_a_bits_source; // @[LazyModule.scala 303:16:freechips.rocketchip.system.DefaultRV32Config.fir@108970.4]
  assign auto_tl_in_d_bits_data = _GEN_3042 ? _GEN_3554 : 32'h0; // @[LazyModule.scala 303:16:freechips.rocketchip.system.DefaultRV32Config.fir@108970.4]
  assign auto_dmi_in_a_ready = auto_dmi_in_d_ready; // @[LazyModule.scala 303:16:freechips.rocketchip.system.DefaultRV32Config.fir@108969.4]
  assign auto_dmi_in_d_valid = auto_dmi_in_a_valid; // @[LazyModule.scala 303:16:freechips.rocketchip.system.DefaultRV32Config.fir@108969.4]
  assign auto_dmi_in_d_bits_opcode = {{2'd0}, _T_380}; // @[LazyModule.scala 303:16:freechips.rocketchip.system.DefaultRV32Config.fir@108969.4]
  assign auto_dmi_in_d_bits_size = auto_dmi_in_a_bits_size; // @[LazyModule.scala 303:16:freechips.rocketchip.system.DefaultRV32Config.fir@108969.4]
  assign auto_dmi_in_d_bits_source = auto_dmi_in_a_bits_source; // @[LazyModule.scala 303:16:freechips.rocketchip.system.DefaultRV32Config.fir@108969.4]
  assign auto_dmi_in_d_bits_data = _GEN_305 ? _GEN_337 : 32'h0; // @[LazyModule.scala 303:16:freechips.rocketchip.system.DefaultRV32Config.fir@108969.4]
  assign io_innerCtrl_ready = 1'h1; // @[Debug.scala 814:24:freechips.rocketchip.system.DefaultRV32Config.fir@109277.4]
  assign io_hgDebugInt_0 = hrDebugInt_0; // @[Debug.scala 1036:19:freechips.rocketchip.system.DefaultRV32Config.fir@109480.4]
  assign TLMonitor_clock = clock; // @[:freechips.rocketchip.system.DefaultRV32Config.fir@108920.4]
  assign TLMonitor_reset = reset; // @[:freechips.rocketchip.system.DefaultRV32Config.fir@108921.4]
  assign TLMonitor_io_in_a_ready = auto_dmi_in_d_ready; // @[Nodes.scala 26:19:freechips.rocketchip.system.DefaultRV32Config.fir@108941.4]
  assign TLMonitor_io_in_a_valid = auto_dmi_in_a_valid; // @[Nodes.scala 26:19:freechips.rocketchip.system.DefaultRV32Config.fir@108940.4]
  assign TLMonitor_io_in_a_bits_opcode = auto_dmi_in_a_bits_opcode; // @[Nodes.scala 26:19:freechips.rocketchip.system.DefaultRV32Config.fir@108939.4]
  assign TLMonitor_io_in_a_bits_param = auto_dmi_in_a_bits_param; // @[Nodes.scala 26:19:freechips.rocketchip.system.DefaultRV32Config.fir@108938.4]
  assign TLMonitor_io_in_a_bits_size = auto_dmi_in_a_bits_size; // @[Nodes.scala 26:19:freechips.rocketchip.system.DefaultRV32Config.fir@108937.4]
  assign TLMonitor_io_in_a_bits_source = auto_dmi_in_a_bits_source; // @[Nodes.scala 26:19:freechips.rocketchip.system.DefaultRV32Config.fir@108936.4]
  assign TLMonitor_io_in_a_bits_address = auto_dmi_in_a_bits_address; // @[Nodes.scala 26:19:freechips.rocketchip.system.DefaultRV32Config.fir@108935.4]
  assign TLMonitor_io_in_a_bits_mask = auto_dmi_in_a_bits_mask; // @[Nodes.scala 26:19:freechips.rocketchip.system.DefaultRV32Config.fir@108934.4]
  assign TLMonitor_io_in_a_bits_corrupt = auto_dmi_in_a_bits_corrupt; // @[Nodes.scala 26:19:freechips.rocketchip.system.DefaultRV32Config.fir@108932.4]
  assign TLMonitor_io_in_d_ready = auto_dmi_in_d_ready; // @[Nodes.scala 26:19:freechips.rocketchip.system.DefaultRV32Config.fir@108931.4]
  assign TLMonitor_io_in_d_valid = auto_dmi_in_a_valid; // @[Nodes.scala 26:19:freechips.rocketchip.system.DefaultRV32Config.fir@108930.4]
  assign TLMonitor_io_in_d_bits_opcode = {{2'd0}, _T_380}; // @[Nodes.scala 26:19:freechips.rocketchip.system.DefaultRV32Config.fir@108929.4]
  assign TLMonitor_io_in_d_bits_size = auto_dmi_in_a_bits_size; // @[Nodes.scala 26:19:freechips.rocketchip.system.DefaultRV32Config.fir@108927.4]
  assign TLMonitor_io_in_d_bits_source = auto_dmi_in_a_bits_source; // @[Nodes.scala 26:19:freechips.rocketchip.system.DefaultRV32Config.fir@108926.4]
  assign TLMonitor_1_clock = clock; // @[:freechips.rocketchip.system.DefaultRV32Config.fir@108945.4]
  assign TLMonitor_1_reset = reset; // @[:freechips.rocketchip.system.DefaultRV32Config.fir@108946.4]
  assign TLMonitor_1_io_in_a_ready = auto_tl_in_d_ready; // @[Nodes.scala 26:19:freechips.rocketchip.system.DefaultRV32Config.fir@108966.4]
  assign TLMonitor_1_io_in_a_valid = auto_tl_in_a_valid; // @[Nodes.scala 26:19:freechips.rocketchip.system.DefaultRV32Config.fir@108965.4]
  assign TLMonitor_1_io_in_a_bits_opcode = auto_tl_in_a_bits_opcode; // @[Nodes.scala 26:19:freechips.rocketchip.system.DefaultRV32Config.fir@108964.4]
  assign TLMonitor_1_io_in_a_bits_param = auto_tl_in_a_bits_param; // @[Nodes.scala 26:19:freechips.rocketchip.system.DefaultRV32Config.fir@108963.4]
  assign TLMonitor_1_io_in_a_bits_size = auto_tl_in_a_bits_size; // @[Nodes.scala 26:19:freechips.rocketchip.system.DefaultRV32Config.fir@108962.4]
  assign TLMonitor_1_io_in_a_bits_source = auto_tl_in_a_bits_source; // @[Nodes.scala 26:19:freechips.rocketchip.system.DefaultRV32Config.fir@108961.4]
  assign TLMonitor_1_io_in_a_bits_address = auto_tl_in_a_bits_address; // @[Nodes.scala 26:19:freechips.rocketchip.system.DefaultRV32Config.fir@108960.4]
  assign TLMonitor_1_io_in_a_bits_mask = auto_tl_in_a_bits_mask; // @[Nodes.scala 26:19:freechips.rocketchip.system.DefaultRV32Config.fir@108959.4]
  assign TLMonitor_1_io_in_a_bits_corrupt = auto_tl_in_a_bits_corrupt; // @[Nodes.scala 26:19:freechips.rocketchip.system.DefaultRV32Config.fir@108957.4]
  assign TLMonitor_1_io_in_d_ready = auto_tl_in_d_ready; // @[Nodes.scala 26:19:freechips.rocketchip.system.DefaultRV32Config.fir@108956.4]
  assign TLMonitor_1_io_in_d_valid = auto_tl_in_a_valid; // @[Nodes.scala 26:19:freechips.rocketchip.system.DefaultRV32Config.fir@108955.4]
  assign TLMonitor_1_io_in_d_bits_opcode = {{2'd0}, _T_6050}; // @[Nodes.scala 26:19:freechips.rocketchip.system.DefaultRV32Config.fir@108954.4]
  assign TLMonitor_1_io_in_d_bits_size = auto_tl_in_a_bits_size; // @[Nodes.scala 26:19:freechips.rocketchip.system.DefaultRV32Config.fir@108952.4]
  assign TLMonitor_1_io_in_d_bits_source = auto_tl_in_a_bits_source; // @[Nodes.scala 26:19:freechips.rocketchip.system.DefaultRV32Config.fir@108951.4]
  assign debug_hartReset_0_clock = clock; // @[:freechips.rocketchip.system.DefaultRV32Config.fir@109293.4]
  assign debug_hartReset_0_reset = reset; // @[:freechips.rocketchip.system.DefaultRV32Config.fir@109294.4]
  assign debug_hartReset_0_io_d = io_hartIsInReset_0; // @[ShiftReg.scala 47:16:freechips.rocketchip.system.DefaultRV32Config.fir@109295.4]
  assign _GEN_3883 = ~_T_13; // @[Debug.scala 1389:15:freechips.rocketchip.system.DefaultRV32Config.fir@115473.12]
  assign _GEN_3884 = ~goAbstract; // @[Debug.scala 1389:15:freechips.rocketchip.system.DefaultRV32Config.fir@115473.12]
  assign _GEN_3885 = _GEN_3883 & _GEN_3884; // @[Debug.scala 1389:15:freechips.rocketchip.system.DefaultRV32Config.fir@115473.12]
  assign _GEN_3886 = _GEN_3885 & hartGoingWrEn; // @[Debug.scala 1389:15:freechips.rocketchip.system.DefaultRV32Config.fir@115473.12]
  assign _GEN_3892 = ~_T_44818; // @[Debug.scala 1653:15:freechips.rocketchip.system.DefaultRV32Config.fir@168777.14]
  assign _GEN_3893 = _T_44785 & _GEN_3892; // @[Debug.scala 1653:15:freechips.rocketchip.system.DefaultRV32Config.fir@168777.14]
  assign _GEN_3894 = _GEN_3893 & _T_44819; // @[Debug.scala 1653:15:freechips.rocketchip.system.DefaultRV32Config.fir@168777.14]
  assign _GEN_3895 = _GEN_3894 & hartExceptionWrEn; // @[Debug.scala 1653:15:freechips.rocketchip.system.DefaultRV32Config.fir@168777.14]
  assign _GEN_3904 = ~_T_44819; // @[Debug.scala 1658:13:freechips.rocketchip.system.DefaultRV32Config.fir@168791.14]
  assign _GEN_3905 = _GEN_3893 & _GEN_3904; // @[Debug.scala 1658:13:freechips.rocketchip.system.DefaultRV32Config.fir@168791.14]
  assign _GEN_3906 = _GEN_3905 & _T_44828; // @[Debug.scala 1658:13:freechips.rocketchip.system.DefaultRV32Config.fir@168791.14]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  haltedBitRegs_0 = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  resumeReqRegs_0 = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  haveResetBitRegs_0 = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  hrmaskReg_0 = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  hrDebugInt_0 = _RAND_4[0:0];
  _RAND_5 = {1{`RANDOM}};
  ABSTRACTCSReg_cmderr = _RAND_5[2:0];
  _RAND_6 = {1{`RANDOM}};
  ctrlStateReg = _RAND_6[1:0];
  _RAND_7 = {1{`RANDOM}};
  COMMANDRdData_cmdtype = _RAND_7[7:0];
  _RAND_8 = {1{`RANDOM}};
  COMMANDRdData_control = _RAND_8[23:0];
  _RAND_9 = {1{`RANDOM}};
  ABSTRACTAUTOReg_autoexecdata = _RAND_9[11:0];
  _RAND_10 = {1{`RANDOM}};
  ABSTRACTAUTOReg_autoexecprogbuf = _RAND_10[15:0];
  _RAND_11 = {1{`RANDOM}};
  abstractDataMem_0 = _RAND_11[7:0];
  _RAND_12 = {1{`RANDOM}};
  abstractDataMem_1 = _RAND_12[7:0];
  _RAND_13 = {1{`RANDOM}};
  abstractDataMem_2 = _RAND_13[7:0];
  _RAND_14 = {1{`RANDOM}};
  abstractDataMem_3 = _RAND_14[7:0];
  _RAND_15 = {1{`RANDOM}};
  programBufferMem_0 = _RAND_15[7:0];
  _RAND_16 = {1{`RANDOM}};
  programBufferMem_1 = _RAND_16[7:0];
  _RAND_17 = {1{`RANDOM}};
  programBufferMem_2 = _RAND_17[7:0];
  _RAND_18 = {1{`RANDOM}};
  programBufferMem_3 = _RAND_18[7:0];
  _RAND_19 = {1{`RANDOM}};
  programBufferMem_4 = _RAND_19[7:0];
  _RAND_20 = {1{`RANDOM}};
  programBufferMem_5 = _RAND_20[7:0];
  _RAND_21 = {1{`RANDOM}};
  programBufferMem_6 = _RAND_21[7:0];
  _RAND_22 = {1{`RANDOM}};
  programBufferMem_7 = _RAND_22[7:0];
  _RAND_23 = {1{`RANDOM}};
  programBufferMem_8 = _RAND_23[7:0];
  _RAND_24 = {1{`RANDOM}};
  programBufferMem_9 = _RAND_24[7:0];
  _RAND_25 = {1{`RANDOM}};
  programBufferMem_10 = _RAND_25[7:0];
  _RAND_26 = {1{`RANDOM}};
  programBufferMem_11 = _RAND_26[7:0];
  _RAND_27 = {1{`RANDOM}};
  programBufferMem_12 = _RAND_27[7:0];
  _RAND_28 = {1{`RANDOM}};
  programBufferMem_13 = _RAND_28[7:0];
  _RAND_29 = {1{`RANDOM}};
  programBufferMem_14 = _RAND_29[7:0];
  _RAND_30 = {1{`RANDOM}};
  programBufferMem_15 = _RAND_30[7:0];
  _RAND_31 = {1{`RANDOM}};
  programBufferMem_16 = _RAND_31[7:0];
  _RAND_32 = {1{`RANDOM}};
  programBufferMem_17 = _RAND_32[7:0];
  _RAND_33 = {1{`RANDOM}};
  programBufferMem_18 = _RAND_33[7:0];
  _RAND_34 = {1{`RANDOM}};
  programBufferMem_19 = _RAND_34[7:0];
  _RAND_35 = {1{`RANDOM}};
  programBufferMem_20 = _RAND_35[7:0];
  _RAND_36 = {1{`RANDOM}};
  programBufferMem_21 = _RAND_36[7:0];
  _RAND_37 = {1{`RANDOM}};
  programBufferMem_22 = _RAND_37[7:0];
  _RAND_38 = {1{`RANDOM}};
  programBufferMem_23 = _RAND_38[7:0];
  _RAND_39 = {1{`RANDOM}};
  programBufferMem_24 = _RAND_39[7:0];
  _RAND_40 = {1{`RANDOM}};
  programBufferMem_25 = _RAND_40[7:0];
  _RAND_41 = {1{`RANDOM}};
  programBufferMem_26 = _RAND_41[7:0];
  _RAND_42 = {1{`RANDOM}};
  programBufferMem_27 = _RAND_42[7:0];
  _RAND_43 = {1{`RANDOM}};
  programBufferMem_28 = _RAND_43[7:0];
  _RAND_44 = {1{`RANDOM}};
  programBufferMem_29 = _RAND_44[7:0];
  _RAND_45 = {1{`RANDOM}};
  programBufferMem_30 = _RAND_45[7:0];
  _RAND_46 = {1{`RANDOM}};
  programBufferMem_31 = _RAND_46[7:0];
  _RAND_47 = {1{`RANDOM}};
  programBufferMem_32 = _RAND_47[7:0];
  _RAND_48 = {1{`RANDOM}};
  programBufferMem_33 = _RAND_48[7:0];
  _RAND_49 = {1{`RANDOM}};
  programBufferMem_34 = _RAND_49[7:0];
  _RAND_50 = {1{`RANDOM}};
  programBufferMem_35 = _RAND_50[7:0];
  _RAND_51 = {1{`RANDOM}};
  programBufferMem_36 = _RAND_51[7:0];
  _RAND_52 = {1{`RANDOM}};
  programBufferMem_37 = _RAND_52[7:0];
  _RAND_53 = {1{`RANDOM}};
  programBufferMem_38 = _RAND_53[7:0];
  _RAND_54 = {1{`RANDOM}};
  programBufferMem_39 = _RAND_54[7:0];
  _RAND_55 = {1{`RANDOM}};
  programBufferMem_40 = _RAND_55[7:0];
  _RAND_56 = {1{`RANDOM}};
  programBufferMem_41 = _RAND_56[7:0];
  _RAND_57 = {1{`RANDOM}};
  programBufferMem_42 = _RAND_57[7:0];
  _RAND_58 = {1{`RANDOM}};
  programBufferMem_43 = _RAND_58[7:0];
  _RAND_59 = {1{`RANDOM}};
  programBufferMem_44 = _RAND_59[7:0];
  _RAND_60 = {1{`RANDOM}};
  programBufferMem_45 = _RAND_60[7:0];
  _RAND_61 = {1{`RANDOM}};
  programBufferMem_46 = _RAND_61[7:0];
  _RAND_62 = {1{`RANDOM}};
  programBufferMem_47 = _RAND_62[7:0];
  _RAND_63 = {1{`RANDOM}};
  programBufferMem_48 = _RAND_63[7:0];
  _RAND_64 = {1{`RANDOM}};
  programBufferMem_49 = _RAND_64[7:0];
  _RAND_65 = {1{`RANDOM}};
  programBufferMem_50 = _RAND_65[7:0];
  _RAND_66 = {1{`RANDOM}};
  programBufferMem_51 = _RAND_66[7:0];
  _RAND_67 = {1{`RANDOM}};
  programBufferMem_52 = _RAND_67[7:0];
  _RAND_68 = {1{`RANDOM}};
  programBufferMem_53 = _RAND_68[7:0];
  _RAND_69 = {1{`RANDOM}};
  programBufferMem_54 = _RAND_69[7:0];
  _RAND_70 = {1{`RANDOM}};
  programBufferMem_55 = _RAND_70[7:0];
  _RAND_71 = {1{`RANDOM}};
  programBufferMem_56 = _RAND_71[7:0];
  _RAND_72 = {1{`RANDOM}};
  programBufferMem_57 = _RAND_72[7:0];
  _RAND_73 = {1{`RANDOM}};
  programBufferMem_58 = _RAND_73[7:0];
  _RAND_74 = {1{`RANDOM}};
  programBufferMem_59 = _RAND_74[7:0];
  _RAND_75 = {1{`RANDOM}};
  programBufferMem_60 = _RAND_75[7:0];
  _RAND_76 = {1{`RANDOM}};
  programBufferMem_61 = _RAND_76[7:0];
  _RAND_77 = {1{`RANDOM}};
  programBufferMem_62 = _RAND_77[7:0];
  _RAND_78 = {1{`RANDOM}};
  programBufferMem_63 = _RAND_78[7:0];
  _RAND_79 = {1{`RANDOM}};
  goReg = _RAND_79[0:0];
  _RAND_80 = {1{`RANDOM}};
  abstractGeneratedMem_0 = _RAND_80[31:0];
  _RAND_81 = {1{`RANDOM}};
  abstractGeneratedMem_1 = _RAND_81[31:0];
`endif // RANDOMIZE_REG_INIT
  if (reset) begin
    hrDebugInt_0 = 1'h0;
  end
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (_T_13) begin
      haltedBitRegs_0 <= 1'h0;
    end else if (hartIsInResetSync_0) begin
      haltedBitRegs_0 <= 1'h0;
    end else begin
      haltedBitRegs_0 <= _GEN_69;
    end
    if (_T_13) begin
      resumeReqRegs_0 <= 1'h0;
    end else begin
      resumeReqRegs_0 <= _GEN_74;
    end
    if (_T_13) begin
      haveResetBitRegs_0 <= 1'h0;
    end else begin
      haveResetBitRegs_0 <= _GEN_35;
    end
    if (reset) begin
      hrmaskReg_0 <= 1'h0;
    end else if (_T_13) begin
      hrmaskReg_0 <= 1'h0;
    end else if (_T_16) begin
      hrmaskReg_0 <= io_innerCtrl_bits_hrmask_0;
    end
    if (_T_13) begin
      ABSTRACTCSReg_cmderr <= 3'h0;
    end else if (errorBusy) begin
      ABSTRACTCSReg_cmderr <= 3'h1;
    end else if (errorException) begin
      ABSTRACTCSReg_cmderr <= 3'h3;
    end else if (errorUnsupported) begin
      ABSTRACTCSReg_cmderr <= 3'h2;
    end else if (errorHaltResume) begin
      ABSTRACTCSReg_cmderr <= 3'h4;
    end else if (ABSTRACTCSWrEn) begin
      ABSTRACTCSReg_cmderr <= _T_84;
    end
    if (_T_13) begin
      ctrlStateReg <= 2'h0;
    end else if (ABSTRACTCSWrEnLegal) begin
      if (_T_44816) begin
        ctrlStateReg <= 2'h1;
      end
    end else if (_T_44818) begin
      if (commandRegIsUnsupported) begin
        ctrlStateReg <= 2'h0;
      end else if (commandRegBadHaltResume) begin
        ctrlStateReg <= 2'h0;
      end else begin
        ctrlStateReg <= 2'h2;
      end
    end else if (_T_44819) begin
      if (hartExceptionWrEn) begin
        ctrlStateReg <= 2'h0;
      end else if (_T_44821) begin
        ctrlStateReg <= 2'h0;
      end
    end
    if (_T_13) begin
      COMMANDRdData_cmdtype <= 8'h0;
    end else if (COMMANDWrEn) begin
      COMMANDRdData_cmdtype <= COMMANDWrData_cmdtype;
    end
    if (_T_13) begin
      COMMANDRdData_control <= 24'h0;
    end else if (COMMANDWrEn) begin
      COMMANDRdData_control <= COMMANDWrData_control;
    end
    if (_T_13) begin
      ABSTRACTAUTOReg_autoexecdata <= 12'h0;
    end else if (_T_93) begin
      ABSTRACTAUTOReg_autoexecdata <= _T_94;
    end
    if (_T_13) begin
      ABSTRACTAUTOReg_autoexecprogbuf <= 16'h0;
    end else if (_T_91) begin
      ABSTRACTAUTOReg_autoexecprogbuf <= ABSTRACTAUTOWrData_autoexecprogbuf;
    end
    if (_T_13) begin
      abstractDataMem_0 <= 8'h0;
    end else if (_T_15806) begin
      abstractDataMem_0 <= auto_tl_in_a_bits_data[7:0];
    end else if (_T_3749) begin
      if (dmiAbstractDataWrEnMaybe_0) begin
        abstractDataMem_0 <= auto_dmi_in_a_bits_data[7:0];
      end
    end
    if (_T_13) begin
      abstractDataMem_1 <= 8'h0;
    end else if (_T_15829) begin
      abstractDataMem_1 <= auto_tl_in_a_bits_data[15:8];
    end else if (_T_3751) begin
      if (dmiAbstractDataWrEnMaybe_1) begin
        abstractDataMem_1 <= auto_dmi_in_a_bits_data[15:8];
      end
    end
    if (_T_13) begin
      abstractDataMem_2 <= 8'h0;
    end else if (_T_15854) begin
      abstractDataMem_2 <= auto_tl_in_a_bits_data[23:16];
    end else if (_T_3753) begin
      if (dmiAbstractDataWrEnMaybe_2) begin
        abstractDataMem_2 <= auto_dmi_in_a_bits_data[23:16];
      end
    end
    if (_T_13) begin
      abstractDataMem_3 <= 8'h0;
    end else if (_T_15879) begin
      abstractDataMem_3 <= auto_tl_in_a_bits_data[31:24];
    end else if (_T_3755) begin
      if (dmiAbstractDataWrEnMaybe_3) begin
        abstractDataMem_3 <= auto_dmi_in_a_bits_data[31:24];
      end
    end
    if (_T_13) begin
      programBufferMem_0 <= 8'h0;
    end else if (_T_21791) begin
      programBufferMem_0 <= auto_tl_in_a_bits_data[7:0];
    end else if (_T_3757) begin
      if (dmiProgramBufferWrEnMaybe_0) begin
        programBufferMem_0 <= auto_dmi_in_a_bits_data[7:0];
      end
    end
    if (_T_13) begin
      programBufferMem_1 <= 8'h0;
    end else if (_T_21814) begin
      programBufferMem_1 <= auto_tl_in_a_bits_data[15:8];
    end else if (_T_3759) begin
      if (dmiProgramBufferWrEnMaybe_1) begin
        programBufferMem_1 <= auto_dmi_in_a_bits_data[15:8];
      end
    end
    if (_T_13) begin
      programBufferMem_2 <= 8'h0;
    end else if (_T_21839) begin
      programBufferMem_2 <= auto_tl_in_a_bits_data[23:16];
    end else if (_T_3761) begin
      if (dmiProgramBufferWrEnMaybe_2) begin
        programBufferMem_2 <= auto_dmi_in_a_bits_data[23:16];
      end
    end
    if (_T_13) begin
      programBufferMem_3 <= 8'h0;
    end else if (_T_21864) begin
      programBufferMem_3 <= auto_tl_in_a_bits_data[31:24];
    end else if (_T_3763) begin
      if (dmiProgramBufferWrEnMaybe_3) begin
        programBufferMem_3 <= auto_dmi_in_a_bits_data[31:24];
      end
    end
    if (_T_13) begin
      programBufferMem_4 <= 8'h0;
    end else if (_T_24446) begin
      programBufferMem_4 <= auto_tl_in_a_bits_data[7:0];
    end else if (_T_3765) begin
      if (dmiProgramBufferWrEnMaybe_4) begin
        programBufferMem_4 <= auto_dmi_in_a_bits_data[7:0];
      end
    end
    if (_T_13) begin
      programBufferMem_5 <= 8'h0;
    end else if (_T_24469) begin
      programBufferMem_5 <= auto_tl_in_a_bits_data[15:8];
    end else if (_T_3767) begin
      if (dmiProgramBufferWrEnMaybe_5) begin
        programBufferMem_5 <= auto_dmi_in_a_bits_data[15:8];
      end
    end
    if (_T_13) begin
      programBufferMem_6 <= 8'h0;
    end else if (_T_24494) begin
      programBufferMem_6 <= auto_tl_in_a_bits_data[23:16];
    end else if (_T_3769) begin
      if (dmiProgramBufferWrEnMaybe_6) begin
        programBufferMem_6 <= auto_dmi_in_a_bits_data[23:16];
      end
    end
    if (_T_13) begin
      programBufferMem_7 <= 8'h0;
    end else if (_T_24519) begin
      programBufferMem_7 <= auto_tl_in_a_bits_data[31:24];
    end else if (_T_3771) begin
      if (dmiProgramBufferWrEnMaybe_7) begin
        programBufferMem_7 <= auto_dmi_in_a_bits_data[31:24];
      end
    end
    if (_T_13) begin
      programBufferMem_8 <= 8'h0;
    end else if (_T_30272) begin
      programBufferMem_8 <= auto_tl_in_a_bits_data[7:0];
    end else if (_T_3773) begin
      if (dmiProgramBufferWrEnMaybe_8) begin
        programBufferMem_8 <= auto_dmi_in_a_bits_data[7:0];
      end
    end
    if (_T_13) begin
      programBufferMem_9 <= 8'h0;
    end else if (_T_30295) begin
      programBufferMem_9 <= auto_tl_in_a_bits_data[15:8];
    end else if (_T_3775) begin
      if (dmiProgramBufferWrEnMaybe_9) begin
        programBufferMem_9 <= auto_dmi_in_a_bits_data[15:8];
      end
    end
    if (_T_13) begin
      programBufferMem_10 <= 8'h0;
    end else if (_T_30320) begin
      programBufferMem_10 <= auto_tl_in_a_bits_data[23:16];
    end else if (_T_3777) begin
      if (dmiProgramBufferWrEnMaybe_10) begin
        programBufferMem_10 <= auto_dmi_in_a_bits_data[23:16];
      end
    end
    if (_T_13) begin
      programBufferMem_11 <= 8'h0;
    end else if (_T_30345) begin
      programBufferMem_11 <= auto_tl_in_a_bits_data[31:24];
    end else if (_T_3779) begin
      if (dmiProgramBufferWrEnMaybe_11) begin
        programBufferMem_11 <= auto_dmi_in_a_bits_data[31:24];
      end
    end
    if (_T_13) begin
      programBufferMem_12 <= 8'h0;
    end else if (_T_11219) begin
      programBufferMem_12 <= auto_tl_in_a_bits_data[7:0];
    end else if (_T_3781) begin
      if (dmiProgramBufferWrEnMaybe_12) begin
        programBufferMem_12 <= auto_dmi_in_a_bits_data[7:0];
      end
    end
    if (_T_13) begin
      programBufferMem_13 <= 8'h0;
    end else if (_T_11242) begin
      programBufferMem_13 <= auto_tl_in_a_bits_data[15:8];
    end else if (_T_3783) begin
      if (dmiProgramBufferWrEnMaybe_13) begin
        programBufferMem_13 <= auto_dmi_in_a_bits_data[15:8];
      end
    end
    if (_T_13) begin
      programBufferMem_14 <= 8'h0;
    end else if (_T_11267) begin
      programBufferMem_14 <= auto_tl_in_a_bits_data[23:16];
    end else if (_T_3785) begin
      if (dmiProgramBufferWrEnMaybe_14) begin
        programBufferMem_14 <= auto_dmi_in_a_bits_data[23:16];
      end
    end
    if (_T_13) begin
      programBufferMem_15 <= 8'h0;
    end else if (_T_11292) begin
      programBufferMem_15 <= auto_tl_in_a_bits_data[31:24];
    end else if (_T_3787) begin
      if (dmiProgramBufferWrEnMaybe_15) begin
        programBufferMem_15 <= auto_dmi_in_a_bits_data[31:24];
      end
    end
    if (_T_13) begin
      programBufferMem_16 <= 8'h0;
    end else if (_T_17254) begin
      programBufferMem_16 <= auto_tl_in_a_bits_data[7:0];
    end else if (_T_3789) begin
      if (dmiProgramBufferWrEnMaybe_16) begin
        programBufferMem_16 <= auto_dmi_in_a_bits_data[7:0];
      end
    end
    if (_T_13) begin
      programBufferMem_17 <= 8'h0;
    end else if (_T_17277) begin
      programBufferMem_17 <= auto_tl_in_a_bits_data[15:8];
    end else if (_T_3791) begin
      if (dmiProgramBufferWrEnMaybe_17) begin
        programBufferMem_17 <= auto_dmi_in_a_bits_data[15:8];
      end
    end
    if (_T_13) begin
      programBufferMem_18 <= 8'h0;
    end else if (_T_17302) begin
      programBufferMem_18 <= auto_tl_in_a_bits_data[23:16];
    end else if (_T_3793) begin
      if (dmiProgramBufferWrEnMaybe_18) begin
        programBufferMem_18 <= auto_dmi_in_a_bits_data[23:16];
      end
    end
    if (_T_13) begin
      programBufferMem_19 <= 8'h0;
    end else if (_T_17327) begin
      programBufferMem_19 <= auto_tl_in_a_bits_data[31:24];
    end else if (_T_3795) begin
      if (dmiProgramBufferWrEnMaybe_19) begin
        programBufferMem_19 <= auto_dmi_in_a_bits_data[31:24];
      end
    end
    if (_T_13) begin
      programBufferMem_20 <= 8'h0;
    end else if (_T_22429) begin
      programBufferMem_20 <= auto_tl_in_a_bits_data[7:0];
    end else if (_T_3797) begin
      if (dmiProgramBufferWrEnMaybe_20) begin
        programBufferMem_20 <= auto_dmi_in_a_bits_data[7:0];
      end
    end
    if (_T_13) begin
      programBufferMem_21 <= 8'h0;
    end else if (_T_22452) begin
      programBufferMem_21 <= auto_tl_in_a_bits_data[15:8];
    end else if (_T_3799) begin
      if (dmiProgramBufferWrEnMaybe_21) begin
        programBufferMem_21 <= auto_dmi_in_a_bits_data[15:8];
      end
    end
    if (_T_13) begin
      programBufferMem_22 <= 8'h0;
    end else if (_T_22477) begin
      programBufferMem_22 <= auto_tl_in_a_bits_data[23:16];
    end else if (_T_3801) begin
      if (dmiProgramBufferWrEnMaybe_22) begin
        programBufferMem_22 <= auto_dmi_in_a_bits_data[23:16];
      end
    end
    if (_T_13) begin
      programBufferMem_23 <= 8'h0;
    end else if (_T_22502) begin
      programBufferMem_23 <= auto_tl_in_a_bits_data[31:24];
    end else if (_T_3803) begin
      if (dmiProgramBufferWrEnMaybe_23) begin
        programBufferMem_23 <= auto_dmi_in_a_bits_data[31:24];
      end
    end
    if (_T_13) begin
      programBufferMem_24 <= 8'h0;
    end else if (_T_29094) begin
      programBufferMem_24 <= auto_tl_in_a_bits_data[7:0];
    end else if (_T_3805) begin
      if (dmiProgramBufferWrEnMaybe_24) begin
        programBufferMem_24 <= auto_dmi_in_a_bits_data[7:0];
      end
    end
    if (_T_13) begin
      programBufferMem_25 <= 8'h0;
    end else if (_T_29117) begin
      programBufferMem_25 <= auto_tl_in_a_bits_data[15:8];
    end else if (_T_3807) begin
      if (dmiProgramBufferWrEnMaybe_25) begin
        programBufferMem_25 <= auto_dmi_in_a_bits_data[15:8];
      end
    end
    if (_T_13) begin
      programBufferMem_26 <= 8'h0;
    end else if (_T_29142) begin
      programBufferMem_26 <= auto_tl_in_a_bits_data[23:16];
    end else if (_T_3809) begin
      if (dmiProgramBufferWrEnMaybe_26) begin
        programBufferMem_26 <= auto_dmi_in_a_bits_data[23:16];
      end
    end
    if (_T_13) begin
      programBufferMem_27 <= 8'h0;
    end else if (_T_29167) begin
      programBufferMem_27 <= auto_tl_in_a_bits_data[31:24];
    end else if (_T_3811) begin
      if (dmiProgramBufferWrEnMaybe_27) begin
        programBufferMem_27 <= auto_dmi_in_a_bits_data[31:24];
      end
    end
    if (_T_13) begin
      programBufferMem_28 <= 8'h0;
    end else if (_T_32890) begin
      programBufferMem_28 <= auto_tl_in_a_bits_data[7:0];
    end else if (_T_3813) begin
      if (dmiProgramBufferWrEnMaybe_28) begin
        programBufferMem_28 <= auto_dmi_in_a_bits_data[7:0];
      end
    end
    if (_T_13) begin
      programBufferMem_29 <= 8'h0;
    end else if (_T_32913) begin
      programBufferMem_29 <= auto_tl_in_a_bits_data[15:8];
    end else if (_T_3815) begin
      if (dmiProgramBufferWrEnMaybe_29) begin
        programBufferMem_29 <= auto_dmi_in_a_bits_data[15:8];
      end
    end
    if (_T_13) begin
      programBufferMem_30 <= 8'h0;
    end else if (_T_32938) begin
      programBufferMem_30 <= auto_tl_in_a_bits_data[23:16];
    end else if (_T_3817) begin
      if (dmiProgramBufferWrEnMaybe_30) begin
        programBufferMem_30 <= auto_dmi_in_a_bits_data[23:16];
      end
    end
    if (_T_13) begin
      programBufferMem_31 <= 8'h0;
    end else if (_T_32963) begin
      programBufferMem_31 <= auto_tl_in_a_bits_data[31:24];
    end else if (_T_3819) begin
      if (dmiProgramBufferWrEnMaybe_31) begin
        programBufferMem_31 <= auto_dmi_in_a_bits_data[31:24];
      end
    end
    if (_T_13) begin
      programBufferMem_32 <= 8'h0;
    end else if (_T_10671) begin
      programBufferMem_32 <= auto_tl_in_a_bits_data[7:0];
    end else if (_T_3821) begin
      if (dmiProgramBufferWrEnMaybe_32) begin
        programBufferMem_32 <= auto_dmi_in_a_bits_data[7:0];
      end
    end
    if (_T_13) begin
      programBufferMem_33 <= 8'h0;
    end else if (_T_10694) begin
      programBufferMem_33 <= auto_tl_in_a_bits_data[15:8];
    end else if (_T_3823) begin
      if (dmiProgramBufferWrEnMaybe_33) begin
        programBufferMem_33 <= auto_dmi_in_a_bits_data[15:8];
      end
    end
    if (_T_13) begin
      programBufferMem_34 <= 8'h0;
    end else if (_T_10719) begin
      programBufferMem_34 <= auto_tl_in_a_bits_data[23:16];
    end else if (_T_3825) begin
      if (dmiProgramBufferWrEnMaybe_34) begin
        programBufferMem_34 <= auto_dmi_in_a_bits_data[23:16];
      end
    end
    if (_T_13) begin
      programBufferMem_35 <= 8'h0;
    end else if (_T_10744) begin
      programBufferMem_35 <= auto_tl_in_a_bits_data[31:24];
    end else if (_T_3827) begin
      if (dmiProgramBufferWrEnMaybe_35) begin
        programBufferMem_35 <= auto_dmi_in_a_bits_data[31:24];
      end
    end
    if (_T_13) begin
      programBufferMem_36 <= 8'h0;
    end else if (_T_7603) begin
      programBufferMem_36 <= auto_tl_in_a_bits_data[7:0];
    end else if (_T_3829) begin
      if (dmiProgramBufferWrEnMaybe_36) begin
        programBufferMem_36 <= auto_dmi_in_a_bits_data[7:0];
      end
    end
    if (_T_13) begin
      programBufferMem_37 <= 8'h0;
    end else if (_T_7626) begin
      programBufferMem_37 <= auto_tl_in_a_bits_data[15:8];
    end else if (_T_3831) begin
      if (dmiProgramBufferWrEnMaybe_37) begin
        programBufferMem_37 <= auto_dmi_in_a_bits_data[15:8];
      end
    end
    if (_T_13) begin
      programBufferMem_38 <= 8'h0;
    end else if (_T_7651) begin
      programBufferMem_38 <= auto_tl_in_a_bits_data[23:16];
    end else if (_T_3833) begin
      if (dmiProgramBufferWrEnMaybe_38) begin
        programBufferMem_38 <= auto_dmi_in_a_bits_data[23:16];
      end
    end
    if (_T_13) begin
      programBufferMem_39 <= 8'h0;
    end else if (_T_7676) begin
      programBufferMem_39 <= auto_tl_in_a_bits_data[31:24];
    end else if (_T_3835) begin
      if (dmiProgramBufferWrEnMaybe_39) begin
        programBufferMem_39 <= auto_dmi_in_a_bits_data[31:24];
      end
    end
    if (_T_13) begin
      programBufferMem_40 <= 8'h0;
    end else if (_T_27445) begin
      programBufferMem_40 <= auto_tl_in_a_bits_data[7:0];
    end else if (_T_3837) begin
      if (dmiProgramBufferWrEnMaybe_40) begin
        programBufferMem_40 <= auto_dmi_in_a_bits_data[7:0];
      end
    end
    if (_T_13) begin
      programBufferMem_41 <= 8'h0;
    end else if (_T_27468) begin
      programBufferMem_41 <= auto_tl_in_a_bits_data[15:8];
    end else if (_T_3839) begin
      if (dmiProgramBufferWrEnMaybe_41) begin
        programBufferMem_41 <= auto_dmi_in_a_bits_data[15:8];
      end
    end
    if (_T_13) begin
      programBufferMem_42 <= 8'h0;
    end else if (_T_27493) begin
      programBufferMem_42 <= auto_tl_in_a_bits_data[23:16];
    end else if (_T_3841) begin
      if (dmiProgramBufferWrEnMaybe_42) begin
        programBufferMem_42 <= auto_dmi_in_a_bits_data[23:16];
      end
    end
    if (_T_13) begin
      programBufferMem_43 <= 8'h0;
    end else if (_T_27518) begin
      programBufferMem_43 <= auto_tl_in_a_bits_data[31:24];
    end else if (_T_3843) begin
      if (dmiProgramBufferWrEnMaybe_43) begin
        programBufferMem_43 <= auto_dmi_in_a_bits_data[31:24];
      end
    end
    if (_T_13) begin
      programBufferMem_44 <= 8'h0;
    end else if (_T_20793) begin
      programBufferMem_44 <= auto_tl_in_a_bits_data[7:0];
    end else if (_T_3845) begin
      if (dmiProgramBufferWrEnMaybe_44) begin
        programBufferMem_44 <= auto_dmi_in_a_bits_data[7:0];
      end
    end
    if (_T_13) begin
      programBufferMem_45 <= 8'h0;
    end else if (_T_20816) begin
      programBufferMem_45 <= auto_tl_in_a_bits_data[15:8];
    end else if (_T_3847) begin
      if (dmiProgramBufferWrEnMaybe_45) begin
        programBufferMem_45 <= auto_dmi_in_a_bits_data[15:8];
      end
    end
    if (_T_13) begin
      programBufferMem_46 <= 8'h0;
    end else if (_T_20841) begin
      programBufferMem_46 <= auto_tl_in_a_bits_data[23:16];
    end else if (_T_3849) begin
      if (dmiProgramBufferWrEnMaybe_46) begin
        programBufferMem_46 <= auto_dmi_in_a_bits_data[23:16];
      end
    end
    if (_T_13) begin
      programBufferMem_47 <= 8'h0;
    end else if (_T_20866) begin
      programBufferMem_47 <= auto_tl_in_a_bits_data[31:24];
    end else if (_T_3851) begin
      if (dmiProgramBufferWrEnMaybe_47) begin
        programBufferMem_47 <= auto_dmi_in_a_bits_data[31:24];
      end
    end
    if (_T_13) begin
      programBufferMem_48 <= 8'h0;
    end else if (_T_13686) begin
      programBufferMem_48 <= auto_tl_in_a_bits_data[7:0];
    end else if (_T_3853) begin
      if (dmiProgramBufferWrEnMaybe_48) begin
        programBufferMem_48 <= auto_dmi_in_a_bits_data[7:0];
      end
    end
    if (_T_13) begin
      programBufferMem_49 <= 8'h0;
    end else if (_T_13709) begin
      programBufferMem_49 <= auto_tl_in_a_bits_data[15:8];
    end else if (_T_3855) begin
      if (dmiProgramBufferWrEnMaybe_49) begin
        programBufferMem_49 <= auto_dmi_in_a_bits_data[15:8];
      end
    end
    if (_T_13) begin
      programBufferMem_50 <= 8'h0;
    end else if (_T_13734) begin
      programBufferMem_50 <= auto_tl_in_a_bits_data[23:16];
    end else if (_T_3857) begin
      if (dmiProgramBufferWrEnMaybe_50) begin
        programBufferMem_50 <= auto_dmi_in_a_bits_data[23:16];
      end
    end
    if (_T_13) begin
      programBufferMem_51 <= 8'h0;
    end else if (_T_13759) begin
      programBufferMem_51 <= auto_tl_in_a_bits_data[31:24];
    end else if (_T_3859) begin
      if (dmiProgramBufferWrEnMaybe_51) begin
        programBufferMem_51 <= auto_dmi_in_a_bits_data[31:24];
      end
    end
    if (_T_13) begin
      programBufferMem_52 <= 8'h0;
    end else if (_T_11947) begin
      programBufferMem_52 <= auto_tl_in_a_bits_data[7:0];
    end else if (_T_3861) begin
      if (dmiProgramBufferWrEnMaybe_52) begin
        programBufferMem_52 <= auto_dmi_in_a_bits_data[7:0];
      end
    end
    if (_T_13) begin
      programBufferMem_53 <= 8'h0;
    end else if (_T_11970) begin
      programBufferMem_53 <= auto_tl_in_a_bits_data[15:8];
    end else if (_T_3863) begin
      if (dmiProgramBufferWrEnMaybe_53) begin
        programBufferMem_53 <= auto_dmi_in_a_bits_data[15:8];
      end
    end
    if (_T_13) begin
      programBufferMem_54 <= 8'h0;
    end else if (_T_11995) begin
      programBufferMem_54 <= auto_tl_in_a_bits_data[23:16];
    end else if (_T_3865) begin
      if (dmiProgramBufferWrEnMaybe_54) begin
        programBufferMem_54 <= auto_dmi_in_a_bits_data[23:16];
      end
    end
    if (_T_13) begin
      programBufferMem_55 <= 8'h0;
    end else if (_T_12020) begin
      programBufferMem_55 <= auto_tl_in_a_bits_data[31:24];
    end else if (_T_3867) begin
      if (dmiProgramBufferWrEnMaybe_55) begin
        programBufferMem_55 <= auto_dmi_in_a_bits_data[31:24];
      end
    end
    if (_T_13) begin
      programBufferMem_56 <= 8'h0;
    end else if (_T_33078) begin
      programBufferMem_56 <= auto_tl_in_a_bits_data[7:0];
    end else if (_T_3869) begin
      if (dmiProgramBufferWrEnMaybe_56) begin
        programBufferMem_56 <= auto_dmi_in_a_bits_data[7:0];
      end
    end
    if (_T_13) begin
      programBufferMem_57 <= 8'h0;
    end else if (_T_33101) begin
      programBufferMem_57 <= auto_tl_in_a_bits_data[15:8];
    end else if (_T_3871) begin
      if (dmiProgramBufferWrEnMaybe_57) begin
        programBufferMem_57 <= auto_dmi_in_a_bits_data[15:8];
      end
    end
    if (_T_13) begin
      programBufferMem_58 <= 8'h0;
    end else if (_T_33126) begin
      programBufferMem_58 <= auto_tl_in_a_bits_data[23:16];
    end else if (_T_3873) begin
      if (dmiProgramBufferWrEnMaybe_58) begin
        programBufferMem_58 <= auto_dmi_in_a_bits_data[23:16];
      end
    end
    if (_T_13) begin
      programBufferMem_59 <= 8'h0;
    end else if (_T_33151) begin
      programBufferMem_59 <= auto_tl_in_a_bits_data[31:24];
    end else if (_T_3875) begin
      if (dmiProgramBufferWrEnMaybe_59) begin
        programBufferMem_59 <= auto_dmi_in_a_bits_data[31:24];
      end
    end
    if (_T_13) begin
      programBufferMem_60 <= 8'h0;
    end else if (_T_23268) begin
      programBufferMem_60 <= auto_tl_in_a_bits_data[7:0];
    end else if (_T_3877) begin
      if (dmiProgramBufferWrEnMaybe_60) begin
        programBufferMem_60 <= auto_dmi_in_a_bits_data[7:0];
      end
    end
    if (_T_13) begin
      programBufferMem_61 <= 8'h0;
    end else if (_T_23291) begin
      programBufferMem_61 <= auto_tl_in_a_bits_data[15:8];
    end else if (_T_3879) begin
      if (dmiProgramBufferWrEnMaybe_61) begin
        programBufferMem_61 <= auto_dmi_in_a_bits_data[15:8];
      end
    end
    if (_T_13) begin
      programBufferMem_62 <= 8'h0;
    end else if (_T_23316) begin
      programBufferMem_62 <= auto_tl_in_a_bits_data[23:16];
    end else if (_T_3881) begin
      if (dmiProgramBufferWrEnMaybe_62) begin
        programBufferMem_62 <= auto_dmi_in_a_bits_data[23:16];
      end
    end
    if (_T_13) begin
      programBufferMem_63 <= 8'h0;
    end else if (_T_23341) begin
      programBufferMem_63 <= auto_tl_in_a_bits_data[31:24];
    end else if (_T_3883) begin
      if (dmiProgramBufferWrEnMaybe_63) begin
        programBufferMem_63 <= auto_dmi_in_a_bits_data[31:24];
      end
    end
    if (_T_13) begin
      goReg <= 1'h0;
    end else begin
      goReg <= _GEN_407;
    end
    if (goAbstract) begin
      if (accessRegisterCommandReg_transfer) begin
        if (accessRegisterCommandReg_write) begin
          abstractGeneratedMem_0 <= _T_3979;
        end else begin
          abstractGeneratedMem_0 <= _T_3984;
        end
      end else begin
        abstractGeneratedMem_0 <= 32'h13;
      end
    end
    if (goAbstract) begin
      if (accessRegisterCommandReg_postexec) begin
        abstractGeneratedMem_1 <= 32'h13;
      end else begin
        abstractGeneratedMem_1 <= 32'h100073;
      end
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_3886 & _T_3938) begin
          $fwrite(32'h80000002,"Assertion failed: Unexpected 'GOING' hart.\n    at Debug.scala:1389 assert(hartGoingId === 0.U, \"Unexpected 'GOING' hart.\")//Chisel3 #540 %%x, expected %%x\", hartGoingId, 0.U)\n"); // @[Debug.scala 1389:15:freechips.rocketchip.system.DefaultRV32Config.fir@115473.12]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_3886 & _T_3938) begin
          $fatal; // @[Debug.scala 1389:15:freechips.rocketchip.system.DefaultRV32Config.fir@115474.12]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_3895 & _T_3938) begin
          $fwrite(32'h80000002,"Assertion failed: Unexpected 'EXCEPTION' hart\n    at Debug.scala:1653 assert(hartExceptionId === 0.U, \"Unexpected 'EXCEPTION' hart\")//Chisel3 #540, %%x, expected %%x\", hartExceptionId, 0.U)\n"); // @[Debug.scala 1653:15:freechips.rocketchip.system.DefaultRV32Config.fir@168777.14]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_3895 & _T_3938) begin
          $fatal; // @[Debug.scala 1653:15:freechips.rocketchip.system.DefaultRV32Config.fir@168778.14]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_3906 & _T_44831) begin
          $fwrite(32'h80000002,"Assertion failed: Should not be in custom state unless we need it.\n    at Debug.scala:1658 assert(needCustom.B, \"Should not be in custom state unless we need it.\")\n"); // @[Debug.scala 1658:13:freechips.rocketchip.system.DefaultRV32Config.fir@168791.14]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_3906 & _T_44831) begin
          $fatal; // @[Debug.scala 1658:13:freechips.rocketchip.system.DefaultRV32Config.fir@168792.14]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_44843) begin
          $fwrite(32'h80000002,"Assertion failed: Unexpected EXCEPTION write: should only get it in Debug Module EXEC state\n    at Debug.scala:1671 assert ((!io.dmactive || !hartExceptionWrEn || ctrlStateReg === CtrlState(Exec)),\n"); // @[Debug.scala 1671:12:freechips.rocketchip.system.DefaultRV32Config.fir@168818.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_44843) begin
          $fatal; // @[Debug.scala 1671:12:freechips.rocketchip.system.DefaultRV32Config.fir@168819.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      hrDebugInt_0 <= 1'h0;
    end else if (_T_13) begin
      hrDebugInt_0 <= 1'h0;
    end else begin
      hrDebugInt_0 <= _T_26;
    end
  end
endmodule
