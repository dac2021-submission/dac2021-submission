module AXI4ToTL( // @[:freechips.rocketchip.system.DefaultRV32Config.fir@39531.2]
  input         clock, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@39532.4]
  input         reset, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@39533.4]
  output        auto_in_aw_ready, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@39534.4]
  input         auto_in_aw_valid, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@39534.4]
  input         auto_in_aw_bits_id, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@39534.4]
  input  [31:0] auto_in_aw_bits_addr, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@39534.4]
  input  [7:0]  auto_in_aw_bits_len, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@39534.4]
  input  [2:0]  auto_in_aw_bits_size, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@39534.4]
  input  [3:0]  auto_in_aw_bits_cache, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@39534.4]
  input  [2:0]  auto_in_aw_bits_prot, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@39534.4]
  output        auto_in_w_ready, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@39534.4]
  input         auto_in_w_valid, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@39534.4]
  input  [63:0] auto_in_w_bits_data, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@39534.4]
  input  [7:0]  auto_in_w_bits_strb, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@39534.4]
  input         auto_in_w_bits_last, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@39534.4]
  input         auto_in_b_ready, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@39534.4]
  output        auto_in_b_valid, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@39534.4]
  output        auto_in_b_bits_id, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@39534.4]
  output [1:0]  auto_in_b_bits_resp, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@39534.4]
  output        auto_in_ar_ready, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@39534.4]
  input         auto_in_ar_valid, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@39534.4]
  input         auto_in_ar_bits_id, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@39534.4]
  input  [31:0] auto_in_ar_bits_addr, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@39534.4]
  input  [7:0]  auto_in_ar_bits_len, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@39534.4]
  input  [2:0]  auto_in_ar_bits_size, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@39534.4]
  input  [3:0]  auto_in_ar_bits_cache, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@39534.4]
  input  [2:0]  auto_in_ar_bits_prot, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@39534.4]
  input         auto_in_r_ready, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@39534.4]
  output        auto_in_r_valid, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@39534.4]
  output        auto_in_r_bits_id, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@39534.4]
  output [63:0] auto_in_r_bits_data, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@39534.4]
  output [1:0]  auto_in_r_bits_resp, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@39534.4]
  output        auto_in_r_bits_last, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@39534.4]
  input         auto_out_a_ready, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@39534.4]
  output        auto_out_a_valid, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@39534.4]
  output [2:0]  auto_out_a_bits_opcode, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@39534.4]
  output [2:0]  auto_out_a_bits_param, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@39534.4]
  output [3:0]  auto_out_a_bits_size, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@39534.4]
  output [3:0]  auto_out_a_bits_source, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@39534.4]
  output [31:0] auto_out_a_bits_address, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@39534.4]
  output        auto_out_a_bits_user_amba_prot_bufferable, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@39534.4]
  output        auto_out_a_bits_user_amba_prot_modifiable, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@39534.4]
  output        auto_out_a_bits_user_amba_prot_readalloc, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@39534.4]
  output        auto_out_a_bits_user_amba_prot_writealloc, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@39534.4]
  output        auto_out_a_bits_user_amba_prot_privileged, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@39534.4]
  output        auto_out_a_bits_user_amba_prot_secure, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@39534.4]
  output        auto_out_a_bits_user_amba_prot_fetch, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@39534.4]
  output [7:0]  auto_out_a_bits_mask, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@39534.4]
  output [63:0] auto_out_a_bits_data, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@39534.4]
  output        auto_out_a_bits_corrupt, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@39534.4]
  output        auto_out_d_ready, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@39534.4]
  input         auto_out_d_valid, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@39534.4]
  input  [2:0]  auto_out_d_bits_opcode, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@39534.4]
  input  [3:0]  auto_out_d_bits_size, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@39534.4]
  input  [3:0]  auto_out_d_bits_source, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@39534.4]
  input         auto_out_d_bits_denied, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@39534.4]
  input  [63:0] auto_out_d_bits_data, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@39534.4]
  input         auto_out_d_bits_corrupt // @[:freechips.rocketchip.system.DefaultRV32Config.fir@39534.4]
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
`endif // RANDOMIZE_REG_INIT
  wire  Queue_clock; // @[Decoupled.scala 287:21:freechips.rocketchip.system.DefaultRV32Config.fir@40414.4]
  wire  Queue_reset; // @[Decoupled.scala 287:21:freechips.rocketchip.system.DefaultRV32Config.fir@40414.4]
  wire  Queue_io_enq_ready; // @[Decoupled.scala 287:21:freechips.rocketchip.system.DefaultRV32Config.fir@40414.4]
  wire  Queue_io_enq_valid; // @[Decoupled.scala 287:21:freechips.rocketchip.system.DefaultRV32Config.fir@40414.4]
  wire  Queue_io_enq_bits_id; // @[Decoupled.scala 287:21:freechips.rocketchip.system.DefaultRV32Config.fir@40414.4]
  wire [63:0] Queue_io_enq_bits_data; // @[Decoupled.scala 287:21:freechips.rocketchip.system.DefaultRV32Config.fir@40414.4]
  wire [1:0] Queue_io_enq_bits_resp; // @[Decoupled.scala 287:21:freechips.rocketchip.system.DefaultRV32Config.fir@40414.4]
  wire  Queue_io_enq_bits_last; // @[Decoupled.scala 287:21:freechips.rocketchip.system.DefaultRV32Config.fir@40414.4]
  wire  Queue_io_deq_ready; // @[Decoupled.scala 287:21:freechips.rocketchip.system.DefaultRV32Config.fir@40414.4]
  wire  Queue_io_deq_valid; // @[Decoupled.scala 287:21:freechips.rocketchip.system.DefaultRV32Config.fir@40414.4]
  wire  Queue_io_deq_bits_id; // @[Decoupled.scala 287:21:freechips.rocketchip.system.DefaultRV32Config.fir@40414.4]
  wire [63:0] Queue_io_deq_bits_data; // @[Decoupled.scala 287:21:freechips.rocketchip.system.DefaultRV32Config.fir@40414.4]
  wire [1:0] Queue_io_deq_bits_resp; // @[Decoupled.scala 287:21:freechips.rocketchip.system.DefaultRV32Config.fir@40414.4]
  wire  Queue_io_deq_bits_last; // @[Decoupled.scala 287:21:freechips.rocketchip.system.DefaultRV32Config.fir@40414.4]
  wire  Queue_1_clock; // @[Decoupled.scala 287:21:freechips.rocketchip.system.DefaultRV32Config.fir@40439.4]
  wire  Queue_1_reset; // @[Decoupled.scala 287:21:freechips.rocketchip.system.DefaultRV32Config.fir@40439.4]
  wire  Queue_1_io_enq_ready; // @[Decoupled.scala 287:21:freechips.rocketchip.system.DefaultRV32Config.fir@40439.4]
  wire  Queue_1_io_enq_valid; // @[Decoupled.scala 287:21:freechips.rocketchip.system.DefaultRV32Config.fir@40439.4]
  wire  Queue_1_io_enq_bits_id; // @[Decoupled.scala 287:21:freechips.rocketchip.system.DefaultRV32Config.fir@40439.4]
  wire [1:0] Queue_1_io_enq_bits_resp; // @[Decoupled.scala 287:21:freechips.rocketchip.system.DefaultRV32Config.fir@40439.4]
  wire  Queue_1_io_deq_ready; // @[Decoupled.scala 287:21:freechips.rocketchip.system.DefaultRV32Config.fir@40439.4]
  wire  Queue_1_io_deq_valid; // @[Decoupled.scala 287:21:freechips.rocketchip.system.DefaultRV32Config.fir@40439.4]
  wire  Queue_1_io_deq_bits_id; // @[Decoupled.scala 287:21:freechips.rocketchip.system.DefaultRV32Config.fir@40439.4]
  wire [1:0] Queue_1_io_deq_bits_resp; // @[Decoupled.scala 287:21:freechips.rocketchip.system.DefaultRV32Config.fir@40439.4]
  wire [15:0] _T_3; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@39547.4]
  wire [22:0] _GEN_16; // @[Bundles.scala 30:21:freechips.rocketchip.system.DefaultRV32Config.fir@39548.4]
  wire [22:0] _T_4; // @[Bundles.scala 30:21:freechips.rocketchip.system.DefaultRV32Config.fir@39548.4]
  wire [15:0] _T_6; // @[package.scala 205:35:freechips.rocketchip.system.DefaultRV32Config.fir@39550.4]
  wire [15:0] _T_7; // @[package.scala 205:40:freechips.rocketchip.system.DefaultRV32Config.fir@39551.4]
  wire [15:0] _T_8; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@39552.4]
  wire [15:0] _T_9; // @[package.scala 205:53:freechips.rocketchip.system.DefaultRV32Config.fir@39553.4]
  wire [15:0] _T_10; // @[package.scala 205:51:freechips.rocketchip.system.DefaultRV32Config.fir@39554.4]
  wire  _T_13; // @[OneHot.scala 32:14:freechips.rocketchip.system.DefaultRV32Config.fir@39557.4]
  wire [7:0] _T_14; // @[OneHot.scala 32:28:freechips.rocketchip.system.DefaultRV32Config.fir@39558.4]
  wire  _T_17; // @[OneHot.scala 32:14:freechips.rocketchip.system.DefaultRV32Config.fir@39561.4]
  wire [3:0] _T_18; // @[OneHot.scala 32:28:freechips.rocketchip.system.DefaultRV32Config.fir@39562.4]
  wire  _T_21; // @[OneHot.scala 32:14:freechips.rocketchip.system.DefaultRV32Config.fir@39565.4]
  wire [1:0] _T_22; // @[OneHot.scala 32:28:freechips.rocketchip.system.DefaultRV32Config.fir@39566.4]
  wire [3:0] _T_26; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@39570.4]
  wire  _T_28; // @[Parameters.scala 93:42:freechips.rocketchip.system.DefaultRV32Config.fir@39572.4]
  wire [31:0] _T_31; // @[Parameters.scala 137:31:freechips.rocketchip.system.DefaultRV32Config.fir@39575.4]
  wire [32:0] _T_32; // @[Parameters.scala 137:49:freechips.rocketchip.system.DefaultRV32Config.fir@39576.4]
  wire [32:0] _T_34; // @[Parameters.scala 137:52:freechips.rocketchip.system.DefaultRV32Config.fir@39578.4]
  wire  _T_35; // @[Parameters.scala 137:67:freechips.rocketchip.system.DefaultRV32Config.fir@39579.4]
  wire  _T_36; // @[Parameters.scala 551:56:freechips.rocketchip.system.DefaultRV32Config.fir@39580.4]
  wire  _T_38; // @[Parameters.scala 93:42:freechips.rocketchip.system.DefaultRV32Config.fir@39582.4]
  wire [32:0] _T_42; // @[Parameters.scala 137:49:freechips.rocketchip.system.DefaultRV32Config.fir@39586.4]
  wire [32:0] _T_44; // @[Parameters.scala 137:52:freechips.rocketchip.system.DefaultRV32Config.fir@39588.4]
  wire  _T_45; // @[Parameters.scala 137:67:freechips.rocketchip.system.DefaultRV32Config.fir@39589.4]
  wire [31:0] _T_46; // @[Parameters.scala 137:31:freechips.rocketchip.system.DefaultRV32Config.fir@39590.4]
  wire [32:0] _T_47; // @[Parameters.scala 137:49:freechips.rocketchip.system.DefaultRV32Config.fir@39591.4]
  wire [32:0] _T_49; // @[Parameters.scala 137:52:freechips.rocketchip.system.DefaultRV32Config.fir@39593.4]
  wire  _T_50; // @[Parameters.scala 137:67:freechips.rocketchip.system.DefaultRV32Config.fir@39594.4]
  wire [31:0] _T_51; // @[Parameters.scala 137:31:freechips.rocketchip.system.DefaultRV32Config.fir@39595.4]
  wire [32:0] _T_52; // @[Parameters.scala 137:49:freechips.rocketchip.system.DefaultRV32Config.fir@39596.4]
  wire [32:0] _T_54; // @[Parameters.scala 137:52:freechips.rocketchip.system.DefaultRV32Config.fir@39598.4]
  wire  _T_55; // @[Parameters.scala 137:67:freechips.rocketchip.system.DefaultRV32Config.fir@39599.4]
  wire [31:0] _T_56; // @[Parameters.scala 137:31:freechips.rocketchip.system.DefaultRV32Config.fir@39600.4]
  wire [32:0] _T_57; // @[Parameters.scala 137:49:freechips.rocketchip.system.DefaultRV32Config.fir@39601.4]
  wire [32:0] _T_59; // @[Parameters.scala 137:52:freechips.rocketchip.system.DefaultRV32Config.fir@39603.4]
  wire  _T_60; // @[Parameters.scala 137:67:freechips.rocketchip.system.DefaultRV32Config.fir@39604.4]
  wire [31:0] _T_61; // @[Parameters.scala 137:31:freechips.rocketchip.system.DefaultRV32Config.fir@39605.4]
  wire [32:0] _T_62; // @[Parameters.scala 137:49:freechips.rocketchip.system.DefaultRV32Config.fir@39606.4]
  wire [32:0] _T_64; // @[Parameters.scala 137:52:freechips.rocketchip.system.DefaultRV32Config.fir@39608.4]
  wire  _T_65; // @[Parameters.scala 137:67:freechips.rocketchip.system.DefaultRV32Config.fir@39609.4]
  wire [31:0] _T_66; // @[Parameters.scala 137:31:freechips.rocketchip.system.DefaultRV32Config.fir@39610.4]
  wire [32:0] _T_67; // @[Parameters.scala 137:49:freechips.rocketchip.system.DefaultRV32Config.fir@39611.4]
  wire [32:0] _T_69; // @[Parameters.scala 137:52:freechips.rocketchip.system.DefaultRV32Config.fir@39613.4]
  wire  _T_70; // @[Parameters.scala 137:67:freechips.rocketchip.system.DefaultRV32Config.fir@39614.4]
  wire  _T_71; // @[Parameters.scala 552:42:freechips.rocketchip.system.DefaultRV32Config.fir@39615.4]
  wire  _T_72; // @[Parameters.scala 552:42:freechips.rocketchip.system.DefaultRV32Config.fir@39616.4]
  wire  _T_73; // @[Parameters.scala 552:42:freechips.rocketchip.system.DefaultRV32Config.fir@39617.4]
  wire  _T_74; // @[Parameters.scala 552:42:freechips.rocketchip.system.DefaultRV32Config.fir@39618.4]
  wire  _T_75; // @[Parameters.scala 552:42:freechips.rocketchip.system.DefaultRV32Config.fir@39619.4]
  wire  _T_76; // @[Parameters.scala 551:56:freechips.rocketchip.system.DefaultRV32Config.fir@39620.4]
  wire  _T_78; // @[Parameters.scala 553:30:freechips.rocketchip.system.DefaultRV32Config.fir@39622.4]
  wire [13:0] _GEN_17; // @[ToTL.scala 89:59:freechips.rocketchip.system.DefaultRV32Config.fir@39624.4]
  wire [13:0] _T_80; // @[ToTL.scala 89:59:freechips.rocketchip.system.DefaultRV32Config.fir@39624.4]
  wire [31:0] _T_81; // @[ToTL.scala 89:23:freechips.rocketchip.system.DefaultRV32Config.fir@39625.4]
  reg [2:0] _T_83_0; // @[ToTL.scala 90:28:freechips.rocketchip.system.DefaultRV32Config.fir@39630.4]
  reg [2:0] _T_83_1; // @[ToTL.scala 90:28:freechips.rocketchip.system.DefaultRV32Config.fir@39630.4]
  wire [2:0] _GEN_1; // @[ToTL.scala 94:50:freechips.rocketchip.system.DefaultRV32Config.fir@39631.4]
  wire  _T_87; // @[ToTL.scala 97:15:freechips.rocketchip.system.DefaultRV32Config.fir@39634.4]
  wire [29:0] _T_89; // @[package.scala 207:77:freechips.rocketchip.system.DefaultRV32Config.fir@39636.4]
  wire [14:0] _T_91; // @[package.scala 207:46:freechips.rocketchip.system.DefaultRV32Config.fir@39638.4]
  wire  _T_92; // @[ToTL.scala 97:39:freechips.rocketchip.system.DefaultRV32Config.fir@39639.4]
  wire  _T_93; // @[ToTL.scala 97:28:freechips.rocketchip.system.DefaultRV32Config.fir@39640.4]
  wire  _T_95; // @[ToTL.scala 97:14:freechips.rocketchip.system.DefaultRV32Config.fir@39642.4]
  wire  _T_96; // @[ToTL.scala 97:14:freechips.rocketchip.system.DefaultRV32Config.fir@39643.4]
  wire [3:0] _T_152; // @[OneHot.scala 65:12:freechips.rocketchip.system.DefaultRV32Config.fir@39711.4]
  wire [2:0] _T_154; // @[Misc.scala 201:81:freechips.rocketchip.system.DefaultRV32Config.fir@39713.4]
  wire  _T_155; // @[Misc.scala 205:21:freechips.rocketchip.system.DefaultRV32Config.fir@39714.4]
  wire  _T_158; // @[Misc.scala 210:20:freechips.rocketchip.system.DefaultRV32Config.fir@39717.4]
  wire  _T_160; // @[Misc.scala 214:38:freechips.rocketchip.system.DefaultRV32Config.fir@39719.4]
  wire  _T_161; // @[Misc.scala 214:29:freechips.rocketchip.system.DefaultRV32Config.fir@39720.4]
  wire  _T_163; // @[Misc.scala 214:38:freechips.rocketchip.system.DefaultRV32Config.fir@39722.4]
  wire  _T_164; // @[Misc.scala 214:29:freechips.rocketchip.system.DefaultRV32Config.fir@39723.4]
  wire  _T_167; // @[Misc.scala 210:20:freechips.rocketchip.system.DefaultRV32Config.fir@39726.4]
  wire  _T_168; // @[Misc.scala 213:27:freechips.rocketchip.system.DefaultRV32Config.fir@39727.4]
  wire  _T_169; // @[Misc.scala 214:38:freechips.rocketchip.system.DefaultRV32Config.fir@39728.4]
  wire  _T_170; // @[Misc.scala 214:29:freechips.rocketchip.system.DefaultRV32Config.fir@39729.4]
  wire  _T_171; // @[Misc.scala 213:27:freechips.rocketchip.system.DefaultRV32Config.fir@39730.4]
  wire  _T_172; // @[Misc.scala 214:38:freechips.rocketchip.system.DefaultRV32Config.fir@39731.4]
  wire  _T_173; // @[Misc.scala 214:29:freechips.rocketchip.system.DefaultRV32Config.fir@39732.4]
  wire  _T_174; // @[Misc.scala 213:27:freechips.rocketchip.system.DefaultRV32Config.fir@39733.4]
  wire  _T_175; // @[Misc.scala 214:38:freechips.rocketchip.system.DefaultRV32Config.fir@39734.4]
  wire  _T_176; // @[Misc.scala 214:29:freechips.rocketchip.system.DefaultRV32Config.fir@39735.4]
  wire  _T_177; // @[Misc.scala 213:27:freechips.rocketchip.system.DefaultRV32Config.fir@39736.4]
  wire  _T_178; // @[Misc.scala 214:38:freechips.rocketchip.system.DefaultRV32Config.fir@39737.4]
  wire  _T_179; // @[Misc.scala 214:29:freechips.rocketchip.system.DefaultRV32Config.fir@39738.4]
  wire  _T_182; // @[Misc.scala 210:20:freechips.rocketchip.system.DefaultRV32Config.fir@39741.4]
  wire  _T_183; // @[Misc.scala 213:27:freechips.rocketchip.system.DefaultRV32Config.fir@39742.4]
  wire  _T_184; // @[Misc.scala 214:38:freechips.rocketchip.system.DefaultRV32Config.fir@39743.4]
  wire  _T_185; // @[Misc.scala 214:29:freechips.rocketchip.system.DefaultRV32Config.fir@39744.4]
  wire  _T_186; // @[Misc.scala 213:27:freechips.rocketchip.system.DefaultRV32Config.fir@39745.4]
  wire  _T_187; // @[Misc.scala 214:38:freechips.rocketchip.system.DefaultRV32Config.fir@39746.4]
  wire  _T_188; // @[Misc.scala 214:29:freechips.rocketchip.system.DefaultRV32Config.fir@39747.4]
  wire  _T_189; // @[Misc.scala 213:27:freechips.rocketchip.system.DefaultRV32Config.fir@39748.4]
  wire  _T_190; // @[Misc.scala 214:38:freechips.rocketchip.system.DefaultRV32Config.fir@39749.4]
  wire  _T_191; // @[Misc.scala 214:29:freechips.rocketchip.system.DefaultRV32Config.fir@39750.4]
  wire  _T_192; // @[Misc.scala 213:27:freechips.rocketchip.system.DefaultRV32Config.fir@39751.4]
  wire  _T_193; // @[Misc.scala 214:38:freechips.rocketchip.system.DefaultRV32Config.fir@39752.4]
  wire  _T_194; // @[Misc.scala 214:29:freechips.rocketchip.system.DefaultRV32Config.fir@39753.4]
  wire  _T_195; // @[Misc.scala 213:27:freechips.rocketchip.system.DefaultRV32Config.fir@39754.4]
  wire  _T_196; // @[Misc.scala 214:38:freechips.rocketchip.system.DefaultRV32Config.fir@39755.4]
  wire  _T_197; // @[Misc.scala 214:29:freechips.rocketchip.system.DefaultRV32Config.fir@39756.4]
  wire  _T_198; // @[Misc.scala 213:27:freechips.rocketchip.system.DefaultRV32Config.fir@39757.4]
  wire  _T_199; // @[Misc.scala 214:38:freechips.rocketchip.system.DefaultRV32Config.fir@39758.4]
  wire  _T_200; // @[Misc.scala 214:29:freechips.rocketchip.system.DefaultRV32Config.fir@39759.4]
  wire  _T_201; // @[Misc.scala 213:27:freechips.rocketchip.system.DefaultRV32Config.fir@39760.4]
  wire  _T_202; // @[Misc.scala 214:38:freechips.rocketchip.system.DefaultRV32Config.fir@39761.4]
  wire  _T_203; // @[Misc.scala 214:29:freechips.rocketchip.system.DefaultRV32Config.fir@39762.4]
  wire  _T_204; // @[Misc.scala 213:27:freechips.rocketchip.system.DefaultRV32Config.fir@39763.4]
  wire  _T_205; // @[Misc.scala 214:38:freechips.rocketchip.system.DefaultRV32Config.fir@39764.4]
  wire  _T_206; // @[Misc.scala 214:29:freechips.rocketchip.system.DefaultRV32Config.fir@39765.4]
  wire  _T_216; // @[ToTL.scala 105:29:freechips.rocketchip.system.DefaultRV32Config.fir@39801.4]
  wire [1:0] _T_223; // @[OneHot.scala 65:12:freechips.rocketchip.system.DefaultRV32Config.fir@39814.4]
  reg [7:0] _T_433; // @[Arbiter.scala 78:30:freechips.rocketchip.system.DefaultRV32Config.fir@40125.4]
  wire  _T_434; // @[Arbiter.scala 79:28:freechips.rocketchip.system.DefaultRV32Config.fir@40126.4]
  wire  _T_348; // @[ToTL.scala 134:34:freechips.rocketchip.system.DefaultRV32Config.fir@39959.4]
  wire [1:0] _T_440; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@40132.4]
  reg [1:0] _T_446; // @[Arbiter.scala 22:23:freechips.rocketchip.system.DefaultRV32Config.fir@40142.4]
  wire [1:0] _T_447; // @[Arbiter.scala 23:30:freechips.rocketchip.system.DefaultRV32Config.fir@40143.4]
  wire [1:0] _T_448; // @[Arbiter.scala 23:28:freechips.rocketchip.system.DefaultRV32Config.fir@40144.4]
  wire [3:0] _T_449; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@40145.4]
  wire [3:0] _GEN_18; // @[package.scala 226:43:freechips.rocketchip.system.DefaultRV32Config.fir@40147.4]
  wire [3:0] _T_451; // @[package.scala 226:43:freechips.rocketchip.system.DefaultRV32Config.fir@40147.4]
  wire [3:0] _T_454; // @[Arbiter.scala 24:66:freechips.rocketchip.system.DefaultRV32Config.fir@40150.4]
  wire [3:0] _GEN_19; // @[Arbiter.scala 24:58:freechips.rocketchip.system.DefaultRV32Config.fir@40151.4]
  wire [3:0] _T_455; // @[Arbiter.scala 24:58:freechips.rocketchip.system.DefaultRV32Config.fir@40151.4]
  wire [1:0] _T_458; // @[Arbiter.scala 25:39:freechips.rocketchip.system.DefaultRV32Config.fir@40154.4]
  wire [1:0] _T_459; // @[Arbiter.scala 25:18:freechips.rocketchip.system.DefaultRV32Config.fir@40155.4]
  reg  _T_513_0; // @[Arbiter.scala 107:26:freechips.rocketchip.system.DefaultRV32Config.fir@40233.4]
  wire  _T_516_0; // @[Arbiter.scala 112:24:freechips.rocketchip.system.DefaultRV32Config.fir@40238.4]
  wire  _T_517; // @[Arbiter.scala 114:31:freechips.rocketchip.system.DefaultRV32Config.fir@40239.4]
  wire  _T_227; // @[Decoupled.scala 40:37:freechips.rocketchip.system.DefaultRV32Config.fir@39818.4]
  wire  _T_228; // @[ToTL.scala 115:28:freechips.rocketchip.system.DefaultRV32Config.fir@39819.4]
  wire [2:0] _T_230; // @[ToTL.scala 115:43:freechips.rocketchip.system.DefaultRV32Config.fir@39822.6]
  wire  _T_232; // @[ToTL.scala 115:28:freechips.rocketchip.system.DefaultRV32Config.fir@39826.4]
  wire [2:0] _T_234; // @[ToTL.scala 115:43:freechips.rocketchip.system.DefaultRV32Config.fir@39829.6]
  wire [15:0] _T_236; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@39834.4]
  wire [22:0] _GEN_20; // @[Bundles.scala 30:21:freechips.rocketchip.system.DefaultRV32Config.fir@39835.4]
  wire [22:0] _T_237; // @[Bundles.scala 30:21:freechips.rocketchip.system.DefaultRV32Config.fir@39835.4]
  wire [15:0] _T_239; // @[package.scala 205:35:freechips.rocketchip.system.DefaultRV32Config.fir@39837.4]
  wire [15:0] _T_240; // @[package.scala 205:40:freechips.rocketchip.system.DefaultRV32Config.fir@39838.4]
  wire [15:0] _T_241; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@39839.4]
  wire [15:0] _T_242; // @[package.scala 205:53:freechips.rocketchip.system.DefaultRV32Config.fir@39840.4]
  wire [15:0] _T_243; // @[package.scala 205:51:freechips.rocketchip.system.DefaultRV32Config.fir@39841.4]
  wire  _T_246; // @[OneHot.scala 32:14:freechips.rocketchip.system.DefaultRV32Config.fir@39844.4]
  wire [7:0] _T_247; // @[OneHot.scala 32:28:freechips.rocketchip.system.DefaultRV32Config.fir@39845.4]
  wire  _T_250; // @[OneHot.scala 32:14:freechips.rocketchip.system.DefaultRV32Config.fir@39848.4]
  wire [3:0] _T_251; // @[OneHot.scala 32:28:freechips.rocketchip.system.DefaultRV32Config.fir@39849.4]
  wire  _T_254; // @[OneHot.scala 32:14:freechips.rocketchip.system.DefaultRV32Config.fir@39852.4]
  wire [1:0] _T_255; // @[OneHot.scala 32:28:freechips.rocketchip.system.DefaultRV32Config.fir@39853.4]
  wire [3:0] _T_259; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@39857.4]
  wire  _T_261; // @[Parameters.scala 93:42:freechips.rocketchip.system.DefaultRV32Config.fir@39859.4]
  wire [31:0] _T_264; // @[Parameters.scala 137:31:freechips.rocketchip.system.DefaultRV32Config.fir@39862.4]
  wire [32:0] _T_265; // @[Parameters.scala 137:49:freechips.rocketchip.system.DefaultRV32Config.fir@39863.4]
  wire [32:0] _T_267; // @[Parameters.scala 137:52:freechips.rocketchip.system.DefaultRV32Config.fir@39865.4]
  wire  _T_268; // @[Parameters.scala 137:67:freechips.rocketchip.system.DefaultRV32Config.fir@39866.4]
  wire  _T_269; // @[Parameters.scala 551:56:freechips.rocketchip.system.DefaultRV32Config.fir@39867.4]
  wire  _T_271; // @[Parameters.scala 93:42:freechips.rocketchip.system.DefaultRV32Config.fir@39869.4]
  wire [32:0] _T_275; // @[Parameters.scala 137:49:freechips.rocketchip.system.DefaultRV32Config.fir@39873.4]
  wire [32:0] _T_277; // @[Parameters.scala 137:52:freechips.rocketchip.system.DefaultRV32Config.fir@39875.4]
  wire  _T_278; // @[Parameters.scala 137:67:freechips.rocketchip.system.DefaultRV32Config.fir@39876.4]
  wire [31:0] _T_279; // @[Parameters.scala 137:31:freechips.rocketchip.system.DefaultRV32Config.fir@39877.4]
  wire [32:0] _T_280; // @[Parameters.scala 137:49:freechips.rocketchip.system.DefaultRV32Config.fir@39878.4]
  wire [32:0] _T_282; // @[Parameters.scala 137:52:freechips.rocketchip.system.DefaultRV32Config.fir@39880.4]
  wire  _T_283; // @[Parameters.scala 137:67:freechips.rocketchip.system.DefaultRV32Config.fir@39881.4]
  wire [31:0] _T_284; // @[Parameters.scala 137:31:freechips.rocketchip.system.DefaultRV32Config.fir@39882.4]
  wire [32:0] _T_285; // @[Parameters.scala 137:49:freechips.rocketchip.system.DefaultRV32Config.fir@39883.4]
  wire [32:0] _T_287; // @[Parameters.scala 137:52:freechips.rocketchip.system.DefaultRV32Config.fir@39885.4]
  wire  _T_288; // @[Parameters.scala 137:67:freechips.rocketchip.system.DefaultRV32Config.fir@39886.4]
  wire [31:0] _T_289; // @[Parameters.scala 137:31:freechips.rocketchip.system.DefaultRV32Config.fir@39887.4]
  wire [32:0] _T_290; // @[Parameters.scala 137:49:freechips.rocketchip.system.DefaultRV32Config.fir@39888.4]
  wire [32:0] _T_292; // @[Parameters.scala 137:52:freechips.rocketchip.system.DefaultRV32Config.fir@39890.4]
  wire  _T_293; // @[Parameters.scala 137:67:freechips.rocketchip.system.DefaultRV32Config.fir@39891.4]
  wire  _T_294; // @[Parameters.scala 552:42:freechips.rocketchip.system.DefaultRV32Config.fir@39892.4]
  wire  _T_295; // @[Parameters.scala 552:42:freechips.rocketchip.system.DefaultRV32Config.fir@39893.4]
  wire  _T_296; // @[Parameters.scala 552:42:freechips.rocketchip.system.DefaultRV32Config.fir@39894.4]
  wire  _T_297; // @[Parameters.scala 551:56:freechips.rocketchip.system.DefaultRV32Config.fir@39895.4]
  wire  _T_306; // @[Parameters.scala 93:42:freechips.rocketchip.system.DefaultRV32Config.fir@39904.4]
  wire [31:0] _T_309; // @[Parameters.scala 137:31:freechips.rocketchip.system.DefaultRV32Config.fir@39907.4]
  wire [32:0] _T_310; // @[Parameters.scala 137:49:freechips.rocketchip.system.DefaultRV32Config.fir@39908.4]
  wire [32:0] _T_312; // @[Parameters.scala 137:52:freechips.rocketchip.system.DefaultRV32Config.fir@39910.4]
  wire  _T_313; // @[Parameters.scala 137:67:freechips.rocketchip.system.DefaultRV32Config.fir@39911.4]
  wire  _T_314; // @[Parameters.scala 551:56:freechips.rocketchip.system.DefaultRV32Config.fir@39912.4]
  wire  _T_316; // @[Parameters.scala 553:30:freechips.rocketchip.system.DefaultRV32Config.fir@39914.4]
  wire  _T_318; // @[Parameters.scala 553:30:freechips.rocketchip.system.DefaultRV32Config.fir@39916.4]
  wire [13:0] _GEN_21; // @[ToTL.scala 122:59:freechips.rocketchip.system.DefaultRV32Config.fir@39918.4]
  wire [13:0] _T_320; // @[ToTL.scala 122:59:freechips.rocketchip.system.DefaultRV32Config.fir@39918.4]
  wire [31:0] _T_321; // @[ToTL.scala 122:23:freechips.rocketchip.system.DefaultRV32Config.fir@39919.4]
  reg [2:0] _T_323_0; // @[ToTL.scala 123:28:freechips.rocketchip.system.DefaultRV32Config.fir@39924.4]
  reg [2:0] _T_323_1; // @[ToTL.scala 123:28:freechips.rocketchip.system.DefaultRV32Config.fir@39924.4]
  wire [2:0] _GEN_5; // @[ToTL.scala 127:50:freechips.rocketchip.system.DefaultRV32Config.fir@39925.4]
  wire  _T_327; // @[ToTL.scala 130:15:freechips.rocketchip.system.DefaultRV32Config.fir@39928.4]
  wire [29:0] _T_329; // @[package.scala 207:77:freechips.rocketchip.system.DefaultRV32Config.fir@39930.4]
  wire [14:0] _T_331; // @[package.scala 207:46:freechips.rocketchip.system.DefaultRV32Config.fir@39932.4]
  wire  _T_332; // @[ToTL.scala 130:39:freechips.rocketchip.system.DefaultRV32Config.fir@39933.4]
  wire  _T_333; // @[ToTL.scala 130:28:freechips.rocketchip.system.DefaultRV32Config.fir@39934.4]
  wire  _T_335; // @[ToTL.scala 130:14:freechips.rocketchip.system.DefaultRV32Config.fir@39936.4]
  wire  _T_336; // @[ToTL.scala 130:14:freechips.rocketchip.system.DefaultRV32Config.fir@39937.4]
  wire  _T_338; // @[ToTL.scala 131:46:freechips.rocketchip.system.DefaultRV32Config.fir@39943.4]
  wire  _T_339; // @[ToTL.scala 131:28:freechips.rocketchip.system.DefaultRV32Config.fir@39944.4]
  wire  _T_340; // @[ToTL.scala 131:77:freechips.rocketchip.system.DefaultRV32Config.fir@39945.4]
  wire  _T_341; // @[ToTL.scala 131:58:freechips.rocketchip.system.DefaultRV32Config.fir@39946.4]
  wire  _T_343; // @[ToTL.scala 131:14:freechips.rocketchip.system.DefaultRV32Config.fir@39948.4]
  wire  _T_344; // @[ToTL.scala 131:14:freechips.rocketchip.system.DefaultRV32Config.fir@39949.4]
  reg  _T_513_1; // @[Arbiter.scala 107:26:freechips.rocketchip.system.DefaultRV32Config.fir@40233.4]
  wire  _T_516_1; // @[Arbiter.scala 112:24:freechips.rocketchip.system.DefaultRV32Config.fir@40238.4]
  wire  _T_518; // @[Arbiter.scala 114:31:freechips.rocketchip.system.DefaultRV32Config.fir@40241.4]
  wire  _T_345; // @[ToTL.scala 132:34:freechips.rocketchip.system.DefaultRV32Config.fir@39954.4]
  wire  _T_346; // @[ToTL.scala 132:48:freechips.rocketchip.system.DefaultRV32Config.fir@39955.4]
  wire  _T_411; // @[ToTL.scala 141:29:freechips.rocketchip.system.DefaultRV32Config.fir@40055.4]
  wire [1:0] _T_418; // @[OneHot.scala 65:12:freechips.rocketchip.system.DefaultRV32Config.fir@40068.4]
  wire  _T_422; // @[Decoupled.scala 40:37:freechips.rocketchip.system.DefaultRV32Config.fir@40072.4]
  wire  _T_423; // @[ToTL.scala 151:28:freechips.rocketchip.system.DefaultRV32Config.fir@40073.4]
  wire [2:0] _T_425; // @[ToTL.scala 151:43:freechips.rocketchip.system.DefaultRV32Config.fir@40076.6]
  wire  _T_427; // @[ToTL.scala 151:28:freechips.rocketchip.system.DefaultRV32Config.fir@40080.4]
  wire [2:0] _T_429; // @[ToTL.scala 151:43:freechips.rocketchip.system.DefaultRV32Config.fir@40083.6]
  wire  _T_435; // @[Arbiter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@40127.4]
  wire  _T_460; // @[Arbiter.scala 26:27:freechips.rocketchip.system.DefaultRV32Config.fir@40156.4]
  wire  _T_461; // @[Arbiter.scala 26:18:freechips.rocketchip.system.DefaultRV32Config.fir@40157.4]
  wire [1:0] _T_462; // @[Arbiter.scala 27:29:freechips.rocketchip.system.DefaultRV32Config.fir@40159.6]
  wire [2:0] _T_463; // @[package.scala 217:48:freechips.rocketchip.system.DefaultRV32Config.fir@40160.6]
  wire [1:0] _T_465; // @[package.scala 217:43:freechips.rocketchip.system.DefaultRV32Config.fir@40162.6]
  wire  _T_471; // @[Arbiter.scala 88:79:freechips.rocketchip.system.DefaultRV32Config.fir@40172.4]
  wire  _T_472; // @[Arbiter.scala 88:79:freechips.rocketchip.system.DefaultRV32Config.fir@40173.4]
  wire  _T_478; // @[Arbiter.scala 95:53:freechips.rocketchip.system.DefaultRV32Config.fir@40183.4]
  wire  _T_480; // @[Arbiter.scala 96:67:freechips.rocketchip.system.DefaultRV32Config.fir@40185.4]
  wire  _T_483; // @[Arbiter.scala 96:67:freechips.rocketchip.system.DefaultRV32Config.fir@40188.4]
  wire  _T_484; // @[Arbiter.scala 96:64:freechips.rocketchip.system.DefaultRV32Config.fir@40189.4]
  wire  _T_487; // @[Arbiter.scala 96:13:freechips.rocketchip.system.DefaultRV32Config.fir@40192.4]
  wire  _T_488; // @[Arbiter.scala 96:13:freechips.rocketchip.system.DefaultRV32Config.fir@40193.4]
  wire  _T_489; // @[Arbiter.scala 98:36:freechips.rocketchip.system.DefaultRV32Config.fir@40198.4]
  wire  _T_490; // @[Arbiter.scala 98:15:freechips.rocketchip.system.DefaultRV32Config.fir@40199.4]
  wire  _T_492; // @[Arbiter.scala 98:41:freechips.rocketchip.system.DefaultRV32Config.fir@40201.4]
  wire  _T_494; // @[Arbiter.scala 98:14:freechips.rocketchip.system.DefaultRV32Config.fir@40203.4]
  wire  _T_495; // @[Arbiter.scala 98:14:freechips.rocketchip.system.DefaultRV32Config.fir@40204.4]
  wire  _T_499; // @[Arbiter.scala 99:41:freechips.rocketchip.system.DefaultRV32Config.fir@40212.4]
  wire  _T_501; // @[Arbiter.scala 99:14:freechips.rocketchip.system.DefaultRV32Config.fir@40214.4]
  wire  _T_502; // @[Arbiter.scala 99:14:freechips.rocketchip.system.DefaultRV32Config.fir@40215.4]
  wire  _T_514_0; // @[Arbiter.scala 108:30:freechips.rocketchip.system.DefaultRV32Config.fir@40234.4]
  wire  _T_514_1; // @[Arbiter.scala 108:30:freechips.rocketchip.system.DefaultRV32Config.fir@40234.4]
  wire  _T_520; // @[Mux.scala 27:72:freechips.rocketchip.system.DefaultRV32Config.fir@40244.4]
  wire  _T_521; // @[Mux.scala 27:72:freechips.rocketchip.system.DefaultRV32Config.fir@40245.4]
  wire  _T_522; // @[Mux.scala 27:72:freechips.rocketchip.system.DefaultRV32Config.fir@40246.4]
  wire  _T_524; // @[Arbiter.scala 116:29:freechips.rocketchip.system.DefaultRV32Config.fir@40249.4]
  wire  _T_508; // @[ReadyValidCancel.scala 52:33:freechips.rocketchip.system.DefaultRV32Config.fir@40225.4]
  wire [7:0] _GEN_22; // @[Arbiter.scala 104:52:freechips.rocketchip.system.DefaultRV32Config.fir@40226.4]
  wire [7:0] _T_510; // @[Arbiter.scala 104:52:freechips.rocketchip.system.DefaultRV32Config.fir@40227.4]
  wire [72:0] _T_530; // @[Mux.scala 27:72:freechips.rocketchip.system.DefaultRV32Config.fir@40258.4]
  wire [76:0] _T_534; // @[Mux.scala 27:72:freechips.rocketchip.system.DefaultRV32Config.fir@40262.4]
  wire [34:0] _T_537; // @[Mux.scala 27:72:freechips.rocketchip.system.DefaultRV32Config.fir@40265.4]
  wire [125:0] _T_542; // @[Mux.scala 27:72:freechips.rocketchip.system.DefaultRV32Config.fir@40270.4]
  wire [125:0] _T_543; // @[Mux.scala 27:72:freechips.rocketchip.system.DefaultRV32Config.fir@40271.4]
  wire [76:0] _T_549; // @[Mux.scala 27:72:freechips.rocketchip.system.DefaultRV32Config.fir@40277.4]
  wire [34:0] _T_552; // @[Mux.scala 27:72:freechips.rocketchip.system.DefaultRV32Config.fir@40280.4]
  wire [125:0] _T_557; // @[Mux.scala 27:72:freechips.rocketchip.system.DefaultRV32Config.fir@40285.4]
  wire [125:0] _T_558; // @[Mux.scala 27:72:freechips.rocketchip.system.DefaultRV32Config.fir@40286.4]
  wire [125:0] _T_559; // @[Mux.scala 27:72:freechips.rocketchip.system.DefaultRV32Config.fir@40287.4]
  wire  _T_582; // @[ToTL.scala 159:42:freechips.rocketchip.system.DefaultRV32Config.fir@40377.4]
  wire  _T_581_ready; // @[ToTL.scala 157:23:freechips.rocketchip.system.DefaultRV32Config.fir@40375.4 Decoupled.scala 290:17:freechips.rocketchip.system.DefaultRV32Config.fir@40422.4]
  wire  _T_580_ready; // @[ToTL.scala 156:23:freechips.rocketchip.system.DefaultRV32Config.fir@40373.4 Decoupled.scala 290:17:freechips.rocketchip.system.DefaultRV32Config.fir@40445.4]
  wire  _T_604; // @[ToTL.scala 163:25:freechips.rocketchip.system.DefaultRV32Config.fir@40402.4]
  wire  _T_585; // @[Decoupled.scala 40:37:freechips.rocketchip.system.DefaultRV32Config.fir@40380.4]
  wire [26:0] _T_587; // @[package.scala 207:77:freechips.rocketchip.system.DefaultRV32Config.fir@40382.4]
  wire [11:0] _T_589; // @[package.scala 207:46:freechips.rocketchip.system.DefaultRV32Config.fir@40384.4]
  wire [8:0] _T_592; // @[Edges.scala 222:14:freechips.rocketchip.system.DefaultRV32Config.fir@40387.4]
  reg [8:0] _T_593; // @[Edges.scala 230:27:freechips.rocketchip.system.DefaultRV32Config.fir@40388.4]
  wire [8:0] _T_595; // @[Edges.scala 231:28:freechips.rocketchip.system.DefaultRV32Config.fir@40390.4]
  wire  _T_596; // @[Edges.scala 232:25:freechips.rocketchip.system.DefaultRV32Config.fir@40391.4]
  wire  _T_597; // @[Edges.scala 233:25:freechips.rocketchip.system.DefaultRV32Config.fir@40392.4]
  wire  _T_598; // @[Edges.scala 233:47:freechips.rocketchip.system.DefaultRV32Config.fir@40393.4]
  wire  _T_606; // @[ToTL.scala 165:36:freechips.rocketchip.system.DefaultRV32Config.fir@40406.4]
  reg [2:0] _T_613_0; // @[ToTL.scala 185:28:freechips.rocketchip.system.DefaultRV32Config.fir@40455.4]
  reg [2:0] _T_613_1; // @[ToTL.scala 185:28:freechips.rocketchip.system.DefaultRV32Config.fir@40455.4]
  wire  _T_611_bits_id; // @[Decoupled.scala 308:19:freechips.rocketchip.system.DefaultRV32Config.fir@40446.4 Decoupled.scala 309:14:freechips.rocketchip.system.DefaultRV32Config.fir@40448.4]
  wire [2:0] _GEN_11; // @[ToTL.scala 186:43:freechips.rocketchip.system.DefaultRV32Config.fir@40456.4]
  wire [2:0] _GEN_13; // @[ToTL.scala 186:43:freechips.rocketchip.system.DefaultRV32Config.fir@40456.4]
  wire  _T_614; // @[ToTL.scala 186:43:freechips.rocketchip.system.DefaultRV32Config.fir@40456.4]
  wire [1:0] _T_616; // @[OneHot.scala 65:12:freechips.rocketchip.system.DefaultRV32Config.fir@40458.4]
  wire  _T_611_valid; // @[Decoupled.scala 308:19:freechips.rocketchip.system.DefaultRV32Config.fir@40446.4 Decoupled.scala 310:15:freechips.rocketchip.system.DefaultRV32Config.fir@40449.4]
  wire  _T_628; // @[ToTL.scala 194:31:freechips.rocketchip.system.DefaultRV32Config.fir@40478.4]
  wire  _T_620; // @[Decoupled.scala 40:37:freechips.rocketchip.system.DefaultRV32Config.fir@40462.4]
  wire  _T_621; // @[ToTL.scala 190:27:freechips.rocketchip.system.DefaultRV32Config.fir@40463.4]
  wire [2:0] _T_623; // @[ToTL.scala 190:42:freechips.rocketchip.system.DefaultRV32Config.fir@40466.6]
  wire  _T_625; // @[ToTL.scala 190:27:freechips.rocketchip.system.DefaultRV32Config.fir@40470.4]
  wire [2:0] _T_627; // @[ToTL.scala 190:42:freechips.rocketchip.system.DefaultRV32Config.fir@40473.6]
  Queue_16 Queue ( // @[Decoupled.scala 287:21:freechips.rocketchip.system.DefaultRV32Config.fir@40414.4]
    .clock(Queue_clock),
    .reset(Queue_reset),
    .io_enq_ready(Queue_io_enq_ready),
    .io_enq_valid(Queue_io_enq_valid),
    .io_enq_bits_id(Queue_io_enq_bits_id),
    .io_enq_bits_data(Queue_io_enq_bits_data),
    .io_enq_bits_resp(Queue_io_enq_bits_resp),
    .io_enq_bits_last(Queue_io_enq_bits_last),
    .io_deq_ready(Queue_io_deq_ready),
    .io_deq_valid(Queue_io_deq_valid),
    .io_deq_bits_id(Queue_io_deq_bits_id),
    .io_deq_bits_data(Queue_io_deq_bits_data),
    .io_deq_bits_resp(Queue_io_deq_bits_resp),
    .io_deq_bits_last(Queue_io_deq_bits_last)
  );
  Queue_17 Queue_1 ( // @[Decoupled.scala 287:21:freechips.rocketchip.system.DefaultRV32Config.fir@40439.4]
    .clock(Queue_1_clock),
    .reset(Queue_1_reset),
    .io_enq_ready(Queue_1_io_enq_ready),
    .io_enq_valid(Queue_1_io_enq_valid),
    .io_enq_bits_id(Queue_1_io_enq_bits_id),
    .io_enq_bits_resp(Queue_1_io_enq_bits_resp),
    .io_deq_ready(Queue_1_io_deq_ready),
    .io_deq_valid(Queue_1_io_deq_valid),
    .io_deq_bits_id(Queue_1_io_deq_bits_id),
    .io_deq_bits_resp(Queue_1_io_deq_bits_resp)
  );
  assign _T_3 = {auto_in_ar_bits_len,8'hff}; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@39547.4]
  assign _GEN_16 = {{7'd0}, _T_3}; // @[Bundles.scala 30:21:freechips.rocketchip.system.DefaultRV32Config.fir@39548.4]
  assign _T_4 = _GEN_16 << auto_in_ar_bits_size; // @[Bundles.scala 30:21:freechips.rocketchip.system.DefaultRV32Config.fir@39548.4]
  assign _T_6 = {_T_4[22:8], 1'h0}; // @[package.scala 205:35:freechips.rocketchip.system.DefaultRV32Config.fir@39550.4]
  assign _T_7 = _T_6 | 16'h1; // @[package.scala 205:40:freechips.rocketchip.system.DefaultRV32Config.fir@39551.4]
  assign _T_8 = {1'h0,_T_4[22:8]}; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@39552.4]
  assign _T_9 = ~_T_8; // @[package.scala 205:53:freechips.rocketchip.system.DefaultRV32Config.fir@39553.4]
  assign _T_10 = _T_7 & _T_9; // @[package.scala 205:51:freechips.rocketchip.system.DefaultRV32Config.fir@39554.4]
  assign _T_13 = |_T_10[15:8]; // @[OneHot.scala 32:14:freechips.rocketchip.system.DefaultRV32Config.fir@39557.4]
  assign _T_14 = _T_10[15:8] | _T_10[7:0]; // @[OneHot.scala 32:28:freechips.rocketchip.system.DefaultRV32Config.fir@39558.4]
  assign _T_17 = |_T_14[7:4]; // @[OneHot.scala 32:14:freechips.rocketchip.system.DefaultRV32Config.fir@39561.4]
  assign _T_18 = _T_14[7:4] | _T_14[3:0]; // @[OneHot.scala 32:28:freechips.rocketchip.system.DefaultRV32Config.fir@39562.4]
  assign _T_21 = |_T_18[3:2]; // @[OneHot.scala 32:14:freechips.rocketchip.system.DefaultRV32Config.fir@39565.4]
  assign _T_22 = _T_18[3:2] | _T_18[1:0]; // @[OneHot.scala 32:28:freechips.rocketchip.system.DefaultRV32Config.fir@39566.4]
  assign _T_26 = {_T_13,_T_17,_T_21,_T_22[1]}; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@39570.4]
  assign _T_28 = _T_26 <= 4'hc; // @[Parameters.scala 93:42:freechips.rocketchip.system.DefaultRV32Config.fir@39572.4]
  assign _T_31 = auto_in_ar_bits_addr ^ 32'h3000; // @[Parameters.scala 137:31:freechips.rocketchip.system.DefaultRV32Config.fir@39575.4]
  assign _T_32 = {1'b0,$signed(_T_31)}; // @[Parameters.scala 137:49:freechips.rocketchip.system.DefaultRV32Config.fir@39576.4]
  assign _T_34 = $signed(_T_32) & -33'sh1000; // @[Parameters.scala 137:52:freechips.rocketchip.system.DefaultRV32Config.fir@39578.4]
  assign _T_35 = $signed(_T_34) == 33'sh0; // @[Parameters.scala 137:67:freechips.rocketchip.system.DefaultRV32Config.fir@39579.4]
  assign _T_36 = _T_28 & _T_35; // @[Parameters.scala 551:56:freechips.rocketchip.system.DefaultRV32Config.fir@39580.4]
  assign _T_38 = _T_26 <= 4'h6; // @[Parameters.scala 93:42:freechips.rocketchip.system.DefaultRV32Config.fir@39582.4]
  assign _T_42 = {1'b0,$signed(auto_in_ar_bits_addr)}; // @[Parameters.scala 137:49:freechips.rocketchip.system.DefaultRV32Config.fir@39586.4]
  assign _T_44 = $signed(_T_42) & -33'sh1000; // @[Parameters.scala 137:52:freechips.rocketchip.system.DefaultRV32Config.fir@39588.4]
  assign _T_45 = $signed(_T_44) == 33'sh0; // @[Parameters.scala 137:67:freechips.rocketchip.system.DefaultRV32Config.fir@39589.4]
  assign _T_46 = auto_in_ar_bits_addr ^ 32'h10000; // @[Parameters.scala 137:31:freechips.rocketchip.system.DefaultRV32Config.fir@39590.4]
  assign _T_47 = {1'b0,$signed(_T_46)}; // @[Parameters.scala 137:49:freechips.rocketchip.system.DefaultRV32Config.fir@39591.4]
  assign _T_49 = $signed(_T_47) & -33'sh10000; // @[Parameters.scala 137:52:freechips.rocketchip.system.DefaultRV32Config.fir@39593.4]
  assign _T_50 = $signed(_T_49) == 33'sh0; // @[Parameters.scala 137:67:freechips.rocketchip.system.DefaultRV32Config.fir@39594.4]
  assign _T_51 = auto_in_ar_bits_addr ^ 32'h2000000; // @[Parameters.scala 137:31:freechips.rocketchip.system.DefaultRV32Config.fir@39595.4]
  assign _T_52 = {1'b0,$signed(_T_51)}; // @[Parameters.scala 137:49:freechips.rocketchip.system.DefaultRV32Config.fir@39596.4]
  assign _T_54 = $signed(_T_52) & -33'sh10000; // @[Parameters.scala 137:52:freechips.rocketchip.system.DefaultRV32Config.fir@39598.4]
  assign _T_55 = $signed(_T_54) == 33'sh0; // @[Parameters.scala 137:67:freechips.rocketchip.system.DefaultRV32Config.fir@39599.4]
  assign _T_56 = auto_in_ar_bits_addr ^ 32'hc000000; // @[Parameters.scala 137:31:freechips.rocketchip.system.DefaultRV32Config.fir@39600.4]
  assign _T_57 = {1'b0,$signed(_T_56)}; // @[Parameters.scala 137:49:freechips.rocketchip.system.DefaultRV32Config.fir@39601.4]
  assign _T_59 = $signed(_T_57) & -33'sh4000000; // @[Parameters.scala 137:52:freechips.rocketchip.system.DefaultRV32Config.fir@39603.4]
  assign _T_60 = $signed(_T_59) == 33'sh0; // @[Parameters.scala 137:67:freechips.rocketchip.system.DefaultRV32Config.fir@39604.4]
  assign _T_61 = auto_in_ar_bits_addr ^ 32'h60000000; // @[Parameters.scala 137:31:freechips.rocketchip.system.DefaultRV32Config.fir@39605.4]
  assign _T_62 = {1'b0,$signed(_T_61)}; // @[Parameters.scala 137:49:freechips.rocketchip.system.DefaultRV32Config.fir@39606.4]
  assign _T_64 = $signed(_T_62) & -33'sh20000000; // @[Parameters.scala 137:52:freechips.rocketchip.system.DefaultRV32Config.fir@39608.4]
  assign _T_65 = $signed(_T_64) == 33'sh0; // @[Parameters.scala 137:67:freechips.rocketchip.system.DefaultRV32Config.fir@39609.4]
  assign _T_66 = auto_in_ar_bits_addr ^ 32'h80000000; // @[Parameters.scala 137:31:freechips.rocketchip.system.DefaultRV32Config.fir@39610.4]
  assign _T_67 = {1'b0,$signed(_T_66)}; // @[Parameters.scala 137:49:freechips.rocketchip.system.DefaultRV32Config.fir@39611.4]
  assign _T_69 = $signed(_T_67) & -33'sh10000000; // @[Parameters.scala 137:52:freechips.rocketchip.system.DefaultRV32Config.fir@39613.4]
  assign _T_70 = $signed(_T_69) == 33'sh0; // @[Parameters.scala 137:67:freechips.rocketchip.system.DefaultRV32Config.fir@39614.4]
  assign _T_71 = _T_45 | _T_50; // @[Parameters.scala 552:42:freechips.rocketchip.system.DefaultRV32Config.fir@39615.4]
  assign _T_72 = _T_71 | _T_55; // @[Parameters.scala 552:42:freechips.rocketchip.system.DefaultRV32Config.fir@39616.4]
  assign _T_73 = _T_72 | _T_60; // @[Parameters.scala 552:42:freechips.rocketchip.system.DefaultRV32Config.fir@39617.4]
  assign _T_74 = _T_73 | _T_65; // @[Parameters.scala 552:42:freechips.rocketchip.system.DefaultRV32Config.fir@39618.4]
  assign _T_75 = _T_74 | _T_70; // @[Parameters.scala 552:42:freechips.rocketchip.system.DefaultRV32Config.fir@39619.4]
  assign _T_76 = _T_38 & _T_75; // @[Parameters.scala 551:56:freechips.rocketchip.system.DefaultRV32Config.fir@39620.4]
  assign _T_78 = _T_36 | _T_76; // @[Parameters.scala 553:30:freechips.rocketchip.system.DefaultRV32Config.fir@39622.4]
  assign _GEN_17 = {{11'd0}, auto_in_ar_bits_addr[2:0]}; // @[ToTL.scala 89:59:freechips.rocketchip.system.DefaultRV32Config.fir@39624.4]
  assign _T_80 = 14'h3000 | _GEN_17; // @[ToTL.scala 89:59:freechips.rocketchip.system.DefaultRV32Config.fir@39624.4]
  assign _T_81 = _T_78 ? auto_in_ar_bits_addr : {{18'd0}, _T_80}; // @[ToTL.scala 89:23:freechips.rocketchip.system.DefaultRV32Config.fir@39625.4]
  assign _GEN_1 = auto_in_ar_bits_id ? _T_83_1 : _T_83_0; // @[ToTL.scala 94:50:freechips.rocketchip.system.DefaultRV32Config.fir@39631.4]
  assign _T_87 = ~auto_in_ar_valid; // @[ToTL.scala 97:15:freechips.rocketchip.system.DefaultRV32Config.fir@39634.4]
  assign _T_89 = 30'h7fff << _T_26; // @[package.scala 207:77:freechips.rocketchip.system.DefaultRV32Config.fir@39636.4]
  assign _T_91 = ~_T_89[14:0]; // @[package.scala 207:46:freechips.rocketchip.system.DefaultRV32Config.fir@39638.4]
  assign _T_92 = _T_4[22:8] == _T_91; // @[ToTL.scala 97:39:freechips.rocketchip.system.DefaultRV32Config.fir@39639.4]
  assign _T_93 = _T_87 | _T_92; // @[ToTL.scala 97:28:freechips.rocketchip.system.DefaultRV32Config.fir@39640.4]
  assign _T_95 = _T_93 | reset; // @[ToTL.scala 97:14:freechips.rocketchip.system.DefaultRV32Config.fir@39642.4]
  assign _T_96 = ~_T_95; // @[ToTL.scala 97:14:freechips.rocketchip.system.DefaultRV32Config.fir@39643.4]
  assign _T_152 = 4'h1 << _T_26[1:0]; // @[OneHot.scala 65:12:freechips.rocketchip.system.DefaultRV32Config.fir@39711.4]
  assign _T_154 = _T_152[2:0] | 3'h1; // @[Misc.scala 201:81:freechips.rocketchip.system.DefaultRV32Config.fir@39713.4]
  assign _T_155 = _T_26 >= 4'h3; // @[Misc.scala 205:21:freechips.rocketchip.system.DefaultRV32Config.fir@39714.4]
  assign _T_158 = ~_T_81[2]; // @[Misc.scala 210:20:freechips.rocketchip.system.DefaultRV32Config.fir@39717.4]
  assign _T_160 = _T_154[2] & _T_158; // @[Misc.scala 214:38:freechips.rocketchip.system.DefaultRV32Config.fir@39719.4]
  assign _T_161 = _T_155 | _T_160; // @[Misc.scala 214:29:freechips.rocketchip.system.DefaultRV32Config.fir@39720.4]
  assign _T_163 = _T_154[2] & _T_81[2]; // @[Misc.scala 214:38:freechips.rocketchip.system.DefaultRV32Config.fir@39722.4]
  assign _T_164 = _T_155 | _T_163; // @[Misc.scala 214:29:freechips.rocketchip.system.DefaultRV32Config.fir@39723.4]
  assign _T_167 = ~_T_81[1]; // @[Misc.scala 210:20:freechips.rocketchip.system.DefaultRV32Config.fir@39726.4]
  assign _T_168 = _T_158 & _T_167; // @[Misc.scala 213:27:freechips.rocketchip.system.DefaultRV32Config.fir@39727.4]
  assign _T_169 = _T_154[1] & _T_168; // @[Misc.scala 214:38:freechips.rocketchip.system.DefaultRV32Config.fir@39728.4]
  assign _T_170 = _T_161 | _T_169; // @[Misc.scala 214:29:freechips.rocketchip.system.DefaultRV32Config.fir@39729.4]
  assign _T_171 = _T_158 & _T_81[1]; // @[Misc.scala 213:27:freechips.rocketchip.system.DefaultRV32Config.fir@39730.4]
  assign _T_172 = _T_154[1] & _T_171; // @[Misc.scala 214:38:freechips.rocketchip.system.DefaultRV32Config.fir@39731.4]
  assign _T_173 = _T_161 | _T_172; // @[Misc.scala 214:29:freechips.rocketchip.system.DefaultRV32Config.fir@39732.4]
  assign _T_174 = _T_81[2] & _T_167; // @[Misc.scala 213:27:freechips.rocketchip.system.DefaultRV32Config.fir@39733.4]
  assign _T_175 = _T_154[1] & _T_174; // @[Misc.scala 214:38:freechips.rocketchip.system.DefaultRV32Config.fir@39734.4]
  assign _T_176 = _T_164 | _T_175; // @[Misc.scala 214:29:freechips.rocketchip.system.DefaultRV32Config.fir@39735.4]
  assign _T_177 = _T_81[2] & _T_81[1]; // @[Misc.scala 213:27:freechips.rocketchip.system.DefaultRV32Config.fir@39736.4]
  assign _T_178 = _T_154[1] & _T_177; // @[Misc.scala 214:38:freechips.rocketchip.system.DefaultRV32Config.fir@39737.4]
  assign _T_179 = _T_164 | _T_178; // @[Misc.scala 214:29:freechips.rocketchip.system.DefaultRV32Config.fir@39738.4]
  assign _T_182 = ~_T_81[0]; // @[Misc.scala 210:20:freechips.rocketchip.system.DefaultRV32Config.fir@39741.4]
  assign _T_183 = _T_168 & _T_182; // @[Misc.scala 213:27:freechips.rocketchip.system.DefaultRV32Config.fir@39742.4]
  assign _T_184 = _T_154[0] & _T_183; // @[Misc.scala 214:38:freechips.rocketchip.system.DefaultRV32Config.fir@39743.4]
  assign _T_185 = _T_170 | _T_184; // @[Misc.scala 214:29:freechips.rocketchip.system.DefaultRV32Config.fir@39744.4]
  assign _T_186 = _T_168 & _T_81[0]; // @[Misc.scala 213:27:freechips.rocketchip.system.DefaultRV32Config.fir@39745.4]
  assign _T_187 = _T_154[0] & _T_186; // @[Misc.scala 214:38:freechips.rocketchip.system.DefaultRV32Config.fir@39746.4]
  assign _T_188 = _T_170 | _T_187; // @[Misc.scala 214:29:freechips.rocketchip.system.DefaultRV32Config.fir@39747.4]
  assign _T_189 = _T_171 & _T_182; // @[Misc.scala 213:27:freechips.rocketchip.system.DefaultRV32Config.fir@39748.4]
  assign _T_190 = _T_154[0] & _T_189; // @[Misc.scala 214:38:freechips.rocketchip.system.DefaultRV32Config.fir@39749.4]
  assign _T_191 = _T_173 | _T_190; // @[Misc.scala 214:29:freechips.rocketchip.system.DefaultRV32Config.fir@39750.4]
  assign _T_192 = _T_171 & _T_81[0]; // @[Misc.scala 213:27:freechips.rocketchip.system.DefaultRV32Config.fir@39751.4]
  assign _T_193 = _T_154[0] & _T_192; // @[Misc.scala 214:38:freechips.rocketchip.system.DefaultRV32Config.fir@39752.4]
  assign _T_194 = _T_173 | _T_193; // @[Misc.scala 214:29:freechips.rocketchip.system.DefaultRV32Config.fir@39753.4]
  assign _T_195 = _T_174 & _T_182; // @[Misc.scala 213:27:freechips.rocketchip.system.DefaultRV32Config.fir@39754.4]
  assign _T_196 = _T_154[0] & _T_195; // @[Misc.scala 214:38:freechips.rocketchip.system.DefaultRV32Config.fir@39755.4]
  assign _T_197 = _T_176 | _T_196; // @[Misc.scala 214:29:freechips.rocketchip.system.DefaultRV32Config.fir@39756.4]
  assign _T_198 = _T_174 & _T_81[0]; // @[Misc.scala 213:27:freechips.rocketchip.system.DefaultRV32Config.fir@39757.4]
  assign _T_199 = _T_154[0] & _T_198; // @[Misc.scala 214:38:freechips.rocketchip.system.DefaultRV32Config.fir@39758.4]
  assign _T_200 = _T_176 | _T_199; // @[Misc.scala 214:29:freechips.rocketchip.system.DefaultRV32Config.fir@39759.4]
  assign _T_201 = _T_177 & _T_182; // @[Misc.scala 213:27:freechips.rocketchip.system.DefaultRV32Config.fir@39760.4]
  assign _T_202 = _T_154[0] & _T_201; // @[Misc.scala 214:38:freechips.rocketchip.system.DefaultRV32Config.fir@39761.4]
  assign _T_203 = _T_179 | _T_202; // @[Misc.scala 214:29:freechips.rocketchip.system.DefaultRV32Config.fir@39762.4]
  assign _T_204 = _T_177 & _T_81[0]; // @[Misc.scala 213:27:freechips.rocketchip.system.DefaultRV32Config.fir@39763.4]
  assign _T_205 = _T_154[0] & _T_204; // @[Misc.scala 214:38:freechips.rocketchip.system.DefaultRV32Config.fir@39764.4]
  assign _T_206 = _T_179 | _T_205; // @[Misc.scala 214:29:freechips.rocketchip.system.DefaultRV32Config.fir@39765.4]
  assign _T_216 = ~auto_in_ar_bits_prot[1]; // @[ToTL.scala 105:29:freechips.rocketchip.system.DefaultRV32Config.fir@39801.4]
  assign _T_223 = 2'h1 << auto_in_ar_bits_id; // @[OneHot.scala 65:12:freechips.rocketchip.system.DefaultRV32Config.fir@39814.4]
  assign _T_434 = _T_433 == 8'h0; // @[Arbiter.scala 79:28:freechips.rocketchip.system.DefaultRV32Config.fir@40126.4]
  assign _T_348 = auto_in_aw_valid & auto_in_w_valid; // @[ToTL.scala 134:34:freechips.rocketchip.system.DefaultRV32Config.fir@39959.4]
  assign _T_440 = {_T_348,auto_in_ar_valid}; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@40132.4]
  assign _T_447 = ~_T_446; // @[Arbiter.scala 23:30:freechips.rocketchip.system.DefaultRV32Config.fir@40143.4]
  assign _T_448 = _T_440 & _T_447; // @[Arbiter.scala 23:28:freechips.rocketchip.system.DefaultRV32Config.fir@40144.4]
  assign _T_449 = {_T_448,_T_348,auto_in_ar_valid}; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@40145.4]
  assign _GEN_18 = {{1'd0}, _T_449[3:1]}; // @[package.scala 226:43:freechips.rocketchip.system.DefaultRV32Config.fir@40147.4]
  assign _T_451 = _T_449 | _GEN_18; // @[package.scala 226:43:freechips.rocketchip.system.DefaultRV32Config.fir@40147.4]
  assign _T_454 = {_T_446, 2'h0}; // @[Arbiter.scala 24:66:freechips.rocketchip.system.DefaultRV32Config.fir@40150.4]
  assign _GEN_19 = {{1'd0}, _T_451[3:1]}; // @[Arbiter.scala 24:58:freechips.rocketchip.system.DefaultRV32Config.fir@40151.4]
  assign _T_455 = _GEN_19 | _T_454; // @[Arbiter.scala 24:58:freechips.rocketchip.system.DefaultRV32Config.fir@40151.4]
  assign _T_458 = _T_455[3:2] & _T_455[1:0]; // @[Arbiter.scala 25:39:freechips.rocketchip.system.DefaultRV32Config.fir@40154.4]
  assign _T_459 = ~_T_458; // @[Arbiter.scala 25:18:freechips.rocketchip.system.DefaultRV32Config.fir@40155.4]
  assign _T_516_0 = _T_434 ? _T_459[0] : _T_513_0; // @[Arbiter.scala 112:24:freechips.rocketchip.system.DefaultRV32Config.fir@40238.4]
  assign _T_517 = auto_out_a_ready & _T_516_0; // @[Arbiter.scala 114:31:freechips.rocketchip.system.DefaultRV32Config.fir@40239.4]
  assign _T_227 = _T_517 & auto_in_ar_valid; // @[Decoupled.scala 40:37:freechips.rocketchip.system.DefaultRV32Config.fir@39818.4]
  assign _T_228 = _T_227 & _T_223[0]; // @[ToTL.scala 115:28:freechips.rocketchip.system.DefaultRV32Config.fir@39819.4]
  assign _T_230 = _T_83_0 + 3'h1; // @[ToTL.scala 115:43:freechips.rocketchip.system.DefaultRV32Config.fir@39822.6]
  assign _T_232 = _T_227 & _T_223[1]; // @[ToTL.scala 115:28:freechips.rocketchip.system.DefaultRV32Config.fir@39826.4]
  assign _T_234 = _T_83_1 + 3'h1; // @[ToTL.scala 115:43:freechips.rocketchip.system.DefaultRV32Config.fir@39829.6]
  assign _T_236 = {auto_in_aw_bits_len,8'hff}; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@39834.4]
  assign _GEN_20 = {{7'd0}, _T_236}; // @[Bundles.scala 30:21:freechips.rocketchip.system.DefaultRV32Config.fir@39835.4]
  assign _T_237 = _GEN_20 << auto_in_aw_bits_size; // @[Bundles.scala 30:21:freechips.rocketchip.system.DefaultRV32Config.fir@39835.4]
  assign _T_239 = {_T_237[22:8], 1'h0}; // @[package.scala 205:35:freechips.rocketchip.system.DefaultRV32Config.fir@39837.4]
  assign _T_240 = _T_239 | 16'h1; // @[package.scala 205:40:freechips.rocketchip.system.DefaultRV32Config.fir@39838.4]
  assign _T_241 = {1'h0,_T_237[22:8]}; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@39839.4]
  assign _T_242 = ~_T_241; // @[package.scala 205:53:freechips.rocketchip.system.DefaultRV32Config.fir@39840.4]
  assign _T_243 = _T_240 & _T_242; // @[package.scala 205:51:freechips.rocketchip.system.DefaultRV32Config.fir@39841.4]
  assign _T_246 = |_T_243[15:8]; // @[OneHot.scala 32:14:freechips.rocketchip.system.DefaultRV32Config.fir@39844.4]
  assign _T_247 = _T_243[15:8] | _T_243[7:0]; // @[OneHot.scala 32:28:freechips.rocketchip.system.DefaultRV32Config.fir@39845.4]
  assign _T_250 = |_T_247[7:4]; // @[OneHot.scala 32:14:freechips.rocketchip.system.DefaultRV32Config.fir@39848.4]
  assign _T_251 = _T_247[7:4] | _T_247[3:0]; // @[OneHot.scala 32:28:freechips.rocketchip.system.DefaultRV32Config.fir@39849.4]
  assign _T_254 = |_T_251[3:2]; // @[OneHot.scala 32:14:freechips.rocketchip.system.DefaultRV32Config.fir@39852.4]
  assign _T_255 = _T_251[3:2] | _T_251[1:0]; // @[OneHot.scala 32:28:freechips.rocketchip.system.DefaultRV32Config.fir@39853.4]
  assign _T_259 = {_T_246,_T_250,_T_254,_T_255[1]}; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@39857.4]
  assign _T_261 = _T_259 <= 4'hc; // @[Parameters.scala 93:42:freechips.rocketchip.system.DefaultRV32Config.fir@39859.4]
  assign _T_264 = auto_in_aw_bits_addr ^ 32'h3000; // @[Parameters.scala 137:31:freechips.rocketchip.system.DefaultRV32Config.fir@39862.4]
  assign _T_265 = {1'b0,$signed(_T_264)}; // @[Parameters.scala 137:49:freechips.rocketchip.system.DefaultRV32Config.fir@39863.4]
  assign _T_267 = $signed(_T_265) & -33'sh1000; // @[Parameters.scala 137:52:freechips.rocketchip.system.DefaultRV32Config.fir@39865.4]
  assign _T_268 = $signed(_T_267) == 33'sh0; // @[Parameters.scala 137:67:freechips.rocketchip.system.DefaultRV32Config.fir@39866.4]
  assign _T_269 = _T_261 & _T_268; // @[Parameters.scala 551:56:freechips.rocketchip.system.DefaultRV32Config.fir@39867.4]
  assign _T_271 = _T_259 <= 4'h6; // @[Parameters.scala 93:42:freechips.rocketchip.system.DefaultRV32Config.fir@39869.4]
  assign _T_275 = {1'b0,$signed(auto_in_aw_bits_addr)}; // @[Parameters.scala 137:49:freechips.rocketchip.system.DefaultRV32Config.fir@39873.4]
  assign _T_277 = $signed(_T_275) & -33'sh1000; // @[Parameters.scala 137:52:freechips.rocketchip.system.DefaultRV32Config.fir@39875.4]
  assign _T_278 = $signed(_T_277) == 33'sh0; // @[Parameters.scala 137:67:freechips.rocketchip.system.DefaultRV32Config.fir@39876.4]
  assign _T_279 = auto_in_aw_bits_addr ^ 32'h2000000; // @[Parameters.scala 137:31:freechips.rocketchip.system.DefaultRV32Config.fir@39877.4]
  assign _T_280 = {1'b0,$signed(_T_279)}; // @[Parameters.scala 137:49:freechips.rocketchip.system.DefaultRV32Config.fir@39878.4]
  assign _T_282 = $signed(_T_280) & -33'sh10000; // @[Parameters.scala 137:52:freechips.rocketchip.system.DefaultRV32Config.fir@39880.4]
  assign _T_283 = $signed(_T_282) == 33'sh0; // @[Parameters.scala 137:67:freechips.rocketchip.system.DefaultRV32Config.fir@39881.4]
  assign _T_284 = auto_in_aw_bits_addr ^ 32'hc000000; // @[Parameters.scala 137:31:freechips.rocketchip.system.DefaultRV32Config.fir@39882.4]
  assign _T_285 = {1'b0,$signed(_T_284)}; // @[Parameters.scala 137:49:freechips.rocketchip.system.DefaultRV32Config.fir@39883.4]
  assign _T_287 = $signed(_T_285) & -33'sh4000000; // @[Parameters.scala 137:52:freechips.rocketchip.system.DefaultRV32Config.fir@39885.4]
  assign _T_288 = $signed(_T_287) == 33'sh0; // @[Parameters.scala 137:67:freechips.rocketchip.system.DefaultRV32Config.fir@39886.4]
  assign _T_289 = auto_in_aw_bits_addr ^ 32'h80000000; // @[Parameters.scala 137:31:freechips.rocketchip.system.DefaultRV32Config.fir@39887.4]
  assign _T_290 = {1'b0,$signed(_T_289)}; // @[Parameters.scala 137:49:freechips.rocketchip.system.DefaultRV32Config.fir@39888.4]
  assign _T_292 = $signed(_T_290) & -33'sh10000000; // @[Parameters.scala 137:52:freechips.rocketchip.system.DefaultRV32Config.fir@39890.4]
  assign _T_293 = $signed(_T_292) == 33'sh0; // @[Parameters.scala 137:67:freechips.rocketchip.system.DefaultRV32Config.fir@39891.4]
  assign _T_294 = _T_278 | _T_283; // @[Parameters.scala 552:42:freechips.rocketchip.system.DefaultRV32Config.fir@39892.4]
  assign _T_295 = _T_294 | _T_288; // @[Parameters.scala 552:42:freechips.rocketchip.system.DefaultRV32Config.fir@39893.4]
  assign _T_296 = _T_295 | _T_293; // @[Parameters.scala 552:42:freechips.rocketchip.system.DefaultRV32Config.fir@39894.4]
  assign _T_297 = _T_271 & _T_296; // @[Parameters.scala 551:56:freechips.rocketchip.system.DefaultRV32Config.fir@39895.4]
  assign _T_306 = _T_259 <= 4'h8; // @[Parameters.scala 93:42:freechips.rocketchip.system.DefaultRV32Config.fir@39904.4]
  assign _T_309 = auto_in_aw_bits_addr ^ 32'h60000000; // @[Parameters.scala 137:31:freechips.rocketchip.system.DefaultRV32Config.fir@39907.4]
  assign _T_310 = {1'b0,$signed(_T_309)}; // @[Parameters.scala 137:49:freechips.rocketchip.system.DefaultRV32Config.fir@39908.4]
  assign _T_312 = $signed(_T_310) & -33'sh20000000; // @[Parameters.scala 137:52:freechips.rocketchip.system.DefaultRV32Config.fir@39910.4]
  assign _T_313 = $signed(_T_312) == 33'sh0; // @[Parameters.scala 137:67:freechips.rocketchip.system.DefaultRV32Config.fir@39911.4]
  assign _T_314 = _T_306 & _T_313; // @[Parameters.scala 551:56:freechips.rocketchip.system.DefaultRV32Config.fir@39912.4]
  assign _T_316 = _T_269 | _T_297; // @[Parameters.scala 553:30:freechips.rocketchip.system.DefaultRV32Config.fir@39914.4]
  assign _T_318 = _T_316 | _T_314; // @[Parameters.scala 553:30:freechips.rocketchip.system.DefaultRV32Config.fir@39916.4]
  assign _GEN_21 = {{11'd0}, auto_in_aw_bits_addr[2:0]}; // @[ToTL.scala 122:59:freechips.rocketchip.system.DefaultRV32Config.fir@39918.4]
  assign _T_320 = 14'h3000 | _GEN_21; // @[ToTL.scala 122:59:freechips.rocketchip.system.DefaultRV32Config.fir@39918.4]
  assign _T_321 = _T_318 ? auto_in_aw_bits_addr : {{18'd0}, _T_320}; // @[ToTL.scala 122:23:freechips.rocketchip.system.DefaultRV32Config.fir@39919.4]
  assign _GEN_5 = auto_in_aw_bits_id ? _T_323_1 : _T_323_0; // @[ToTL.scala 127:50:freechips.rocketchip.system.DefaultRV32Config.fir@39925.4]
  assign _T_327 = ~auto_in_aw_valid; // @[ToTL.scala 130:15:freechips.rocketchip.system.DefaultRV32Config.fir@39928.4]
  assign _T_329 = 30'h7fff << _T_259; // @[package.scala 207:77:freechips.rocketchip.system.DefaultRV32Config.fir@39930.4]
  assign _T_331 = ~_T_329[14:0]; // @[package.scala 207:46:freechips.rocketchip.system.DefaultRV32Config.fir@39932.4]
  assign _T_332 = _T_237[22:8] == _T_331; // @[ToTL.scala 130:39:freechips.rocketchip.system.DefaultRV32Config.fir@39933.4]
  assign _T_333 = _T_327 | _T_332; // @[ToTL.scala 130:28:freechips.rocketchip.system.DefaultRV32Config.fir@39934.4]
  assign _T_335 = _T_333 | reset; // @[ToTL.scala 130:14:freechips.rocketchip.system.DefaultRV32Config.fir@39936.4]
  assign _T_336 = ~_T_335; // @[ToTL.scala 130:14:freechips.rocketchip.system.DefaultRV32Config.fir@39937.4]
  assign _T_338 = auto_in_aw_bits_len == 8'h0; // @[ToTL.scala 131:46:freechips.rocketchip.system.DefaultRV32Config.fir@39943.4]
  assign _T_339 = _T_327 | _T_338; // @[ToTL.scala 131:28:freechips.rocketchip.system.DefaultRV32Config.fir@39944.4]
  assign _T_340 = auto_in_aw_bits_size == 3'h3; // @[ToTL.scala 131:77:freechips.rocketchip.system.DefaultRV32Config.fir@39945.4]
  assign _T_341 = _T_339 | _T_340; // @[ToTL.scala 131:58:freechips.rocketchip.system.DefaultRV32Config.fir@39946.4]
  assign _T_343 = _T_341 | reset; // @[ToTL.scala 131:14:freechips.rocketchip.system.DefaultRV32Config.fir@39948.4]
  assign _T_344 = ~_T_343; // @[ToTL.scala 131:14:freechips.rocketchip.system.DefaultRV32Config.fir@39949.4]
  assign _T_516_1 = _T_434 ? _T_459[1] : _T_513_1; // @[Arbiter.scala 112:24:freechips.rocketchip.system.DefaultRV32Config.fir@40238.4]
  assign _T_518 = auto_out_a_ready & _T_516_1; // @[Arbiter.scala 114:31:freechips.rocketchip.system.DefaultRV32Config.fir@40241.4]
  assign _T_345 = _T_518 & auto_in_w_valid; // @[ToTL.scala 132:34:freechips.rocketchip.system.DefaultRV32Config.fir@39954.4]
  assign _T_346 = _T_345 & auto_in_w_bits_last; // @[ToTL.scala 132:48:freechips.rocketchip.system.DefaultRV32Config.fir@39955.4]
  assign _T_411 = ~auto_in_aw_bits_prot[1]; // @[ToTL.scala 141:29:freechips.rocketchip.system.DefaultRV32Config.fir@40055.4]
  assign _T_418 = 2'h1 << auto_in_aw_bits_id; // @[OneHot.scala 65:12:freechips.rocketchip.system.DefaultRV32Config.fir@40068.4]
  assign _T_422 = _T_346 & auto_in_aw_valid; // @[Decoupled.scala 40:37:freechips.rocketchip.system.DefaultRV32Config.fir@40072.4]
  assign _T_423 = _T_422 & _T_418[0]; // @[ToTL.scala 151:28:freechips.rocketchip.system.DefaultRV32Config.fir@40073.4]
  assign _T_425 = _T_323_0 + 3'h1; // @[ToTL.scala 151:43:freechips.rocketchip.system.DefaultRV32Config.fir@40076.6]
  assign _T_427 = _T_422 & _T_418[1]; // @[ToTL.scala 151:28:freechips.rocketchip.system.DefaultRV32Config.fir@40080.4]
  assign _T_429 = _T_323_1 + 3'h1; // @[ToTL.scala 151:43:freechips.rocketchip.system.DefaultRV32Config.fir@40083.6]
  assign _T_435 = _T_434 & auto_out_a_ready; // @[Arbiter.scala 80:24:freechips.rocketchip.system.DefaultRV32Config.fir@40127.4]
  assign _T_460 = |_T_440; // @[Arbiter.scala 26:27:freechips.rocketchip.system.DefaultRV32Config.fir@40156.4]
  assign _T_461 = _T_435 & _T_460; // @[Arbiter.scala 26:18:freechips.rocketchip.system.DefaultRV32Config.fir@40157.4]
  assign _T_462 = _T_459 & _T_440; // @[Arbiter.scala 27:29:freechips.rocketchip.system.DefaultRV32Config.fir@40159.6]
  assign _T_463 = {_T_462, 1'h0}; // @[package.scala 217:48:freechips.rocketchip.system.DefaultRV32Config.fir@40160.6]
  assign _T_465 = _T_462 | _T_463[1:0]; // @[package.scala 217:43:freechips.rocketchip.system.DefaultRV32Config.fir@40162.6]
  assign _T_471 = _T_459[0] & auto_in_ar_valid; // @[Arbiter.scala 88:79:freechips.rocketchip.system.DefaultRV32Config.fir@40172.4]
  assign _T_472 = _T_459[1] & _T_348; // @[Arbiter.scala 88:79:freechips.rocketchip.system.DefaultRV32Config.fir@40173.4]
  assign _T_478 = _T_471 | _T_472; // @[Arbiter.scala 95:53:freechips.rocketchip.system.DefaultRV32Config.fir@40183.4]
  assign _T_480 = ~_T_471; // @[Arbiter.scala 96:67:freechips.rocketchip.system.DefaultRV32Config.fir@40185.4]
  assign _T_483 = ~_T_472; // @[Arbiter.scala 96:67:freechips.rocketchip.system.DefaultRV32Config.fir@40188.4]
  assign _T_484 = _T_480 | _T_483; // @[Arbiter.scala 96:64:freechips.rocketchip.system.DefaultRV32Config.fir@40189.4]
  assign _T_487 = _T_484 | reset; // @[Arbiter.scala 96:13:freechips.rocketchip.system.DefaultRV32Config.fir@40192.4]
  assign _T_488 = ~_T_487; // @[Arbiter.scala 96:13:freechips.rocketchip.system.DefaultRV32Config.fir@40193.4]
  assign _T_489 = auto_in_ar_valid | _T_348; // @[Arbiter.scala 98:36:freechips.rocketchip.system.DefaultRV32Config.fir@40198.4]
  assign _T_490 = ~_T_489; // @[Arbiter.scala 98:15:freechips.rocketchip.system.DefaultRV32Config.fir@40199.4]
  assign _T_492 = _T_490 | _T_478; // @[Arbiter.scala 98:41:freechips.rocketchip.system.DefaultRV32Config.fir@40201.4]
  assign _T_494 = _T_492 | reset; // @[Arbiter.scala 98:14:freechips.rocketchip.system.DefaultRV32Config.fir@40203.4]
  assign _T_495 = ~_T_494; // @[Arbiter.scala 98:14:freechips.rocketchip.system.DefaultRV32Config.fir@40204.4]
  assign _T_499 = _T_490 | _T_489; // @[Arbiter.scala 99:41:freechips.rocketchip.system.DefaultRV32Config.fir@40212.4]
  assign _T_501 = _T_499 | reset; // @[Arbiter.scala 99:14:freechips.rocketchip.system.DefaultRV32Config.fir@40214.4]
  assign _T_502 = ~_T_501; // @[Arbiter.scala 99:14:freechips.rocketchip.system.DefaultRV32Config.fir@40215.4]
  assign _T_514_0 = _T_434 ? _T_471 : _T_513_0; // @[Arbiter.scala 108:30:freechips.rocketchip.system.DefaultRV32Config.fir@40234.4]
  assign _T_514_1 = _T_434 ? _T_472 : _T_513_1; // @[Arbiter.scala 108:30:freechips.rocketchip.system.DefaultRV32Config.fir@40234.4]
  assign _T_520 = _T_513_0 & auto_in_ar_valid; // @[Mux.scala 27:72:freechips.rocketchip.system.DefaultRV32Config.fir@40244.4]
  assign _T_521 = _T_513_1 & _T_348; // @[Mux.scala 27:72:freechips.rocketchip.system.DefaultRV32Config.fir@40245.4]
  assign _T_522 = _T_520 | _T_521; // @[Mux.scala 27:72:freechips.rocketchip.system.DefaultRV32Config.fir@40246.4]
  assign _T_524 = _T_434 ? _T_489 : _T_522; // @[Arbiter.scala 116:29:freechips.rocketchip.system.DefaultRV32Config.fir@40249.4]
  assign _T_508 = auto_out_a_ready & _T_524; // @[ReadyValidCancel.scala 52:33:freechips.rocketchip.system.DefaultRV32Config.fir@40225.4]
  assign _GEN_22 = {{7'd0}, _T_508}; // @[Arbiter.scala 104:52:freechips.rocketchip.system.DefaultRV32Config.fir@40226.4]
  assign _T_510 = _T_433 - _GEN_22; // @[Arbiter.scala 104:52:freechips.rocketchip.system.DefaultRV32Config.fir@40227.4]
  assign _T_530 = {_T_206,_T_203,_T_200,_T_197,_T_194,_T_191,_T_188,_T_185,64'h0,1'h0}; // @[Mux.scala 27:72:freechips.rocketchip.system.DefaultRV32Config.fir@40258.4]
  assign _T_534 = {auto_in_ar_bits_cache[3],auto_in_ar_bits_prot[0],_T_216,auto_in_ar_bits_prot[2],_T_530}; // @[Mux.scala 27:72:freechips.rocketchip.system.DefaultRV32Config.fir@40262.4]
  assign _T_537 = {_T_81,auto_in_ar_bits_cache[0],auto_in_ar_bits_cache[1],auto_in_ar_bits_cache[2]}; // @[Mux.scala 27:72:freechips.rocketchip.system.DefaultRV32Config.fir@40265.4]
  assign _T_542 = {6'h20,_T_13,_T_17,_T_21,_T_22[1],auto_in_ar_bits_id,_GEN_1[1:0],1'h0,_T_537,_T_534}; // @[Mux.scala 27:72:freechips.rocketchip.system.DefaultRV32Config.fir@40270.4]
  assign _T_543 = _T_514_0 ? _T_542 : 126'h0; // @[Mux.scala 27:72:freechips.rocketchip.system.DefaultRV32Config.fir@40271.4]
  assign _T_549 = {auto_in_aw_bits_cache[3],auto_in_aw_bits_prot[0],_T_411,auto_in_aw_bits_prot[2],auto_in_w_bits_strb,auto_in_w_bits_data,1'h0}; // @[Mux.scala 27:72:freechips.rocketchip.system.DefaultRV32Config.fir@40277.4]
  assign _T_552 = {_T_321,auto_in_aw_bits_cache[0],auto_in_aw_bits_cache[1],auto_in_aw_bits_cache[2]}; // @[Mux.scala 27:72:freechips.rocketchip.system.DefaultRV32Config.fir@40280.4]
  assign _T_557 = {6'h8,_T_246,_T_250,_T_254,_T_255[1],auto_in_aw_bits_id,_GEN_5[1:0],1'h1,_T_552,_T_549}; // @[Mux.scala 27:72:freechips.rocketchip.system.DefaultRV32Config.fir@40285.4]
  assign _T_558 = _T_514_1 ? _T_557 : 126'h0; // @[Mux.scala 27:72:freechips.rocketchip.system.DefaultRV32Config.fir@40286.4]
  assign _T_559 = _T_543 | _T_558; // @[Mux.scala 27:72:freechips.rocketchip.system.DefaultRV32Config.fir@40287.4]
  assign _T_582 = auto_out_d_bits_denied | auto_out_d_bits_corrupt; // @[ToTL.scala 159:42:freechips.rocketchip.system.DefaultRV32Config.fir@40377.4]
  assign _T_581_ready = Queue_io_enq_ready; // @[ToTL.scala 157:23:freechips.rocketchip.system.DefaultRV32Config.fir@40375.4 Decoupled.scala 290:17:freechips.rocketchip.system.DefaultRV32Config.fir@40422.4]
  assign _T_580_ready = Queue_1_io_enq_ready; // @[ToTL.scala 156:23:freechips.rocketchip.system.DefaultRV32Config.fir@40373.4 Decoupled.scala 290:17:freechips.rocketchip.system.DefaultRV32Config.fir@40445.4]
  assign _T_604 = auto_out_d_bits_opcode[0] ? _T_581_ready : _T_580_ready; // @[ToTL.scala 163:25:freechips.rocketchip.system.DefaultRV32Config.fir@40402.4]
  assign _T_585 = _T_604 & auto_out_d_valid; // @[Decoupled.scala 40:37:freechips.rocketchip.system.DefaultRV32Config.fir@40380.4]
  assign _T_587 = 27'hfff << auto_out_d_bits_size; // @[package.scala 207:77:freechips.rocketchip.system.DefaultRV32Config.fir@40382.4]
  assign _T_589 = ~_T_587[11:0]; // @[package.scala 207:46:freechips.rocketchip.system.DefaultRV32Config.fir@40384.4]
  assign _T_592 = auto_out_d_bits_opcode[0] ? _T_589[11:3] : 9'h0; // @[Edges.scala 222:14:freechips.rocketchip.system.DefaultRV32Config.fir@40387.4]
  assign _T_595 = _T_593 - 9'h1; // @[Edges.scala 231:28:freechips.rocketchip.system.DefaultRV32Config.fir@40390.4]
  assign _T_596 = _T_593 == 9'h0; // @[Edges.scala 232:25:freechips.rocketchip.system.DefaultRV32Config.fir@40391.4]
  assign _T_597 = _T_593 == 9'h1; // @[Edges.scala 233:25:freechips.rocketchip.system.DefaultRV32Config.fir@40392.4]
  assign _T_598 = _T_592 == 9'h0; // @[Edges.scala 233:47:freechips.rocketchip.system.DefaultRV32Config.fir@40393.4]
  assign _T_606 = ~auto_out_d_bits_opcode[0]; // @[ToTL.scala 165:36:freechips.rocketchip.system.DefaultRV32Config.fir@40406.4]
  assign _T_611_bits_id = Queue_1_io_deq_bits_id; // @[Decoupled.scala 308:19:freechips.rocketchip.system.DefaultRV32Config.fir@40446.4 Decoupled.scala 309:14:freechips.rocketchip.system.DefaultRV32Config.fir@40448.4]
  assign _GEN_11 = _T_611_bits_id ? _T_613_1 : _T_613_0; // @[ToTL.scala 186:43:freechips.rocketchip.system.DefaultRV32Config.fir@40456.4]
  assign _GEN_13 = _T_611_bits_id ? _T_323_1 : _T_323_0; // @[ToTL.scala 186:43:freechips.rocketchip.system.DefaultRV32Config.fir@40456.4]
  assign _T_614 = _GEN_11 != _GEN_13; // @[ToTL.scala 186:43:freechips.rocketchip.system.DefaultRV32Config.fir@40456.4]
  assign _T_616 = 2'h1 << _T_611_bits_id; // @[OneHot.scala 65:12:freechips.rocketchip.system.DefaultRV32Config.fir@40458.4]
  assign _T_611_valid = Queue_1_io_deq_valid; // @[Decoupled.scala 308:19:freechips.rocketchip.system.DefaultRV32Config.fir@40446.4 Decoupled.scala 310:15:freechips.rocketchip.system.DefaultRV32Config.fir@40449.4]
  assign _T_628 = _T_611_valid & _T_614; // @[ToTL.scala 194:31:freechips.rocketchip.system.DefaultRV32Config.fir@40478.4]
  assign _T_620 = auto_in_b_ready & _T_628; // @[Decoupled.scala 40:37:freechips.rocketchip.system.DefaultRV32Config.fir@40462.4]
  assign _T_621 = _T_620 & _T_616[0]; // @[ToTL.scala 190:27:freechips.rocketchip.system.DefaultRV32Config.fir@40463.4]
  assign _T_623 = _T_613_0 + 3'h1; // @[ToTL.scala 190:42:freechips.rocketchip.system.DefaultRV32Config.fir@40466.6]
  assign _T_625 = _T_620 & _T_616[1]; // @[ToTL.scala 190:27:freechips.rocketchip.system.DefaultRV32Config.fir@40470.4]
  assign _T_627 = _T_613_1 + 3'h1; // @[ToTL.scala 190:42:freechips.rocketchip.system.DefaultRV32Config.fir@40473.6]
  assign auto_in_aw_ready = _T_345 & auto_in_w_bits_last; // @[LazyModule.scala 303:16:freechips.rocketchip.system.DefaultRV32Config.fir@39544.4]
  assign auto_in_w_ready = _T_518 & auto_in_aw_valid; // @[LazyModule.scala 303:16:freechips.rocketchip.system.DefaultRV32Config.fir@39544.4]
  assign auto_in_b_valid = _T_611_valid & _T_614; // @[LazyModule.scala 303:16:freechips.rocketchip.system.DefaultRV32Config.fir@39544.4]
  assign auto_in_b_bits_id = Queue_1_io_deq_bits_id; // @[LazyModule.scala 303:16:freechips.rocketchip.system.DefaultRV32Config.fir@39544.4]
  assign auto_in_b_bits_resp = Queue_1_io_deq_bits_resp; // @[LazyModule.scala 303:16:freechips.rocketchip.system.DefaultRV32Config.fir@39544.4]
  assign auto_in_ar_ready = auto_out_a_ready & _T_516_0; // @[LazyModule.scala 303:16:freechips.rocketchip.system.DefaultRV32Config.fir@39544.4]
  assign auto_in_r_valid = Queue_io_deq_valid; // @[LazyModule.scala 303:16:freechips.rocketchip.system.DefaultRV32Config.fir@39544.4]
  assign auto_in_r_bits_id = Queue_io_deq_bits_id; // @[LazyModule.scala 303:16:freechips.rocketchip.system.DefaultRV32Config.fir@39544.4]
  assign auto_in_r_bits_data = Queue_io_deq_bits_data; // @[LazyModule.scala 303:16:freechips.rocketchip.system.DefaultRV32Config.fir@39544.4]
  assign auto_in_r_bits_resp = Queue_io_deq_bits_resp; // @[LazyModule.scala 303:16:freechips.rocketchip.system.DefaultRV32Config.fir@39544.4]
  assign auto_in_r_bits_last = Queue_io_deq_bits_last; // @[LazyModule.scala 303:16:freechips.rocketchip.system.DefaultRV32Config.fir@39544.4]
  assign auto_out_a_valid = _T_434 ? _T_489 : _T_522; // @[LazyModule.scala 305:12:freechips.rocketchip.system.DefaultRV32Config.fir@39543.4]
  assign auto_out_a_bits_opcode = _T_559[125:123]; // @[LazyModule.scala 305:12:freechips.rocketchip.system.DefaultRV32Config.fir@39543.4]
  assign auto_out_a_bits_param = _T_559[122:120]; // @[LazyModule.scala 305:12:freechips.rocketchip.system.DefaultRV32Config.fir@39543.4]
  assign auto_out_a_bits_size = _T_559[119:116]; // @[LazyModule.scala 305:12:freechips.rocketchip.system.DefaultRV32Config.fir@39543.4]
  assign auto_out_a_bits_source = _T_559[115:112]; // @[LazyModule.scala 305:12:freechips.rocketchip.system.DefaultRV32Config.fir@39543.4]
  assign auto_out_a_bits_address = _T_559[111:80]; // @[LazyModule.scala 305:12:freechips.rocketchip.system.DefaultRV32Config.fir@39543.4]
  assign auto_out_a_bits_user_amba_prot_bufferable = _T_559[79]; // @[LazyModule.scala 305:12:freechips.rocketchip.system.DefaultRV32Config.fir@39543.4]
  assign auto_out_a_bits_user_amba_prot_modifiable = _T_559[78]; // @[LazyModule.scala 305:12:freechips.rocketchip.system.DefaultRV32Config.fir@39543.4]
  assign auto_out_a_bits_user_amba_prot_readalloc = _T_559[77]; // @[LazyModule.scala 305:12:freechips.rocketchip.system.DefaultRV32Config.fir@39543.4]
  assign auto_out_a_bits_user_amba_prot_writealloc = _T_559[76]; // @[LazyModule.scala 305:12:freechips.rocketchip.system.DefaultRV32Config.fir@39543.4]
  assign auto_out_a_bits_user_amba_prot_privileged = _T_559[75]; // @[LazyModule.scala 305:12:freechips.rocketchip.system.DefaultRV32Config.fir@39543.4]
  assign auto_out_a_bits_user_amba_prot_secure = _T_559[74]; // @[LazyModule.scala 305:12:freechips.rocketchip.system.DefaultRV32Config.fir@39543.4]
  assign auto_out_a_bits_user_amba_prot_fetch = _T_559[73]; // @[LazyModule.scala 305:12:freechips.rocketchip.system.DefaultRV32Config.fir@39543.4]
  assign auto_out_a_bits_mask = _T_559[72:65]; // @[LazyModule.scala 305:12:freechips.rocketchip.system.DefaultRV32Config.fir@39543.4]
  assign auto_out_a_bits_data = _T_559[64:1]; // @[LazyModule.scala 305:12:freechips.rocketchip.system.DefaultRV32Config.fir@39543.4]
  assign auto_out_a_bits_corrupt = _T_559[0]; // @[LazyModule.scala 305:12:freechips.rocketchip.system.DefaultRV32Config.fir@39543.4]
  assign auto_out_d_ready = auto_out_d_bits_opcode[0] ? _T_581_ready : _T_580_ready; // @[LazyModule.scala 305:12:freechips.rocketchip.system.DefaultRV32Config.fir@39543.4]
  assign Queue_clock = clock; // @[:freechips.rocketchip.system.DefaultRV32Config.fir@40415.4]
  assign Queue_reset = reset; // @[:freechips.rocketchip.system.DefaultRV32Config.fir@40416.4]
  assign Queue_io_enq_valid = auto_out_d_valid & auto_out_d_bits_opcode[0]; // @[Decoupled.scala 288:22:freechips.rocketchip.system.DefaultRV32Config.fir@40417.4]
  assign Queue_io_enq_bits_id = auto_out_d_bits_source[3]; // @[Decoupled.scala 289:21:freechips.rocketchip.system.DefaultRV32Config.fir@40421.4]
  assign Queue_io_enq_bits_data = auto_out_d_bits_data; // @[Decoupled.scala 289:21:freechips.rocketchip.system.DefaultRV32Config.fir@40420.4]
  assign Queue_io_enq_bits_resp = _T_582 ? 2'h2 : 2'h0; // @[Decoupled.scala 289:21:freechips.rocketchip.system.DefaultRV32Config.fir@40419.4]
  assign Queue_io_enq_bits_last = _T_597 | _T_598; // @[Decoupled.scala 289:21:freechips.rocketchip.system.DefaultRV32Config.fir@40418.4]
  assign Queue_io_deq_ready = auto_in_r_ready; // @[Decoupled.scala 311:15:freechips.rocketchip.system.DefaultRV32Config.fir@40429.4]
  assign Queue_1_clock = clock; // @[:freechips.rocketchip.system.DefaultRV32Config.fir@40440.4]
  assign Queue_1_reset = reset; // @[:freechips.rocketchip.system.DefaultRV32Config.fir@40441.4]
  assign Queue_1_io_enq_valid = auto_out_d_valid & _T_606; // @[Decoupled.scala 288:22:freechips.rocketchip.system.DefaultRV32Config.fir@40442.4]
  assign Queue_1_io_enq_bits_id = auto_out_d_bits_source[3]; // @[Decoupled.scala 289:21:freechips.rocketchip.system.DefaultRV32Config.fir@40444.4]
  assign Queue_1_io_enq_bits_resp = _T_582 ? 2'h2 : 2'h0; // @[Decoupled.scala 289:21:freechips.rocketchip.system.DefaultRV32Config.fir@40443.4]
  assign Queue_1_io_deq_ready = auto_in_b_ready & _T_614; // @[Decoupled.scala 311:15:freechips.rocketchip.system.DefaultRV32Config.fir@40450.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_83_0 = _RAND_0[2:0];
  _RAND_1 = {1{`RANDOM}};
  _T_83_1 = _RAND_1[2:0];
  _RAND_2 = {1{`RANDOM}};
  _T_433 = _RAND_2[7:0];
  _RAND_3 = {1{`RANDOM}};
  _T_446 = _RAND_3[1:0];
  _RAND_4 = {1{`RANDOM}};
  _T_513_0 = _RAND_4[0:0];
  _RAND_5 = {1{`RANDOM}};
  _T_323_0 = _RAND_5[2:0];
  _RAND_6 = {1{`RANDOM}};
  _T_323_1 = _RAND_6[2:0];
  _RAND_7 = {1{`RANDOM}};
  _T_513_1 = _RAND_7[0:0];
  _RAND_8 = {1{`RANDOM}};
  _T_593 = _RAND_8[8:0];
  _RAND_9 = {1{`RANDOM}};
  _T_613_0 = _RAND_9[2:0];
  _RAND_10 = {1{`RANDOM}};
  _T_613_1 = _RAND_10[2:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      _T_83_0 <= 3'h0;
    end else if (_T_228) begin
      _T_83_0 <= _T_230;
    end
    if (reset) begin
      _T_83_1 <= 3'h0;
    end else if (_T_232) begin
      _T_83_1 <= _T_234;
    end
    if (reset) begin
      _T_433 <= 8'h0;
    end else if (_T_435) begin
      if (_T_472) begin
        _T_433 <= auto_in_aw_bits_len;
      end else begin
        _T_433 <= 8'h0;
      end
    end else begin
      _T_433 <= _T_510;
    end
    if (reset) begin
      _T_446 <= 2'h3;
    end else if (_T_461) begin
      _T_446 <= _T_465;
    end
    if (reset) begin
      _T_513_0 <= 1'h0;
    end else if (_T_434) begin
      _T_513_0 <= _T_471;
    end
    if (reset) begin
      _T_323_0 <= 3'h0;
    end else if (_T_423) begin
      _T_323_0 <= _T_425;
    end
    if (reset) begin
      _T_323_1 <= 3'h0;
    end else if (_T_427) begin
      _T_323_1 <= _T_429;
    end
    if (reset) begin
      _T_513_1 <= 1'h0;
    end else if (_T_434) begin
      _T_513_1 <= _T_472;
    end
    if (reset) begin
      _T_593 <= 9'h0;
    end else if (_T_585) begin
      if (_T_596) begin
        if (auto_out_d_bits_opcode[0]) begin
          _T_593 <= _T_589[11:3];
        end else begin
          _T_593 <= 9'h0;
        end
      end else begin
        _T_593 <= _T_595;
      end
    end
    if (reset) begin
      _T_613_0 <= 3'h0;
    end else if (_T_621) begin
      _T_613_0 <= _T_623;
    end
    if (reset) begin
      _T_613_1 <= 3'h0;
    end else if (_T_625) begin
      _T_613_1 <= _T_627;
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_96) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToTL.scala:97 assert (!in.ar.valid || r_size1 === UIntToOH1(r_size, beatCountBits)) // because aligned\n"); // @[ToTL.scala 97:14:freechips.rocketchip.system.DefaultRV32Config.fir@39645.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_96) begin
          $fatal; // @[ToTL.scala 97:14:freechips.rocketchip.system.DefaultRV32Config.fir@39646.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_336) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToTL.scala:130 assert (!in.aw.valid || w_size1 === UIntToOH1(w_size, beatCountBits)) // because aligned\n"); // @[ToTL.scala 130:14:freechips.rocketchip.system.DefaultRV32Config.fir@39939.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_336) begin
          $fatal; // @[ToTL.scala 130:14:freechips.rocketchip.system.DefaultRV32Config.fir@39940.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_344) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToTL.scala:131 assert (!in.aw.valid || in.aw.bits.len === UInt(0) || in.aw.bits.size === UInt(log2Ceil(beatBytes))) // because aligned\n"); // @[ToTL.scala 131:14:freechips.rocketchip.system.DefaultRV32Config.fir@39951.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_344) begin
          $fatal; // @[ToTL.scala 131:14:freechips.rocketchip.system.DefaultRV32Config.fir@39952.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_488) begin
          $fwrite(32'h80000002,"Assertion failed\n    at Arbiter.scala:96 assert((prefixOR zip earlyWinner) map { case (p,w) => !p || !w } reduce {_ && _})\n"); // @[Arbiter.scala 96:13:freechips.rocketchip.system.DefaultRV32Config.fir@40195.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_488) begin
          $fatal; // @[Arbiter.scala 96:13:freechips.rocketchip.system.DefaultRV32Config.fir@40196.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_495) begin
          $fwrite(32'h80000002,"Assertion failed\n    at Arbiter.scala:98 assert (!earlyValids.reduce(_||_) || earlyWinner.reduce(_||_))\n"); // @[Arbiter.scala 98:14:freechips.rocketchip.system.DefaultRV32Config.fir@40206.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_495) begin
          $fatal; // @[Arbiter.scala 98:14:freechips.rocketchip.system.DefaultRV32Config.fir@40207.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_502) begin
          $fwrite(32'h80000002,"Assertion failed\n    at Arbiter.scala:99 assert (!validQuals .reduce(_||_) || validQuals .reduce(_||_))\n"); // @[Arbiter.scala 99:14:freechips.rocketchip.system.DefaultRV32Config.fir@40217.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_502) begin
          $fatal; // @[Arbiter.scala 99:14:freechips.rocketchip.system.DefaultRV32Config.fir@40218.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
  end
endmodule
