module AXI4UserYanker_2( // @[:freechips.rocketchip.system.DefaultRV32Config.fir@71894.2]
  input         clock, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@71895.4]
  input         reset, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@71896.4]
  output        auto_in_aw_ready, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@71897.4]
  input         auto_in_aw_valid, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@71897.4]
  input  [3:0]  auto_in_aw_bits_id, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@71897.4]
  input  [31:0] auto_in_aw_bits_addr, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@71897.4]
  input  [7:0]  auto_in_aw_bits_len, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@71897.4]
  input  [2:0]  auto_in_aw_bits_size, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@71897.4]
  input  [1:0]  auto_in_aw_bits_burst, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@71897.4]
  input         auto_in_aw_bits_lock, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@71897.4]
  input  [3:0]  auto_in_aw_bits_cache, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@71897.4]
  input  [2:0]  auto_in_aw_bits_prot, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@71897.4]
  input  [3:0]  auto_in_aw_bits_qos, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@71897.4]
  input  [3:0]  auto_in_aw_bits_echo_tl_state_size, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@71897.4]
  input  [1:0]  auto_in_aw_bits_echo_tl_state_source, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@71897.4]
  output        auto_in_w_ready, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@71897.4]
  input         auto_in_w_valid, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@71897.4]
  input  [31:0] auto_in_w_bits_data, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@71897.4]
  input  [3:0]  auto_in_w_bits_strb, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@71897.4]
  input         auto_in_w_bits_last, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@71897.4]
  input         auto_in_b_ready, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@71897.4]
  output        auto_in_b_valid, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@71897.4]
  output [3:0]  auto_in_b_bits_id, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@71897.4]
  output [1:0]  auto_in_b_bits_resp, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@71897.4]
  output [3:0]  auto_in_b_bits_echo_tl_state_size, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@71897.4]
  output [1:0]  auto_in_b_bits_echo_tl_state_source, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@71897.4]
  output        auto_in_ar_ready, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@71897.4]
  input         auto_in_ar_valid, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@71897.4]
  input  [3:0]  auto_in_ar_bits_id, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@71897.4]
  input  [31:0] auto_in_ar_bits_addr, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@71897.4]
  input  [7:0]  auto_in_ar_bits_len, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@71897.4]
  input  [2:0]  auto_in_ar_bits_size, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@71897.4]
  input  [1:0]  auto_in_ar_bits_burst, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@71897.4]
  input         auto_in_ar_bits_lock, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@71897.4]
  input  [3:0]  auto_in_ar_bits_cache, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@71897.4]
  input  [2:0]  auto_in_ar_bits_prot, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@71897.4]
  input  [3:0]  auto_in_ar_bits_qos, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@71897.4]
  input  [3:0]  auto_in_ar_bits_echo_tl_state_size, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@71897.4]
  input  [1:0]  auto_in_ar_bits_echo_tl_state_source, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@71897.4]
  input         auto_in_r_ready, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@71897.4]
  output        auto_in_r_valid, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@71897.4]
  output [3:0]  auto_in_r_bits_id, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@71897.4]
  output [31:0] auto_in_r_bits_data, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@71897.4]
  output [1:0]  auto_in_r_bits_resp, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@71897.4]
  output [3:0]  auto_in_r_bits_echo_tl_state_size, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@71897.4]
  output [1:0]  auto_in_r_bits_echo_tl_state_source, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@71897.4]
  output        auto_in_r_bits_last, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@71897.4]
  input         auto_out_aw_ready, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@71897.4]
  output        auto_out_aw_valid, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@71897.4]
  output [3:0]  auto_out_aw_bits_id, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@71897.4]
  output [31:0] auto_out_aw_bits_addr, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@71897.4]
  output [7:0]  auto_out_aw_bits_len, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@71897.4]
  output [2:0]  auto_out_aw_bits_size, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@71897.4]
  output [1:0]  auto_out_aw_bits_burst, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@71897.4]
  output        auto_out_aw_bits_lock, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@71897.4]
  output [3:0]  auto_out_aw_bits_cache, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@71897.4]
  output [2:0]  auto_out_aw_bits_prot, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@71897.4]
  output [3:0]  auto_out_aw_bits_qos, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@71897.4]
  input         auto_out_w_ready, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@71897.4]
  output        auto_out_w_valid, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@71897.4]
  output [31:0] auto_out_w_bits_data, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@71897.4]
  output [3:0]  auto_out_w_bits_strb, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@71897.4]
  output        auto_out_w_bits_last, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@71897.4]
  output        auto_out_b_ready, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@71897.4]
  input         auto_out_b_valid, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@71897.4]
  input  [3:0]  auto_out_b_bits_id, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@71897.4]
  input  [1:0]  auto_out_b_bits_resp, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@71897.4]
  input         auto_out_ar_ready, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@71897.4]
  output        auto_out_ar_valid, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@71897.4]
  output [3:0]  auto_out_ar_bits_id, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@71897.4]
  output [31:0] auto_out_ar_bits_addr, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@71897.4]
  output [7:0]  auto_out_ar_bits_len, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@71897.4]
  output [2:0]  auto_out_ar_bits_size, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@71897.4]
  output [1:0]  auto_out_ar_bits_burst, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@71897.4]
  output        auto_out_ar_bits_lock, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@71897.4]
  output [3:0]  auto_out_ar_bits_cache, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@71897.4]
  output [2:0]  auto_out_ar_bits_prot, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@71897.4]
  output [3:0]  auto_out_ar_bits_qos, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@71897.4]
  output        auto_out_r_ready, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@71897.4]
  input         auto_out_r_valid, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@71897.4]
  input  [3:0]  auto_out_r_bits_id, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@71897.4]
  input  [31:0] auto_out_r_bits_data, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@71897.4]
  input  [1:0]  auto_out_r_bits_resp, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@71897.4]
  input         auto_out_r_bits_last // @[:freechips.rocketchip.system.DefaultRV32Config.fir@71897.4]
);
  wire  QueueCompatibility_clock; // @[UserYanker.scala 39:17:freechips.rocketchip.system.DefaultRV32Config.fir@71908.4]
  wire  QueueCompatibility_reset; // @[UserYanker.scala 39:17:freechips.rocketchip.system.DefaultRV32Config.fir@71908.4]
  wire  QueueCompatibility_io_enq_ready; // @[UserYanker.scala 39:17:freechips.rocketchip.system.DefaultRV32Config.fir@71908.4]
  wire  QueueCompatibility_io_enq_valid; // @[UserYanker.scala 39:17:freechips.rocketchip.system.DefaultRV32Config.fir@71908.4]
  wire [3:0] QueueCompatibility_io_enq_bits_tl_state_size; // @[UserYanker.scala 39:17:freechips.rocketchip.system.DefaultRV32Config.fir@71908.4]
  wire [1:0] QueueCompatibility_io_enq_bits_tl_state_source; // @[UserYanker.scala 39:17:freechips.rocketchip.system.DefaultRV32Config.fir@71908.4]
  wire  QueueCompatibility_io_deq_ready; // @[UserYanker.scala 39:17:freechips.rocketchip.system.DefaultRV32Config.fir@71908.4]
  wire  QueueCompatibility_io_deq_valid; // @[UserYanker.scala 39:17:freechips.rocketchip.system.DefaultRV32Config.fir@71908.4]
  wire [3:0] QueueCompatibility_io_deq_bits_tl_state_size; // @[UserYanker.scala 39:17:freechips.rocketchip.system.DefaultRV32Config.fir@71908.4]
  wire [1:0] QueueCompatibility_io_deq_bits_tl_state_source; // @[UserYanker.scala 39:17:freechips.rocketchip.system.DefaultRV32Config.fir@71908.4]
  wire  QueueCompatibility_1_clock; // @[UserYanker.scala 39:17:freechips.rocketchip.system.DefaultRV32Config.fir@71912.4]
  wire  QueueCompatibility_1_reset; // @[UserYanker.scala 39:17:freechips.rocketchip.system.DefaultRV32Config.fir@71912.4]
  wire  QueueCompatibility_1_io_enq_ready; // @[UserYanker.scala 39:17:freechips.rocketchip.system.DefaultRV32Config.fir@71912.4]
  wire  QueueCompatibility_1_io_enq_valid; // @[UserYanker.scala 39:17:freechips.rocketchip.system.DefaultRV32Config.fir@71912.4]
  wire [3:0] QueueCompatibility_1_io_enq_bits_tl_state_size; // @[UserYanker.scala 39:17:freechips.rocketchip.system.DefaultRV32Config.fir@71912.4]
  wire [1:0] QueueCompatibility_1_io_enq_bits_tl_state_source; // @[UserYanker.scala 39:17:freechips.rocketchip.system.DefaultRV32Config.fir@71912.4]
  wire  QueueCompatibility_1_io_deq_ready; // @[UserYanker.scala 39:17:freechips.rocketchip.system.DefaultRV32Config.fir@71912.4]
  wire  QueueCompatibility_1_io_deq_valid; // @[UserYanker.scala 39:17:freechips.rocketchip.system.DefaultRV32Config.fir@71912.4]
  wire [3:0] QueueCompatibility_1_io_deq_bits_tl_state_size; // @[UserYanker.scala 39:17:freechips.rocketchip.system.DefaultRV32Config.fir@71912.4]
  wire [1:0] QueueCompatibility_1_io_deq_bits_tl_state_source; // @[UserYanker.scala 39:17:freechips.rocketchip.system.DefaultRV32Config.fir@71912.4]
  wire  QueueCompatibility_2_clock; // @[UserYanker.scala 39:17:freechips.rocketchip.system.DefaultRV32Config.fir@71916.4]
  wire  QueueCompatibility_2_reset; // @[UserYanker.scala 39:17:freechips.rocketchip.system.DefaultRV32Config.fir@71916.4]
  wire  QueueCompatibility_2_io_enq_ready; // @[UserYanker.scala 39:17:freechips.rocketchip.system.DefaultRV32Config.fir@71916.4]
  wire  QueueCompatibility_2_io_enq_valid; // @[UserYanker.scala 39:17:freechips.rocketchip.system.DefaultRV32Config.fir@71916.4]
  wire [3:0] QueueCompatibility_2_io_enq_bits_tl_state_size; // @[UserYanker.scala 39:17:freechips.rocketchip.system.DefaultRV32Config.fir@71916.4]
  wire [1:0] QueueCompatibility_2_io_enq_bits_tl_state_source; // @[UserYanker.scala 39:17:freechips.rocketchip.system.DefaultRV32Config.fir@71916.4]
  wire  QueueCompatibility_2_io_deq_ready; // @[UserYanker.scala 39:17:freechips.rocketchip.system.DefaultRV32Config.fir@71916.4]
  wire  QueueCompatibility_2_io_deq_valid; // @[UserYanker.scala 39:17:freechips.rocketchip.system.DefaultRV32Config.fir@71916.4]
  wire [3:0] QueueCompatibility_2_io_deq_bits_tl_state_size; // @[UserYanker.scala 39:17:freechips.rocketchip.system.DefaultRV32Config.fir@71916.4]
  wire [1:0] QueueCompatibility_2_io_deq_bits_tl_state_source; // @[UserYanker.scala 39:17:freechips.rocketchip.system.DefaultRV32Config.fir@71916.4]
  wire  QueueCompatibility_3_clock; // @[UserYanker.scala 39:17:freechips.rocketchip.system.DefaultRV32Config.fir@71920.4]
  wire  QueueCompatibility_3_reset; // @[UserYanker.scala 39:17:freechips.rocketchip.system.DefaultRV32Config.fir@71920.4]
  wire  QueueCompatibility_3_io_enq_ready; // @[UserYanker.scala 39:17:freechips.rocketchip.system.DefaultRV32Config.fir@71920.4]
  wire  QueueCompatibility_3_io_enq_valid; // @[UserYanker.scala 39:17:freechips.rocketchip.system.DefaultRV32Config.fir@71920.4]
  wire [3:0] QueueCompatibility_3_io_enq_bits_tl_state_size; // @[UserYanker.scala 39:17:freechips.rocketchip.system.DefaultRV32Config.fir@71920.4]
  wire [1:0] QueueCompatibility_3_io_enq_bits_tl_state_source; // @[UserYanker.scala 39:17:freechips.rocketchip.system.DefaultRV32Config.fir@71920.4]
  wire  QueueCompatibility_3_io_deq_ready; // @[UserYanker.scala 39:17:freechips.rocketchip.system.DefaultRV32Config.fir@71920.4]
  wire  QueueCompatibility_3_io_deq_valid; // @[UserYanker.scala 39:17:freechips.rocketchip.system.DefaultRV32Config.fir@71920.4]
  wire [3:0] QueueCompatibility_3_io_deq_bits_tl_state_size; // @[UserYanker.scala 39:17:freechips.rocketchip.system.DefaultRV32Config.fir@71920.4]
  wire [1:0] QueueCompatibility_3_io_deq_bits_tl_state_source; // @[UserYanker.scala 39:17:freechips.rocketchip.system.DefaultRV32Config.fir@71920.4]
  wire  QueueCompatibility_4_clock; // @[UserYanker.scala 39:17:freechips.rocketchip.system.DefaultRV32Config.fir@71948.4]
  wire  QueueCompatibility_4_reset; // @[UserYanker.scala 39:17:freechips.rocketchip.system.DefaultRV32Config.fir@71948.4]
  wire  QueueCompatibility_4_io_enq_ready; // @[UserYanker.scala 39:17:freechips.rocketchip.system.DefaultRV32Config.fir@71948.4]
  wire  QueueCompatibility_4_io_enq_valid; // @[UserYanker.scala 39:17:freechips.rocketchip.system.DefaultRV32Config.fir@71948.4]
  wire [3:0] QueueCompatibility_4_io_enq_bits_tl_state_size; // @[UserYanker.scala 39:17:freechips.rocketchip.system.DefaultRV32Config.fir@71948.4]
  wire [1:0] QueueCompatibility_4_io_enq_bits_tl_state_source; // @[UserYanker.scala 39:17:freechips.rocketchip.system.DefaultRV32Config.fir@71948.4]
  wire  QueueCompatibility_4_io_deq_ready; // @[UserYanker.scala 39:17:freechips.rocketchip.system.DefaultRV32Config.fir@71948.4]
  wire  QueueCompatibility_4_io_deq_valid; // @[UserYanker.scala 39:17:freechips.rocketchip.system.DefaultRV32Config.fir@71948.4]
  wire [3:0] QueueCompatibility_4_io_deq_bits_tl_state_size; // @[UserYanker.scala 39:17:freechips.rocketchip.system.DefaultRV32Config.fir@71948.4]
  wire [1:0] QueueCompatibility_4_io_deq_bits_tl_state_source; // @[UserYanker.scala 39:17:freechips.rocketchip.system.DefaultRV32Config.fir@71948.4]
  wire  QueueCompatibility_5_clock; // @[UserYanker.scala 39:17:freechips.rocketchip.system.DefaultRV32Config.fir@71952.4]
  wire  QueueCompatibility_5_reset; // @[UserYanker.scala 39:17:freechips.rocketchip.system.DefaultRV32Config.fir@71952.4]
  wire  QueueCompatibility_5_io_enq_ready; // @[UserYanker.scala 39:17:freechips.rocketchip.system.DefaultRV32Config.fir@71952.4]
  wire  QueueCompatibility_5_io_enq_valid; // @[UserYanker.scala 39:17:freechips.rocketchip.system.DefaultRV32Config.fir@71952.4]
  wire [3:0] QueueCompatibility_5_io_enq_bits_tl_state_size; // @[UserYanker.scala 39:17:freechips.rocketchip.system.DefaultRV32Config.fir@71952.4]
  wire [1:0] QueueCompatibility_5_io_enq_bits_tl_state_source; // @[UserYanker.scala 39:17:freechips.rocketchip.system.DefaultRV32Config.fir@71952.4]
  wire  QueueCompatibility_5_io_deq_ready; // @[UserYanker.scala 39:17:freechips.rocketchip.system.DefaultRV32Config.fir@71952.4]
  wire  QueueCompatibility_5_io_deq_valid; // @[UserYanker.scala 39:17:freechips.rocketchip.system.DefaultRV32Config.fir@71952.4]
  wire [3:0] QueueCompatibility_5_io_deq_bits_tl_state_size; // @[UserYanker.scala 39:17:freechips.rocketchip.system.DefaultRV32Config.fir@71952.4]
  wire [1:0] QueueCompatibility_5_io_deq_bits_tl_state_source; // @[UserYanker.scala 39:17:freechips.rocketchip.system.DefaultRV32Config.fir@71952.4]
  wire  QueueCompatibility_6_clock; // @[UserYanker.scala 39:17:freechips.rocketchip.system.DefaultRV32Config.fir@71956.4]
  wire  QueueCompatibility_6_reset; // @[UserYanker.scala 39:17:freechips.rocketchip.system.DefaultRV32Config.fir@71956.4]
  wire  QueueCompatibility_6_io_enq_ready; // @[UserYanker.scala 39:17:freechips.rocketchip.system.DefaultRV32Config.fir@71956.4]
  wire  QueueCompatibility_6_io_enq_valid; // @[UserYanker.scala 39:17:freechips.rocketchip.system.DefaultRV32Config.fir@71956.4]
  wire [3:0] QueueCompatibility_6_io_enq_bits_tl_state_size; // @[UserYanker.scala 39:17:freechips.rocketchip.system.DefaultRV32Config.fir@71956.4]
  wire [1:0] QueueCompatibility_6_io_enq_bits_tl_state_source; // @[UserYanker.scala 39:17:freechips.rocketchip.system.DefaultRV32Config.fir@71956.4]
  wire  QueueCompatibility_6_io_deq_ready; // @[UserYanker.scala 39:17:freechips.rocketchip.system.DefaultRV32Config.fir@71956.4]
  wire  QueueCompatibility_6_io_deq_valid; // @[UserYanker.scala 39:17:freechips.rocketchip.system.DefaultRV32Config.fir@71956.4]
  wire [3:0] QueueCompatibility_6_io_deq_bits_tl_state_size; // @[UserYanker.scala 39:17:freechips.rocketchip.system.DefaultRV32Config.fir@71956.4]
  wire [1:0] QueueCompatibility_6_io_deq_bits_tl_state_source; // @[UserYanker.scala 39:17:freechips.rocketchip.system.DefaultRV32Config.fir@71956.4]
  wire  QueueCompatibility_7_clock; // @[UserYanker.scala 39:17:freechips.rocketchip.system.DefaultRV32Config.fir@71960.4]
  wire  QueueCompatibility_7_reset; // @[UserYanker.scala 39:17:freechips.rocketchip.system.DefaultRV32Config.fir@71960.4]
  wire  QueueCompatibility_7_io_enq_ready; // @[UserYanker.scala 39:17:freechips.rocketchip.system.DefaultRV32Config.fir@71960.4]
  wire  QueueCompatibility_7_io_enq_valid; // @[UserYanker.scala 39:17:freechips.rocketchip.system.DefaultRV32Config.fir@71960.4]
  wire [3:0] QueueCompatibility_7_io_enq_bits_tl_state_size; // @[UserYanker.scala 39:17:freechips.rocketchip.system.DefaultRV32Config.fir@71960.4]
  wire [1:0] QueueCompatibility_7_io_enq_bits_tl_state_source; // @[UserYanker.scala 39:17:freechips.rocketchip.system.DefaultRV32Config.fir@71960.4]
  wire  QueueCompatibility_7_io_deq_ready; // @[UserYanker.scala 39:17:freechips.rocketchip.system.DefaultRV32Config.fir@71960.4]
  wire  QueueCompatibility_7_io_deq_valid; // @[UserYanker.scala 39:17:freechips.rocketchip.system.DefaultRV32Config.fir@71960.4]
  wire [3:0] QueueCompatibility_7_io_deq_bits_tl_state_size; // @[UserYanker.scala 39:17:freechips.rocketchip.system.DefaultRV32Config.fir@71960.4]
  wire [1:0] QueueCompatibility_7_io_deq_bits_tl_state_source; // @[UserYanker.scala 39:17:freechips.rocketchip.system.DefaultRV32Config.fir@71960.4]
  wire  _T_26_0; // @[UserYanker.scala 47:25:freechips.rocketchip.system.DefaultRV32Config.fir@71988.4 UserYanker.scala 47:25:freechips.rocketchip.system.DefaultRV32Config.fir@71990.4]
  wire  _T_26_1; // @[UserYanker.scala 47:25:freechips.rocketchip.system.DefaultRV32Config.fir@71988.4 UserYanker.scala 47:25:freechips.rocketchip.system.DefaultRV32Config.fir@71991.4]
  wire  _GEN_1; // @[UserYanker.scala 48:36:freechips.rocketchip.system.DefaultRV32Config.fir@72006.4]
  wire  _T_26_2; // @[UserYanker.scala 47:25:freechips.rocketchip.system.DefaultRV32Config.fir@71988.4 UserYanker.scala 47:25:freechips.rocketchip.system.DefaultRV32Config.fir@71992.4]
  wire  _GEN_2; // @[UserYanker.scala 48:36:freechips.rocketchip.system.DefaultRV32Config.fir@72006.4]
  wire  _T_26_3; // @[UserYanker.scala 47:25:freechips.rocketchip.system.DefaultRV32Config.fir@71988.4 UserYanker.scala 47:25:freechips.rocketchip.system.DefaultRV32Config.fir@71993.4]
  wire  _GEN_3; // @[UserYanker.scala 48:36:freechips.rocketchip.system.DefaultRV32Config.fir@72006.4]
  wire  _GEN_4; // @[UserYanker.scala 48:36:freechips.rocketchip.system.DefaultRV32Config.fir@72006.4]
  wire  _GEN_5; // @[UserYanker.scala 48:36:freechips.rocketchip.system.DefaultRV32Config.fir@72006.4]
  wire  _GEN_6; // @[UserYanker.scala 48:36:freechips.rocketchip.system.DefaultRV32Config.fir@72006.4]
  wire  _GEN_7; // @[UserYanker.scala 48:36:freechips.rocketchip.system.DefaultRV32Config.fir@72006.4]
  wire  _GEN_8; // @[UserYanker.scala 48:36:freechips.rocketchip.system.DefaultRV32Config.fir@72006.4]
  wire  _GEN_9; // @[UserYanker.scala 48:36:freechips.rocketchip.system.DefaultRV32Config.fir@72006.4]
  wire  _GEN_10; // @[UserYanker.scala 48:36:freechips.rocketchip.system.DefaultRV32Config.fir@72006.4]
  wire  _GEN_11; // @[UserYanker.scala 48:36:freechips.rocketchip.system.DefaultRV32Config.fir@72006.4]
  wire  _GEN_12; // @[UserYanker.scala 48:36:freechips.rocketchip.system.DefaultRV32Config.fir@72006.4]
  wire  _GEN_13; // @[UserYanker.scala 48:36:freechips.rocketchip.system.DefaultRV32Config.fir@72006.4]
  wire  _GEN_14; // @[UserYanker.scala 48:36:freechips.rocketchip.system.DefaultRV32Config.fir@72006.4]
  wire  _GEN_15; // @[UserYanker.scala 48:36:freechips.rocketchip.system.DefaultRV32Config.fir@72006.4]
  wire  _T_31; // @[UserYanker.scala 55:15:freechips.rocketchip.system.DefaultRV32Config.fir@72055.4]
  wire  _T_29_0; // @[UserYanker.scala 53:24:freechips.rocketchip.system.DefaultRV32Config.fir@72019.4 UserYanker.scala 53:24:freechips.rocketchip.system.DefaultRV32Config.fir@72021.4]
  wire  _T_29_1; // @[UserYanker.scala 53:24:freechips.rocketchip.system.DefaultRV32Config.fir@72019.4 UserYanker.scala 53:24:freechips.rocketchip.system.DefaultRV32Config.fir@72022.4]
  wire  _GEN_17; // @[UserYanker.scala 55:28:freechips.rocketchip.system.DefaultRV32Config.fir@72056.4]
  wire  _T_29_2; // @[UserYanker.scala 53:24:freechips.rocketchip.system.DefaultRV32Config.fir@72019.4 UserYanker.scala 53:24:freechips.rocketchip.system.DefaultRV32Config.fir@72023.4]
  wire  _GEN_18; // @[UserYanker.scala 55:28:freechips.rocketchip.system.DefaultRV32Config.fir@72056.4]
  wire  _T_29_3; // @[UserYanker.scala 53:24:freechips.rocketchip.system.DefaultRV32Config.fir@72019.4 UserYanker.scala 53:24:freechips.rocketchip.system.DefaultRV32Config.fir@72024.4]
  wire  _GEN_19; // @[UserYanker.scala 55:28:freechips.rocketchip.system.DefaultRV32Config.fir@72056.4]
  wire  _GEN_20; // @[UserYanker.scala 55:28:freechips.rocketchip.system.DefaultRV32Config.fir@72056.4]
  wire  _GEN_21; // @[UserYanker.scala 55:28:freechips.rocketchip.system.DefaultRV32Config.fir@72056.4]
  wire  _GEN_22; // @[UserYanker.scala 55:28:freechips.rocketchip.system.DefaultRV32Config.fir@72056.4]
  wire  _GEN_23; // @[UserYanker.scala 55:28:freechips.rocketchip.system.DefaultRV32Config.fir@72056.4]
  wire  _GEN_24; // @[UserYanker.scala 55:28:freechips.rocketchip.system.DefaultRV32Config.fir@72056.4]
  wire  _GEN_25; // @[UserYanker.scala 55:28:freechips.rocketchip.system.DefaultRV32Config.fir@72056.4]
  wire  _GEN_26; // @[UserYanker.scala 55:28:freechips.rocketchip.system.DefaultRV32Config.fir@72056.4]
  wire  _GEN_27; // @[UserYanker.scala 55:28:freechips.rocketchip.system.DefaultRV32Config.fir@72056.4]
  wire  _GEN_28; // @[UserYanker.scala 55:28:freechips.rocketchip.system.DefaultRV32Config.fir@72056.4]
  wire  _GEN_29; // @[UserYanker.scala 55:28:freechips.rocketchip.system.DefaultRV32Config.fir@72056.4]
  wire  _GEN_30; // @[UserYanker.scala 55:28:freechips.rocketchip.system.DefaultRV32Config.fir@72056.4]
  wire  _GEN_31; // @[UserYanker.scala 55:28:freechips.rocketchip.system.DefaultRV32Config.fir@72056.4]
  wire  _T_32; // @[UserYanker.scala 55:28:freechips.rocketchip.system.DefaultRV32Config.fir@72056.4]
  wire  _T_34; // @[UserYanker.scala 55:14:freechips.rocketchip.system.DefaultRV32Config.fir@72058.4]
  wire  _T_35; // @[UserYanker.scala 55:14:freechips.rocketchip.system.DefaultRV32Config.fir@72059.4]
  wire [3:0] _T_30_0_tl_state_size; // @[UserYanker.scala 54:23:freechips.rocketchip.system.DefaultRV32Config.fir@72037.4 UserYanker.scala 54:23:freechips.rocketchip.system.DefaultRV32Config.fir@72039.4]
  wire [1:0] _T_30_0_tl_state_source; // @[UserYanker.scala 54:23:freechips.rocketchip.system.DefaultRV32Config.fir@72037.4 UserYanker.scala 54:23:freechips.rocketchip.system.DefaultRV32Config.fir@72039.4]
  wire [3:0] _T_30_1_tl_state_size; // @[UserYanker.scala 54:23:freechips.rocketchip.system.DefaultRV32Config.fir@72037.4 UserYanker.scala 54:23:freechips.rocketchip.system.DefaultRV32Config.fir@72040.4]
  wire [3:0] _GEN_34; // @[BundleMap.scala 248:19:freechips.rocketchip.system.DefaultRV32Config.fir@72072.4]
  wire [1:0] _T_30_1_tl_state_source; // @[UserYanker.scala 54:23:freechips.rocketchip.system.DefaultRV32Config.fir@72037.4 UserYanker.scala 54:23:freechips.rocketchip.system.DefaultRV32Config.fir@72040.4]
  wire [1:0] _GEN_35; // @[BundleMap.scala 248:19:freechips.rocketchip.system.DefaultRV32Config.fir@72072.4]
  wire [3:0] _T_30_2_tl_state_size; // @[UserYanker.scala 54:23:freechips.rocketchip.system.DefaultRV32Config.fir@72037.4 UserYanker.scala 54:23:freechips.rocketchip.system.DefaultRV32Config.fir@72041.4]
  wire [3:0] _GEN_36; // @[BundleMap.scala 248:19:freechips.rocketchip.system.DefaultRV32Config.fir@72072.4]
  wire [1:0] _T_30_2_tl_state_source; // @[UserYanker.scala 54:23:freechips.rocketchip.system.DefaultRV32Config.fir@72037.4 UserYanker.scala 54:23:freechips.rocketchip.system.DefaultRV32Config.fir@72041.4]
  wire [1:0] _GEN_37; // @[BundleMap.scala 248:19:freechips.rocketchip.system.DefaultRV32Config.fir@72072.4]
  wire [3:0] _T_30_3_tl_state_size; // @[UserYanker.scala 54:23:freechips.rocketchip.system.DefaultRV32Config.fir@72037.4 UserYanker.scala 54:23:freechips.rocketchip.system.DefaultRV32Config.fir@72042.4]
  wire [3:0] _GEN_38; // @[BundleMap.scala 248:19:freechips.rocketchip.system.DefaultRV32Config.fir@72072.4]
  wire [1:0] _T_30_3_tl_state_source; // @[UserYanker.scala 54:23:freechips.rocketchip.system.DefaultRV32Config.fir@72037.4 UserYanker.scala 54:23:freechips.rocketchip.system.DefaultRV32Config.fir@72042.4]
  wire [1:0] _GEN_39; // @[BundleMap.scala 248:19:freechips.rocketchip.system.DefaultRV32Config.fir@72072.4]
  wire [3:0] _GEN_40; // @[BundleMap.scala 248:19:freechips.rocketchip.system.DefaultRV32Config.fir@72072.4]
  wire [1:0] _GEN_41; // @[BundleMap.scala 248:19:freechips.rocketchip.system.DefaultRV32Config.fir@72072.4]
  wire [3:0] _GEN_42; // @[BundleMap.scala 248:19:freechips.rocketchip.system.DefaultRV32Config.fir@72072.4]
  wire [1:0] _GEN_43; // @[BundleMap.scala 248:19:freechips.rocketchip.system.DefaultRV32Config.fir@72072.4]
  wire [3:0] _GEN_44; // @[BundleMap.scala 248:19:freechips.rocketchip.system.DefaultRV32Config.fir@72072.4]
  wire [1:0] _GEN_45; // @[BundleMap.scala 248:19:freechips.rocketchip.system.DefaultRV32Config.fir@72072.4]
  wire [3:0] _GEN_46; // @[BundleMap.scala 248:19:freechips.rocketchip.system.DefaultRV32Config.fir@72072.4]
  wire [1:0] _GEN_47; // @[BundleMap.scala 248:19:freechips.rocketchip.system.DefaultRV32Config.fir@72072.4]
  wire [3:0] _GEN_48; // @[BundleMap.scala 248:19:freechips.rocketchip.system.DefaultRV32Config.fir@72072.4]
  wire [1:0] _GEN_49; // @[BundleMap.scala 248:19:freechips.rocketchip.system.DefaultRV32Config.fir@72072.4]
  wire [3:0] _GEN_50; // @[BundleMap.scala 248:19:freechips.rocketchip.system.DefaultRV32Config.fir@72072.4]
  wire [1:0] _GEN_51; // @[BundleMap.scala 248:19:freechips.rocketchip.system.DefaultRV32Config.fir@72072.4]
  wire [3:0] _GEN_52; // @[BundleMap.scala 248:19:freechips.rocketchip.system.DefaultRV32Config.fir@72072.4]
  wire [1:0] _GEN_53; // @[BundleMap.scala 248:19:freechips.rocketchip.system.DefaultRV32Config.fir@72072.4]
  wire [3:0] _GEN_54; // @[BundleMap.scala 248:19:freechips.rocketchip.system.DefaultRV32Config.fir@72072.4]
  wire [1:0] _GEN_55; // @[BundleMap.scala 248:19:freechips.rocketchip.system.DefaultRV32Config.fir@72072.4]
  wire [3:0] _GEN_56; // @[BundleMap.scala 248:19:freechips.rocketchip.system.DefaultRV32Config.fir@72072.4]
  wire [1:0] _GEN_57; // @[BundleMap.scala 248:19:freechips.rocketchip.system.DefaultRV32Config.fir@72072.4]
  wire [3:0] _GEN_58; // @[BundleMap.scala 248:19:freechips.rocketchip.system.DefaultRV32Config.fir@72072.4]
  wire [1:0] _GEN_59; // @[BundleMap.scala 248:19:freechips.rocketchip.system.DefaultRV32Config.fir@72072.4]
  wire [3:0] _GEN_60; // @[BundleMap.scala 248:19:freechips.rocketchip.system.DefaultRV32Config.fir@72072.4]
  wire [1:0] _GEN_61; // @[BundleMap.scala 248:19:freechips.rocketchip.system.DefaultRV32Config.fir@72072.4]
  wire [15:0] _T_37; // @[OneHot.scala 65:12:freechips.rocketchip.system.DefaultRV32Config.fir@72075.4]
  wire [15:0] _T_56; // @[OneHot.scala 65:12:freechips.rocketchip.system.DefaultRV32Config.fir@72094.4]
  wire  _T_74; // @[UserYanker.scala 62:37:freechips.rocketchip.system.DefaultRV32Config.fir@72112.4]
  wire  _T_75; // @[UserYanker.scala 62:53:freechips.rocketchip.system.DefaultRV32Config.fir@72113.4]
  wire  _T_77; // @[UserYanker.scala 63:37:freechips.rocketchip.system.DefaultRV32Config.fir@72116.4]
  wire  _T_80; // @[UserYanker.scala 62:53:freechips.rocketchip.system.DefaultRV32Config.fir@72122.4]
  wire  _T_85; // @[UserYanker.scala 62:53:freechips.rocketchip.system.DefaultRV32Config.fir@72131.4]
  wire  _T_90; // @[UserYanker.scala 62:53:freechips.rocketchip.system.DefaultRV32Config.fir@72140.4]
  wire  _T_154_0; // @[UserYanker.scala 68:25:freechips.rocketchip.system.DefaultRV32Config.fir@72256.4 UserYanker.scala 68:25:freechips.rocketchip.system.DefaultRV32Config.fir@72258.4]
  wire  _T_154_1; // @[UserYanker.scala 68:25:freechips.rocketchip.system.DefaultRV32Config.fir@72256.4 UserYanker.scala 68:25:freechips.rocketchip.system.DefaultRV32Config.fir@72259.4]
  wire  _GEN_65; // @[UserYanker.scala 69:36:freechips.rocketchip.system.DefaultRV32Config.fir@72274.4]
  wire  _T_154_2; // @[UserYanker.scala 68:25:freechips.rocketchip.system.DefaultRV32Config.fir@72256.4 UserYanker.scala 68:25:freechips.rocketchip.system.DefaultRV32Config.fir@72260.4]
  wire  _GEN_66; // @[UserYanker.scala 69:36:freechips.rocketchip.system.DefaultRV32Config.fir@72274.4]
  wire  _T_154_3; // @[UserYanker.scala 68:25:freechips.rocketchip.system.DefaultRV32Config.fir@72256.4 UserYanker.scala 68:25:freechips.rocketchip.system.DefaultRV32Config.fir@72261.4]
  wire  _GEN_67; // @[UserYanker.scala 69:36:freechips.rocketchip.system.DefaultRV32Config.fir@72274.4]
  wire  _GEN_68; // @[UserYanker.scala 69:36:freechips.rocketchip.system.DefaultRV32Config.fir@72274.4]
  wire  _GEN_69; // @[UserYanker.scala 69:36:freechips.rocketchip.system.DefaultRV32Config.fir@72274.4]
  wire  _GEN_70; // @[UserYanker.scala 69:36:freechips.rocketchip.system.DefaultRV32Config.fir@72274.4]
  wire  _GEN_71; // @[UserYanker.scala 69:36:freechips.rocketchip.system.DefaultRV32Config.fir@72274.4]
  wire  _GEN_72; // @[UserYanker.scala 69:36:freechips.rocketchip.system.DefaultRV32Config.fir@72274.4]
  wire  _GEN_73; // @[UserYanker.scala 69:36:freechips.rocketchip.system.DefaultRV32Config.fir@72274.4]
  wire  _GEN_74; // @[UserYanker.scala 69:36:freechips.rocketchip.system.DefaultRV32Config.fir@72274.4]
  wire  _GEN_75; // @[UserYanker.scala 69:36:freechips.rocketchip.system.DefaultRV32Config.fir@72274.4]
  wire  _GEN_76; // @[UserYanker.scala 69:36:freechips.rocketchip.system.DefaultRV32Config.fir@72274.4]
  wire  _GEN_77; // @[UserYanker.scala 69:36:freechips.rocketchip.system.DefaultRV32Config.fir@72274.4]
  wire  _GEN_78; // @[UserYanker.scala 69:36:freechips.rocketchip.system.DefaultRV32Config.fir@72274.4]
  wire  _GEN_79; // @[UserYanker.scala 69:36:freechips.rocketchip.system.DefaultRV32Config.fir@72274.4]
  wire  _T_159; // @[UserYanker.scala 76:15:freechips.rocketchip.system.DefaultRV32Config.fir@72323.4]
  wire  _T_157_0; // @[UserYanker.scala 74:24:freechips.rocketchip.system.DefaultRV32Config.fir@72287.4 UserYanker.scala 74:24:freechips.rocketchip.system.DefaultRV32Config.fir@72289.4]
  wire  _T_157_1; // @[UserYanker.scala 74:24:freechips.rocketchip.system.DefaultRV32Config.fir@72287.4 UserYanker.scala 74:24:freechips.rocketchip.system.DefaultRV32Config.fir@72290.4]
  wire  _GEN_81; // @[UserYanker.scala 76:28:freechips.rocketchip.system.DefaultRV32Config.fir@72324.4]
  wire  _T_157_2; // @[UserYanker.scala 74:24:freechips.rocketchip.system.DefaultRV32Config.fir@72287.4 UserYanker.scala 74:24:freechips.rocketchip.system.DefaultRV32Config.fir@72291.4]
  wire  _GEN_82; // @[UserYanker.scala 76:28:freechips.rocketchip.system.DefaultRV32Config.fir@72324.4]
  wire  _T_157_3; // @[UserYanker.scala 74:24:freechips.rocketchip.system.DefaultRV32Config.fir@72287.4 UserYanker.scala 74:24:freechips.rocketchip.system.DefaultRV32Config.fir@72292.4]
  wire  _GEN_83; // @[UserYanker.scala 76:28:freechips.rocketchip.system.DefaultRV32Config.fir@72324.4]
  wire  _GEN_84; // @[UserYanker.scala 76:28:freechips.rocketchip.system.DefaultRV32Config.fir@72324.4]
  wire  _GEN_85; // @[UserYanker.scala 76:28:freechips.rocketchip.system.DefaultRV32Config.fir@72324.4]
  wire  _GEN_86; // @[UserYanker.scala 76:28:freechips.rocketchip.system.DefaultRV32Config.fir@72324.4]
  wire  _GEN_87; // @[UserYanker.scala 76:28:freechips.rocketchip.system.DefaultRV32Config.fir@72324.4]
  wire  _GEN_88; // @[UserYanker.scala 76:28:freechips.rocketchip.system.DefaultRV32Config.fir@72324.4]
  wire  _GEN_89; // @[UserYanker.scala 76:28:freechips.rocketchip.system.DefaultRV32Config.fir@72324.4]
  wire  _GEN_90; // @[UserYanker.scala 76:28:freechips.rocketchip.system.DefaultRV32Config.fir@72324.4]
  wire  _GEN_91; // @[UserYanker.scala 76:28:freechips.rocketchip.system.DefaultRV32Config.fir@72324.4]
  wire  _GEN_92; // @[UserYanker.scala 76:28:freechips.rocketchip.system.DefaultRV32Config.fir@72324.4]
  wire  _GEN_93; // @[UserYanker.scala 76:28:freechips.rocketchip.system.DefaultRV32Config.fir@72324.4]
  wire  _GEN_94; // @[UserYanker.scala 76:28:freechips.rocketchip.system.DefaultRV32Config.fir@72324.4]
  wire  _GEN_95; // @[UserYanker.scala 76:28:freechips.rocketchip.system.DefaultRV32Config.fir@72324.4]
  wire  _T_160; // @[UserYanker.scala 76:28:freechips.rocketchip.system.DefaultRV32Config.fir@72324.4]
  wire  _T_162; // @[UserYanker.scala 76:14:freechips.rocketchip.system.DefaultRV32Config.fir@72326.4]
  wire  _T_163; // @[UserYanker.scala 76:14:freechips.rocketchip.system.DefaultRV32Config.fir@72327.4]
  wire [3:0] _T_158_0_tl_state_size; // @[UserYanker.scala 75:23:freechips.rocketchip.system.DefaultRV32Config.fir@72305.4 UserYanker.scala 75:23:freechips.rocketchip.system.DefaultRV32Config.fir@72307.4]
  wire [1:0] _T_158_0_tl_state_source; // @[UserYanker.scala 75:23:freechips.rocketchip.system.DefaultRV32Config.fir@72305.4 UserYanker.scala 75:23:freechips.rocketchip.system.DefaultRV32Config.fir@72307.4]
  wire [3:0] _T_158_1_tl_state_size; // @[UserYanker.scala 75:23:freechips.rocketchip.system.DefaultRV32Config.fir@72305.4 UserYanker.scala 75:23:freechips.rocketchip.system.DefaultRV32Config.fir@72308.4]
  wire [3:0] _GEN_98; // @[BundleMap.scala 248:19:freechips.rocketchip.system.DefaultRV32Config.fir@72338.4]
  wire [1:0] _T_158_1_tl_state_source; // @[UserYanker.scala 75:23:freechips.rocketchip.system.DefaultRV32Config.fir@72305.4 UserYanker.scala 75:23:freechips.rocketchip.system.DefaultRV32Config.fir@72308.4]
  wire [1:0] _GEN_99; // @[BundleMap.scala 248:19:freechips.rocketchip.system.DefaultRV32Config.fir@72338.4]
  wire [3:0] _T_158_2_tl_state_size; // @[UserYanker.scala 75:23:freechips.rocketchip.system.DefaultRV32Config.fir@72305.4 UserYanker.scala 75:23:freechips.rocketchip.system.DefaultRV32Config.fir@72309.4]
  wire [3:0] _GEN_100; // @[BundleMap.scala 248:19:freechips.rocketchip.system.DefaultRV32Config.fir@72338.4]
  wire [1:0] _T_158_2_tl_state_source; // @[UserYanker.scala 75:23:freechips.rocketchip.system.DefaultRV32Config.fir@72305.4 UserYanker.scala 75:23:freechips.rocketchip.system.DefaultRV32Config.fir@72309.4]
  wire [1:0] _GEN_101; // @[BundleMap.scala 248:19:freechips.rocketchip.system.DefaultRV32Config.fir@72338.4]
  wire [3:0] _T_158_3_tl_state_size; // @[UserYanker.scala 75:23:freechips.rocketchip.system.DefaultRV32Config.fir@72305.4 UserYanker.scala 75:23:freechips.rocketchip.system.DefaultRV32Config.fir@72310.4]
  wire [3:0] _GEN_102; // @[BundleMap.scala 248:19:freechips.rocketchip.system.DefaultRV32Config.fir@72338.4]
  wire [1:0] _T_158_3_tl_state_source; // @[UserYanker.scala 75:23:freechips.rocketchip.system.DefaultRV32Config.fir@72305.4 UserYanker.scala 75:23:freechips.rocketchip.system.DefaultRV32Config.fir@72310.4]
  wire [1:0] _GEN_103; // @[BundleMap.scala 248:19:freechips.rocketchip.system.DefaultRV32Config.fir@72338.4]
  wire [3:0] _GEN_104; // @[BundleMap.scala 248:19:freechips.rocketchip.system.DefaultRV32Config.fir@72338.4]
  wire [1:0] _GEN_105; // @[BundleMap.scala 248:19:freechips.rocketchip.system.DefaultRV32Config.fir@72338.4]
  wire [3:0] _GEN_106; // @[BundleMap.scala 248:19:freechips.rocketchip.system.DefaultRV32Config.fir@72338.4]
  wire [1:0] _GEN_107; // @[BundleMap.scala 248:19:freechips.rocketchip.system.DefaultRV32Config.fir@72338.4]
  wire [3:0] _GEN_108; // @[BundleMap.scala 248:19:freechips.rocketchip.system.DefaultRV32Config.fir@72338.4]
  wire [1:0] _GEN_109; // @[BundleMap.scala 248:19:freechips.rocketchip.system.DefaultRV32Config.fir@72338.4]
  wire [3:0] _GEN_110; // @[BundleMap.scala 248:19:freechips.rocketchip.system.DefaultRV32Config.fir@72338.4]
  wire [1:0] _GEN_111; // @[BundleMap.scala 248:19:freechips.rocketchip.system.DefaultRV32Config.fir@72338.4]
  wire [3:0] _GEN_112; // @[BundleMap.scala 248:19:freechips.rocketchip.system.DefaultRV32Config.fir@72338.4]
  wire [1:0] _GEN_113; // @[BundleMap.scala 248:19:freechips.rocketchip.system.DefaultRV32Config.fir@72338.4]
  wire [3:0] _GEN_114; // @[BundleMap.scala 248:19:freechips.rocketchip.system.DefaultRV32Config.fir@72338.4]
  wire [1:0] _GEN_115; // @[BundleMap.scala 248:19:freechips.rocketchip.system.DefaultRV32Config.fir@72338.4]
  wire [3:0] _GEN_116; // @[BundleMap.scala 248:19:freechips.rocketchip.system.DefaultRV32Config.fir@72338.4]
  wire [1:0] _GEN_117; // @[BundleMap.scala 248:19:freechips.rocketchip.system.DefaultRV32Config.fir@72338.4]
  wire [3:0] _GEN_118; // @[BundleMap.scala 248:19:freechips.rocketchip.system.DefaultRV32Config.fir@72338.4]
  wire [1:0] _GEN_119; // @[BundleMap.scala 248:19:freechips.rocketchip.system.DefaultRV32Config.fir@72338.4]
  wire [3:0] _GEN_120; // @[BundleMap.scala 248:19:freechips.rocketchip.system.DefaultRV32Config.fir@72338.4]
  wire [1:0] _GEN_121; // @[BundleMap.scala 248:19:freechips.rocketchip.system.DefaultRV32Config.fir@72338.4]
  wire [3:0] _GEN_122; // @[BundleMap.scala 248:19:freechips.rocketchip.system.DefaultRV32Config.fir@72338.4]
  wire [1:0] _GEN_123; // @[BundleMap.scala 248:19:freechips.rocketchip.system.DefaultRV32Config.fir@72338.4]
  wire [3:0] _GEN_124; // @[BundleMap.scala 248:19:freechips.rocketchip.system.DefaultRV32Config.fir@72338.4]
  wire [1:0] _GEN_125; // @[BundleMap.scala 248:19:freechips.rocketchip.system.DefaultRV32Config.fir@72338.4]
  wire [15:0] _T_165; // @[OneHot.scala 65:12:freechips.rocketchip.system.DefaultRV32Config.fir@72341.4]
  wire [15:0] _T_184; // @[OneHot.scala 65:12:freechips.rocketchip.system.DefaultRV32Config.fir@72360.4]
  wire  _T_202; // @[UserYanker.scala 83:37:freechips.rocketchip.system.DefaultRV32Config.fir@72378.4]
  wire  _T_204; // @[UserYanker.scala 84:37:freechips.rocketchip.system.DefaultRV32Config.fir@72381.4]
  QueueCompatibility_14 QueueCompatibility ( // @[UserYanker.scala 39:17:freechips.rocketchip.system.DefaultRV32Config.fir@71908.4]
    .clock(QueueCompatibility_clock),
    .reset(QueueCompatibility_reset),
    .io_enq_ready(QueueCompatibility_io_enq_ready),
    .io_enq_valid(QueueCompatibility_io_enq_valid),
    .io_enq_bits_tl_state_size(QueueCompatibility_io_enq_bits_tl_state_size),
    .io_enq_bits_tl_state_source(QueueCompatibility_io_enq_bits_tl_state_source),
    .io_deq_ready(QueueCompatibility_io_deq_ready),
    .io_deq_valid(QueueCompatibility_io_deq_valid),
    .io_deq_bits_tl_state_size(QueueCompatibility_io_deq_bits_tl_state_size),
    .io_deq_bits_tl_state_source(QueueCompatibility_io_deq_bits_tl_state_source)
  );
  QueueCompatibility_14 QueueCompatibility_1 ( // @[UserYanker.scala 39:17:freechips.rocketchip.system.DefaultRV32Config.fir@71912.4]
    .clock(QueueCompatibility_1_clock),
    .reset(QueueCompatibility_1_reset),
    .io_enq_ready(QueueCompatibility_1_io_enq_ready),
    .io_enq_valid(QueueCompatibility_1_io_enq_valid),
    .io_enq_bits_tl_state_size(QueueCompatibility_1_io_enq_bits_tl_state_size),
    .io_enq_bits_tl_state_source(QueueCompatibility_1_io_enq_bits_tl_state_source),
    .io_deq_ready(QueueCompatibility_1_io_deq_ready),
    .io_deq_valid(QueueCompatibility_1_io_deq_valid),
    .io_deq_bits_tl_state_size(QueueCompatibility_1_io_deq_bits_tl_state_size),
    .io_deq_bits_tl_state_source(QueueCompatibility_1_io_deq_bits_tl_state_source)
  );
  QueueCompatibility_14 QueueCompatibility_2 ( // @[UserYanker.scala 39:17:freechips.rocketchip.system.DefaultRV32Config.fir@71916.4]
    .clock(QueueCompatibility_2_clock),
    .reset(QueueCompatibility_2_reset),
    .io_enq_ready(QueueCompatibility_2_io_enq_ready),
    .io_enq_valid(QueueCompatibility_2_io_enq_valid),
    .io_enq_bits_tl_state_size(QueueCompatibility_2_io_enq_bits_tl_state_size),
    .io_enq_bits_tl_state_source(QueueCompatibility_2_io_enq_bits_tl_state_source),
    .io_deq_ready(QueueCompatibility_2_io_deq_ready),
    .io_deq_valid(QueueCompatibility_2_io_deq_valid),
    .io_deq_bits_tl_state_size(QueueCompatibility_2_io_deq_bits_tl_state_size),
    .io_deq_bits_tl_state_source(QueueCompatibility_2_io_deq_bits_tl_state_source)
  );
  QueueCompatibility_14 QueueCompatibility_3 ( // @[UserYanker.scala 39:17:freechips.rocketchip.system.DefaultRV32Config.fir@71920.4]
    .clock(QueueCompatibility_3_clock),
    .reset(QueueCompatibility_3_reset),
    .io_enq_ready(QueueCompatibility_3_io_enq_ready),
    .io_enq_valid(QueueCompatibility_3_io_enq_valid),
    .io_enq_bits_tl_state_size(QueueCompatibility_3_io_enq_bits_tl_state_size),
    .io_enq_bits_tl_state_source(QueueCompatibility_3_io_enq_bits_tl_state_source),
    .io_deq_ready(QueueCompatibility_3_io_deq_ready),
    .io_deq_valid(QueueCompatibility_3_io_deq_valid),
    .io_deq_bits_tl_state_size(QueueCompatibility_3_io_deq_bits_tl_state_size),
    .io_deq_bits_tl_state_source(QueueCompatibility_3_io_deq_bits_tl_state_source)
  );
  QueueCompatibility_14 QueueCompatibility_4 ( // @[UserYanker.scala 39:17:freechips.rocketchip.system.DefaultRV32Config.fir@71948.4]
    .clock(QueueCompatibility_4_clock),
    .reset(QueueCompatibility_4_reset),
    .io_enq_ready(QueueCompatibility_4_io_enq_ready),
    .io_enq_valid(QueueCompatibility_4_io_enq_valid),
    .io_enq_bits_tl_state_size(QueueCompatibility_4_io_enq_bits_tl_state_size),
    .io_enq_bits_tl_state_source(QueueCompatibility_4_io_enq_bits_tl_state_source),
    .io_deq_ready(QueueCompatibility_4_io_deq_ready),
    .io_deq_valid(QueueCompatibility_4_io_deq_valid),
    .io_deq_bits_tl_state_size(QueueCompatibility_4_io_deq_bits_tl_state_size),
    .io_deq_bits_tl_state_source(QueueCompatibility_4_io_deq_bits_tl_state_source)
  );
  QueueCompatibility_14 QueueCompatibility_5 ( // @[UserYanker.scala 39:17:freechips.rocketchip.system.DefaultRV32Config.fir@71952.4]
    .clock(QueueCompatibility_5_clock),
    .reset(QueueCompatibility_5_reset),
    .io_enq_ready(QueueCompatibility_5_io_enq_ready),
    .io_enq_valid(QueueCompatibility_5_io_enq_valid),
    .io_enq_bits_tl_state_size(QueueCompatibility_5_io_enq_bits_tl_state_size),
    .io_enq_bits_tl_state_source(QueueCompatibility_5_io_enq_bits_tl_state_source),
    .io_deq_ready(QueueCompatibility_5_io_deq_ready),
    .io_deq_valid(QueueCompatibility_5_io_deq_valid),
    .io_deq_bits_tl_state_size(QueueCompatibility_5_io_deq_bits_tl_state_size),
    .io_deq_bits_tl_state_source(QueueCompatibility_5_io_deq_bits_tl_state_source)
  );
  QueueCompatibility_14 QueueCompatibility_6 ( // @[UserYanker.scala 39:17:freechips.rocketchip.system.DefaultRV32Config.fir@71956.4]
    .clock(QueueCompatibility_6_clock),
    .reset(QueueCompatibility_6_reset),
    .io_enq_ready(QueueCompatibility_6_io_enq_ready),
    .io_enq_valid(QueueCompatibility_6_io_enq_valid),
    .io_enq_bits_tl_state_size(QueueCompatibility_6_io_enq_bits_tl_state_size),
    .io_enq_bits_tl_state_source(QueueCompatibility_6_io_enq_bits_tl_state_source),
    .io_deq_ready(QueueCompatibility_6_io_deq_ready),
    .io_deq_valid(QueueCompatibility_6_io_deq_valid),
    .io_deq_bits_tl_state_size(QueueCompatibility_6_io_deq_bits_tl_state_size),
    .io_deq_bits_tl_state_source(QueueCompatibility_6_io_deq_bits_tl_state_source)
  );
  QueueCompatibility_14 QueueCompatibility_7 ( // @[UserYanker.scala 39:17:freechips.rocketchip.system.DefaultRV32Config.fir@71960.4]
    .clock(QueueCompatibility_7_clock),
    .reset(QueueCompatibility_7_reset),
    .io_enq_ready(QueueCompatibility_7_io_enq_ready),
    .io_enq_valid(QueueCompatibility_7_io_enq_valid),
    .io_enq_bits_tl_state_size(QueueCompatibility_7_io_enq_bits_tl_state_size),
    .io_enq_bits_tl_state_source(QueueCompatibility_7_io_enq_bits_tl_state_source),
    .io_deq_ready(QueueCompatibility_7_io_deq_ready),
    .io_deq_valid(QueueCompatibility_7_io_deq_valid),
    .io_deq_bits_tl_state_size(QueueCompatibility_7_io_deq_bits_tl_state_size),
    .io_deq_bits_tl_state_source(QueueCompatibility_7_io_deq_bits_tl_state_source)
  );
  assign _T_26_0 = QueueCompatibility_io_enq_ready; // @[UserYanker.scala 47:25:freechips.rocketchip.system.DefaultRV32Config.fir@71988.4 UserYanker.scala 47:25:freechips.rocketchip.system.DefaultRV32Config.fir@71990.4]
  assign _T_26_1 = QueueCompatibility_1_io_enq_ready; // @[UserYanker.scala 47:25:freechips.rocketchip.system.DefaultRV32Config.fir@71988.4 UserYanker.scala 47:25:freechips.rocketchip.system.DefaultRV32Config.fir@71991.4]
  assign _GEN_1 = 4'h1 == auto_in_ar_bits_id ? _T_26_1 : _T_26_0; // @[UserYanker.scala 48:36:freechips.rocketchip.system.DefaultRV32Config.fir@72006.4]
  assign _T_26_2 = QueueCompatibility_2_io_enq_ready; // @[UserYanker.scala 47:25:freechips.rocketchip.system.DefaultRV32Config.fir@71988.4 UserYanker.scala 47:25:freechips.rocketchip.system.DefaultRV32Config.fir@71992.4]
  assign _GEN_2 = 4'h2 == auto_in_ar_bits_id ? _T_26_2 : _GEN_1; // @[UserYanker.scala 48:36:freechips.rocketchip.system.DefaultRV32Config.fir@72006.4]
  assign _T_26_3 = QueueCompatibility_3_io_enq_ready; // @[UserYanker.scala 47:25:freechips.rocketchip.system.DefaultRV32Config.fir@71988.4 UserYanker.scala 47:25:freechips.rocketchip.system.DefaultRV32Config.fir@71993.4]
  assign _GEN_3 = 4'h3 == auto_in_ar_bits_id ? _T_26_3 : _GEN_2; // @[UserYanker.scala 48:36:freechips.rocketchip.system.DefaultRV32Config.fir@72006.4]
  assign _GEN_4 = 4'h4 == auto_in_ar_bits_id ? 1'h0 : _GEN_3; // @[UserYanker.scala 48:36:freechips.rocketchip.system.DefaultRV32Config.fir@72006.4]
  assign _GEN_5 = 4'h5 == auto_in_ar_bits_id ? 1'h0 : _GEN_4; // @[UserYanker.scala 48:36:freechips.rocketchip.system.DefaultRV32Config.fir@72006.4]
  assign _GEN_6 = 4'h6 == auto_in_ar_bits_id ? 1'h0 : _GEN_5; // @[UserYanker.scala 48:36:freechips.rocketchip.system.DefaultRV32Config.fir@72006.4]
  assign _GEN_7 = 4'h7 == auto_in_ar_bits_id ? 1'h0 : _GEN_6; // @[UserYanker.scala 48:36:freechips.rocketchip.system.DefaultRV32Config.fir@72006.4]
  assign _GEN_8 = 4'h8 == auto_in_ar_bits_id ? 1'h0 : _GEN_7; // @[UserYanker.scala 48:36:freechips.rocketchip.system.DefaultRV32Config.fir@72006.4]
  assign _GEN_9 = 4'h9 == auto_in_ar_bits_id ? 1'h0 : _GEN_8; // @[UserYanker.scala 48:36:freechips.rocketchip.system.DefaultRV32Config.fir@72006.4]
  assign _GEN_10 = 4'ha == auto_in_ar_bits_id ? 1'h0 : _GEN_9; // @[UserYanker.scala 48:36:freechips.rocketchip.system.DefaultRV32Config.fir@72006.4]
  assign _GEN_11 = 4'hb == auto_in_ar_bits_id ? 1'h0 : _GEN_10; // @[UserYanker.scala 48:36:freechips.rocketchip.system.DefaultRV32Config.fir@72006.4]
  assign _GEN_12 = 4'hc == auto_in_ar_bits_id ? 1'h0 : _GEN_11; // @[UserYanker.scala 48:36:freechips.rocketchip.system.DefaultRV32Config.fir@72006.4]
  assign _GEN_13 = 4'hd == auto_in_ar_bits_id ? 1'h0 : _GEN_12; // @[UserYanker.scala 48:36:freechips.rocketchip.system.DefaultRV32Config.fir@72006.4]
  assign _GEN_14 = 4'he == auto_in_ar_bits_id ? 1'h0 : _GEN_13; // @[UserYanker.scala 48:36:freechips.rocketchip.system.DefaultRV32Config.fir@72006.4]
  assign _GEN_15 = 4'hf == auto_in_ar_bits_id ? 1'h0 : _GEN_14; // @[UserYanker.scala 48:36:freechips.rocketchip.system.DefaultRV32Config.fir@72006.4]
  assign _T_31 = ~auto_out_r_valid; // @[UserYanker.scala 55:15:freechips.rocketchip.system.DefaultRV32Config.fir@72055.4]
  assign _T_29_0 = QueueCompatibility_io_deq_valid; // @[UserYanker.scala 53:24:freechips.rocketchip.system.DefaultRV32Config.fir@72019.4 UserYanker.scala 53:24:freechips.rocketchip.system.DefaultRV32Config.fir@72021.4]
  assign _T_29_1 = QueueCompatibility_1_io_deq_valid; // @[UserYanker.scala 53:24:freechips.rocketchip.system.DefaultRV32Config.fir@72019.4 UserYanker.scala 53:24:freechips.rocketchip.system.DefaultRV32Config.fir@72022.4]
  assign _GEN_17 = 4'h1 == auto_out_r_bits_id ? _T_29_1 : _T_29_0; // @[UserYanker.scala 55:28:freechips.rocketchip.system.DefaultRV32Config.fir@72056.4]
  assign _T_29_2 = QueueCompatibility_2_io_deq_valid; // @[UserYanker.scala 53:24:freechips.rocketchip.system.DefaultRV32Config.fir@72019.4 UserYanker.scala 53:24:freechips.rocketchip.system.DefaultRV32Config.fir@72023.4]
  assign _GEN_18 = 4'h2 == auto_out_r_bits_id ? _T_29_2 : _GEN_17; // @[UserYanker.scala 55:28:freechips.rocketchip.system.DefaultRV32Config.fir@72056.4]
  assign _T_29_3 = QueueCompatibility_3_io_deq_valid; // @[UserYanker.scala 53:24:freechips.rocketchip.system.DefaultRV32Config.fir@72019.4 UserYanker.scala 53:24:freechips.rocketchip.system.DefaultRV32Config.fir@72024.4]
  assign _GEN_19 = 4'h3 == auto_out_r_bits_id ? _T_29_3 : _GEN_18; // @[UserYanker.scala 55:28:freechips.rocketchip.system.DefaultRV32Config.fir@72056.4]
  assign _GEN_20 = 4'h4 == auto_out_r_bits_id ? 1'h0 : _GEN_19; // @[UserYanker.scala 55:28:freechips.rocketchip.system.DefaultRV32Config.fir@72056.4]
  assign _GEN_21 = 4'h5 == auto_out_r_bits_id ? 1'h0 : _GEN_20; // @[UserYanker.scala 55:28:freechips.rocketchip.system.DefaultRV32Config.fir@72056.4]
  assign _GEN_22 = 4'h6 == auto_out_r_bits_id ? 1'h0 : _GEN_21; // @[UserYanker.scala 55:28:freechips.rocketchip.system.DefaultRV32Config.fir@72056.4]
  assign _GEN_23 = 4'h7 == auto_out_r_bits_id ? 1'h0 : _GEN_22; // @[UserYanker.scala 55:28:freechips.rocketchip.system.DefaultRV32Config.fir@72056.4]
  assign _GEN_24 = 4'h8 == auto_out_r_bits_id ? 1'h0 : _GEN_23; // @[UserYanker.scala 55:28:freechips.rocketchip.system.DefaultRV32Config.fir@72056.4]
  assign _GEN_25 = 4'h9 == auto_out_r_bits_id ? 1'h0 : _GEN_24; // @[UserYanker.scala 55:28:freechips.rocketchip.system.DefaultRV32Config.fir@72056.4]
  assign _GEN_26 = 4'ha == auto_out_r_bits_id ? 1'h0 : _GEN_25; // @[UserYanker.scala 55:28:freechips.rocketchip.system.DefaultRV32Config.fir@72056.4]
  assign _GEN_27 = 4'hb == auto_out_r_bits_id ? 1'h0 : _GEN_26; // @[UserYanker.scala 55:28:freechips.rocketchip.system.DefaultRV32Config.fir@72056.4]
  assign _GEN_28 = 4'hc == auto_out_r_bits_id ? 1'h0 : _GEN_27; // @[UserYanker.scala 55:28:freechips.rocketchip.system.DefaultRV32Config.fir@72056.4]
  assign _GEN_29 = 4'hd == auto_out_r_bits_id ? 1'h0 : _GEN_28; // @[UserYanker.scala 55:28:freechips.rocketchip.system.DefaultRV32Config.fir@72056.4]
  assign _GEN_30 = 4'he == auto_out_r_bits_id ? 1'h0 : _GEN_29; // @[UserYanker.scala 55:28:freechips.rocketchip.system.DefaultRV32Config.fir@72056.4]
  assign _GEN_31 = 4'hf == auto_out_r_bits_id ? 1'h0 : _GEN_30; // @[UserYanker.scala 55:28:freechips.rocketchip.system.DefaultRV32Config.fir@72056.4]
  assign _T_32 = _T_31 | _GEN_31; // @[UserYanker.scala 55:28:freechips.rocketchip.system.DefaultRV32Config.fir@72056.4]
  assign _T_34 = _T_32 | reset; // @[UserYanker.scala 55:14:freechips.rocketchip.system.DefaultRV32Config.fir@72058.4]
  assign _T_35 = ~_T_34; // @[UserYanker.scala 55:14:freechips.rocketchip.system.DefaultRV32Config.fir@72059.4]
  assign _T_30_0_tl_state_size = QueueCompatibility_io_deq_bits_tl_state_size; // @[UserYanker.scala 54:23:freechips.rocketchip.system.DefaultRV32Config.fir@72037.4 UserYanker.scala 54:23:freechips.rocketchip.system.DefaultRV32Config.fir@72039.4]
  assign _T_30_0_tl_state_source = QueueCompatibility_io_deq_bits_tl_state_source; // @[UserYanker.scala 54:23:freechips.rocketchip.system.DefaultRV32Config.fir@72037.4 UserYanker.scala 54:23:freechips.rocketchip.system.DefaultRV32Config.fir@72039.4]
  assign _T_30_1_tl_state_size = QueueCompatibility_1_io_deq_bits_tl_state_size; // @[UserYanker.scala 54:23:freechips.rocketchip.system.DefaultRV32Config.fir@72037.4 UserYanker.scala 54:23:freechips.rocketchip.system.DefaultRV32Config.fir@72040.4]
  assign _GEN_34 = 4'h1 == auto_out_r_bits_id ? _T_30_1_tl_state_size : _T_30_0_tl_state_size; // @[BundleMap.scala 248:19:freechips.rocketchip.system.DefaultRV32Config.fir@72072.4]
  assign _T_30_1_tl_state_source = QueueCompatibility_1_io_deq_bits_tl_state_source; // @[UserYanker.scala 54:23:freechips.rocketchip.system.DefaultRV32Config.fir@72037.4 UserYanker.scala 54:23:freechips.rocketchip.system.DefaultRV32Config.fir@72040.4]
  assign _GEN_35 = 4'h1 == auto_out_r_bits_id ? _T_30_1_tl_state_source : _T_30_0_tl_state_source; // @[BundleMap.scala 248:19:freechips.rocketchip.system.DefaultRV32Config.fir@72072.4]
  assign _T_30_2_tl_state_size = QueueCompatibility_2_io_deq_bits_tl_state_size; // @[UserYanker.scala 54:23:freechips.rocketchip.system.DefaultRV32Config.fir@72037.4 UserYanker.scala 54:23:freechips.rocketchip.system.DefaultRV32Config.fir@72041.4]
  assign _GEN_36 = 4'h2 == auto_out_r_bits_id ? _T_30_2_tl_state_size : _GEN_34; // @[BundleMap.scala 248:19:freechips.rocketchip.system.DefaultRV32Config.fir@72072.4]
  assign _T_30_2_tl_state_source = QueueCompatibility_2_io_deq_bits_tl_state_source; // @[UserYanker.scala 54:23:freechips.rocketchip.system.DefaultRV32Config.fir@72037.4 UserYanker.scala 54:23:freechips.rocketchip.system.DefaultRV32Config.fir@72041.4]
  assign _GEN_37 = 4'h2 == auto_out_r_bits_id ? _T_30_2_tl_state_source : _GEN_35; // @[BundleMap.scala 248:19:freechips.rocketchip.system.DefaultRV32Config.fir@72072.4]
  assign _T_30_3_tl_state_size = QueueCompatibility_3_io_deq_bits_tl_state_size; // @[UserYanker.scala 54:23:freechips.rocketchip.system.DefaultRV32Config.fir@72037.4 UserYanker.scala 54:23:freechips.rocketchip.system.DefaultRV32Config.fir@72042.4]
  assign _GEN_38 = 4'h3 == auto_out_r_bits_id ? _T_30_3_tl_state_size : _GEN_36; // @[BundleMap.scala 248:19:freechips.rocketchip.system.DefaultRV32Config.fir@72072.4]
  assign _T_30_3_tl_state_source = QueueCompatibility_3_io_deq_bits_tl_state_source; // @[UserYanker.scala 54:23:freechips.rocketchip.system.DefaultRV32Config.fir@72037.4 UserYanker.scala 54:23:freechips.rocketchip.system.DefaultRV32Config.fir@72042.4]
  assign _GEN_39 = 4'h3 == auto_out_r_bits_id ? _T_30_3_tl_state_source : _GEN_37; // @[BundleMap.scala 248:19:freechips.rocketchip.system.DefaultRV32Config.fir@72072.4]
  assign _GEN_40 = 4'h4 == auto_out_r_bits_id ? 4'h0 : _GEN_38; // @[BundleMap.scala 248:19:freechips.rocketchip.system.DefaultRV32Config.fir@72072.4]
  assign _GEN_41 = 4'h4 == auto_out_r_bits_id ? 2'h0 : _GEN_39; // @[BundleMap.scala 248:19:freechips.rocketchip.system.DefaultRV32Config.fir@72072.4]
  assign _GEN_42 = 4'h5 == auto_out_r_bits_id ? 4'h0 : _GEN_40; // @[BundleMap.scala 248:19:freechips.rocketchip.system.DefaultRV32Config.fir@72072.4]
  assign _GEN_43 = 4'h5 == auto_out_r_bits_id ? 2'h0 : _GEN_41; // @[BundleMap.scala 248:19:freechips.rocketchip.system.DefaultRV32Config.fir@72072.4]
  assign _GEN_44 = 4'h6 == auto_out_r_bits_id ? 4'h0 : _GEN_42; // @[BundleMap.scala 248:19:freechips.rocketchip.system.DefaultRV32Config.fir@72072.4]
  assign _GEN_45 = 4'h6 == auto_out_r_bits_id ? 2'h0 : _GEN_43; // @[BundleMap.scala 248:19:freechips.rocketchip.system.DefaultRV32Config.fir@72072.4]
  assign _GEN_46 = 4'h7 == auto_out_r_bits_id ? 4'h0 : _GEN_44; // @[BundleMap.scala 248:19:freechips.rocketchip.system.DefaultRV32Config.fir@72072.4]
  assign _GEN_47 = 4'h7 == auto_out_r_bits_id ? 2'h0 : _GEN_45; // @[BundleMap.scala 248:19:freechips.rocketchip.system.DefaultRV32Config.fir@72072.4]
  assign _GEN_48 = 4'h8 == auto_out_r_bits_id ? 4'h0 : _GEN_46; // @[BundleMap.scala 248:19:freechips.rocketchip.system.DefaultRV32Config.fir@72072.4]
  assign _GEN_49 = 4'h8 == auto_out_r_bits_id ? 2'h0 : _GEN_47; // @[BundleMap.scala 248:19:freechips.rocketchip.system.DefaultRV32Config.fir@72072.4]
  assign _GEN_50 = 4'h9 == auto_out_r_bits_id ? 4'h0 : _GEN_48; // @[BundleMap.scala 248:19:freechips.rocketchip.system.DefaultRV32Config.fir@72072.4]
  assign _GEN_51 = 4'h9 == auto_out_r_bits_id ? 2'h0 : _GEN_49; // @[BundleMap.scala 248:19:freechips.rocketchip.system.DefaultRV32Config.fir@72072.4]
  assign _GEN_52 = 4'ha == auto_out_r_bits_id ? 4'h0 : _GEN_50; // @[BundleMap.scala 248:19:freechips.rocketchip.system.DefaultRV32Config.fir@72072.4]
  assign _GEN_53 = 4'ha == auto_out_r_bits_id ? 2'h0 : _GEN_51; // @[BundleMap.scala 248:19:freechips.rocketchip.system.DefaultRV32Config.fir@72072.4]
  assign _GEN_54 = 4'hb == auto_out_r_bits_id ? 4'h0 : _GEN_52; // @[BundleMap.scala 248:19:freechips.rocketchip.system.DefaultRV32Config.fir@72072.4]
  assign _GEN_55 = 4'hb == auto_out_r_bits_id ? 2'h0 : _GEN_53; // @[BundleMap.scala 248:19:freechips.rocketchip.system.DefaultRV32Config.fir@72072.4]
  assign _GEN_56 = 4'hc == auto_out_r_bits_id ? 4'h0 : _GEN_54; // @[BundleMap.scala 248:19:freechips.rocketchip.system.DefaultRV32Config.fir@72072.4]
  assign _GEN_57 = 4'hc == auto_out_r_bits_id ? 2'h0 : _GEN_55; // @[BundleMap.scala 248:19:freechips.rocketchip.system.DefaultRV32Config.fir@72072.4]
  assign _GEN_58 = 4'hd == auto_out_r_bits_id ? 4'h0 : _GEN_56; // @[BundleMap.scala 248:19:freechips.rocketchip.system.DefaultRV32Config.fir@72072.4]
  assign _GEN_59 = 4'hd == auto_out_r_bits_id ? 2'h0 : _GEN_57; // @[BundleMap.scala 248:19:freechips.rocketchip.system.DefaultRV32Config.fir@72072.4]
  assign _GEN_60 = 4'he == auto_out_r_bits_id ? 4'h0 : _GEN_58; // @[BundleMap.scala 248:19:freechips.rocketchip.system.DefaultRV32Config.fir@72072.4]
  assign _GEN_61 = 4'he == auto_out_r_bits_id ? 2'h0 : _GEN_59; // @[BundleMap.scala 248:19:freechips.rocketchip.system.DefaultRV32Config.fir@72072.4]
  assign _T_37 = 16'h1 << auto_in_ar_bits_id; // @[OneHot.scala 65:12:freechips.rocketchip.system.DefaultRV32Config.fir@72075.4]
  assign _T_56 = 16'h1 << auto_out_r_bits_id; // @[OneHot.scala 65:12:freechips.rocketchip.system.DefaultRV32Config.fir@72094.4]
  assign _T_74 = auto_out_r_valid & auto_in_r_ready; // @[UserYanker.scala 62:37:freechips.rocketchip.system.DefaultRV32Config.fir@72112.4]
  assign _T_75 = _T_74 & _T_56[0]; // @[UserYanker.scala 62:53:freechips.rocketchip.system.DefaultRV32Config.fir@72113.4]
  assign _T_77 = auto_in_ar_valid & auto_out_ar_ready; // @[UserYanker.scala 63:37:freechips.rocketchip.system.DefaultRV32Config.fir@72116.4]
  assign _T_80 = _T_74 & _T_56[1]; // @[UserYanker.scala 62:53:freechips.rocketchip.system.DefaultRV32Config.fir@72122.4]
  assign _T_85 = _T_74 & _T_56[2]; // @[UserYanker.scala 62:53:freechips.rocketchip.system.DefaultRV32Config.fir@72131.4]
  assign _T_90 = _T_74 & _T_56[3]; // @[UserYanker.scala 62:53:freechips.rocketchip.system.DefaultRV32Config.fir@72140.4]
  assign _T_154_0 = QueueCompatibility_4_io_enq_ready; // @[UserYanker.scala 68:25:freechips.rocketchip.system.DefaultRV32Config.fir@72256.4 UserYanker.scala 68:25:freechips.rocketchip.system.DefaultRV32Config.fir@72258.4]
  assign _T_154_1 = QueueCompatibility_5_io_enq_ready; // @[UserYanker.scala 68:25:freechips.rocketchip.system.DefaultRV32Config.fir@72256.4 UserYanker.scala 68:25:freechips.rocketchip.system.DefaultRV32Config.fir@72259.4]
  assign _GEN_65 = 4'h1 == auto_in_aw_bits_id ? _T_154_1 : _T_154_0; // @[UserYanker.scala 69:36:freechips.rocketchip.system.DefaultRV32Config.fir@72274.4]
  assign _T_154_2 = QueueCompatibility_6_io_enq_ready; // @[UserYanker.scala 68:25:freechips.rocketchip.system.DefaultRV32Config.fir@72256.4 UserYanker.scala 68:25:freechips.rocketchip.system.DefaultRV32Config.fir@72260.4]
  assign _GEN_66 = 4'h2 == auto_in_aw_bits_id ? _T_154_2 : _GEN_65; // @[UserYanker.scala 69:36:freechips.rocketchip.system.DefaultRV32Config.fir@72274.4]
  assign _T_154_3 = QueueCompatibility_7_io_enq_ready; // @[UserYanker.scala 68:25:freechips.rocketchip.system.DefaultRV32Config.fir@72256.4 UserYanker.scala 68:25:freechips.rocketchip.system.DefaultRV32Config.fir@72261.4]
  assign _GEN_67 = 4'h3 == auto_in_aw_bits_id ? _T_154_3 : _GEN_66; // @[UserYanker.scala 69:36:freechips.rocketchip.system.DefaultRV32Config.fir@72274.4]
  assign _GEN_68 = 4'h4 == auto_in_aw_bits_id ? 1'h0 : _GEN_67; // @[UserYanker.scala 69:36:freechips.rocketchip.system.DefaultRV32Config.fir@72274.4]
  assign _GEN_69 = 4'h5 == auto_in_aw_bits_id ? 1'h0 : _GEN_68; // @[UserYanker.scala 69:36:freechips.rocketchip.system.DefaultRV32Config.fir@72274.4]
  assign _GEN_70 = 4'h6 == auto_in_aw_bits_id ? 1'h0 : _GEN_69; // @[UserYanker.scala 69:36:freechips.rocketchip.system.DefaultRV32Config.fir@72274.4]
  assign _GEN_71 = 4'h7 == auto_in_aw_bits_id ? 1'h0 : _GEN_70; // @[UserYanker.scala 69:36:freechips.rocketchip.system.DefaultRV32Config.fir@72274.4]
  assign _GEN_72 = 4'h8 == auto_in_aw_bits_id ? 1'h0 : _GEN_71; // @[UserYanker.scala 69:36:freechips.rocketchip.system.DefaultRV32Config.fir@72274.4]
  assign _GEN_73 = 4'h9 == auto_in_aw_bits_id ? 1'h0 : _GEN_72; // @[UserYanker.scala 69:36:freechips.rocketchip.system.DefaultRV32Config.fir@72274.4]
  assign _GEN_74 = 4'ha == auto_in_aw_bits_id ? 1'h0 : _GEN_73; // @[UserYanker.scala 69:36:freechips.rocketchip.system.DefaultRV32Config.fir@72274.4]
  assign _GEN_75 = 4'hb == auto_in_aw_bits_id ? 1'h0 : _GEN_74; // @[UserYanker.scala 69:36:freechips.rocketchip.system.DefaultRV32Config.fir@72274.4]
  assign _GEN_76 = 4'hc == auto_in_aw_bits_id ? 1'h0 : _GEN_75; // @[UserYanker.scala 69:36:freechips.rocketchip.system.DefaultRV32Config.fir@72274.4]
  assign _GEN_77 = 4'hd == auto_in_aw_bits_id ? 1'h0 : _GEN_76; // @[UserYanker.scala 69:36:freechips.rocketchip.system.DefaultRV32Config.fir@72274.4]
  assign _GEN_78 = 4'he == auto_in_aw_bits_id ? 1'h0 : _GEN_77; // @[UserYanker.scala 69:36:freechips.rocketchip.system.DefaultRV32Config.fir@72274.4]
  assign _GEN_79 = 4'hf == auto_in_aw_bits_id ? 1'h0 : _GEN_78; // @[UserYanker.scala 69:36:freechips.rocketchip.system.DefaultRV32Config.fir@72274.4]
  assign _T_159 = ~auto_out_b_valid; // @[UserYanker.scala 76:15:freechips.rocketchip.system.DefaultRV32Config.fir@72323.4]
  assign _T_157_0 = QueueCompatibility_4_io_deq_valid; // @[UserYanker.scala 74:24:freechips.rocketchip.system.DefaultRV32Config.fir@72287.4 UserYanker.scala 74:24:freechips.rocketchip.system.DefaultRV32Config.fir@72289.4]
  assign _T_157_1 = QueueCompatibility_5_io_deq_valid; // @[UserYanker.scala 74:24:freechips.rocketchip.system.DefaultRV32Config.fir@72287.4 UserYanker.scala 74:24:freechips.rocketchip.system.DefaultRV32Config.fir@72290.4]
  assign _GEN_81 = 4'h1 == auto_out_b_bits_id ? _T_157_1 : _T_157_0; // @[UserYanker.scala 76:28:freechips.rocketchip.system.DefaultRV32Config.fir@72324.4]
  assign _T_157_2 = QueueCompatibility_6_io_deq_valid; // @[UserYanker.scala 74:24:freechips.rocketchip.system.DefaultRV32Config.fir@72287.4 UserYanker.scala 74:24:freechips.rocketchip.system.DefaultRV32Config.fir@72291.4]
  assign _GEN_82 = 4'h2 == auto_out_b_bits_id ? _T_157_2 : _GEN_81; // @[UserYanker.scala 76:28:freechips.rocketchip.system.DefaultRV32Config.fir@72324.4]
  assign _T_157_3 = QueueCompatibility_7_io_deq_valid; // @[UserYanker.scala 74:24:freechips.rocketchip.system.DefaultRV32Config.fir@72287.4 UserYanker.scala 74:24:freechips.rocketchip.system.DefaultRV32Config.fir@72292.4]
  assign _GEN_83 = 4'h3 == auto_out_b_bits_id ? _T_157_3 : _GEN_82; // @[UserYanker.scala 76:28:freechips.rocketchip.system.DefaultRV32Config.fir@72324.4]
  assign _GEN_84 = 4'h4 == auto_out_b_bits_id ? 1'h0 : _GEN_83; // @[UserYanker.scala 76:28:freechips.rocketchip.system.DefaultRV32Config.fir@72324.4]
  assign _GEN_85 = 4'h5 == auto_out_b_bits_id ? 1'h0 : _GEN_84; // @[UserYanker.scala 76:28:freechips.rocketchip.system.DefaultRV32Config.fir@72324.4]
  assign _GEN_86 = 4'h6 == auto_out_b_bits_id ? 1'h0 : _GEN_85; // @[UserYanker.scala 76:28:freechips.rocketchip.system.DefaultRV32Config.fir@72324.4]
  assign _GEN_87 = 4'h7 == auto_out_b_bits_id ? 1'h0 : _GEN_86; // @[UserYanker.scala 76:28:freechips.rocketchip.system.DefaultRV32Config.fir@72324.4]
  assign _GEN_88 = 4'h8 == auto_out_b_bits_id ? 1'h0 : _GEN_87; // @[UserYanker.scala 76:28:freechips.rocketchip.system.DefaultRV32Config.fir@72324.4]
  assign _GEN_89 = 4'h9 == auto_out_b_bits_id ? 1'h0 : _GEN_88; // @[UserYanker.scala 76:28:freechips.rocketchip.system.DefaultRV32Config.fir@72324.4]
  assign _GEN_90 = 4'ha == auto_out_b_bits_id ? 1'h0 : _GEN_89; // @[UserYanker.scala 76:28:freechips.rocketchip.system.DefaultRV32Config.fir@72324.4]
  assign _GEN_91 = 4'hb == auto_out_b_bits_id ? 1'h0 : _GEN_90; // @[UserYanker.scala 76:28:freechips.rocketchip.system.DefaultRV32Config.fir@72324.4]
  assign _GEN_92 = 4'hc == auto_out_b_bits_id ? 1'h0 : _GEN_91; // @[UserYanker.scala 76:28:freechips.rocketchip.system.DefaultRV32Config.fir@72324.4]
  assign _GEN_93 = 4'hd == auto_out_b_bits_id ? 1'h0 : _GEN_92; // @[UserYanker.scala 76:28:freechips.rocketchip.system.DefaultRV32Config.fir@72324.4]
  assign _GEN_94 = 4'he == auto_out_b_bits_id ? 1'h0 : _GEN_93; // @[UserYanker.scala 76:28:freechips.rocketchip.system.DefaultRV32Config.fir@72324.4]
  assign _GEN_95 = 4'hf == auto_out_b_bits_id ? 1'h0 : _GEN_94; // @[UserYanker.scala 76:28:freechips.rocketchip.system.DefaultRV32Config.fir@72324.4]
  assign _T_160 = _T_159 | _GEN_95; // @[UserYanker.scala 76:28:freechips.rocketchip.system.DefaultRV32Config.fir@72324.4]
  assign _T_162 = _T_160 | reset; // @[UserYanker.scala 76:14:freechips.rocketchip.system.DefaultRV32Config.fir@72326.4]
  assign _T_163 = ~_T_162; // @[UserYanker.scala 76:14:freechips.rocketchip.system.DefaultRV32Config.fir@72327.4]
  assign _T_158_0_tl_state_size = QueueCompatibility_4_io_deq_bits_tl_state_size; // @[UserYanker.scala 75:23:freechips.rocketchip.system.DefaultRV32Config.fir@72305.4 UserYanker.scala 75:23:freechips.rocketchip.system.DefaultRV32Config.fir@72307.4]
  assign _T_158_0_tl_state_source = QueueCompatibility_4_io_deq_bits_tl_state_source; // @[UserYanker.scala 75:23:freechips.rocketchip.system.DefaultRV32Config.fir@72305.4 UserYanker.scala 75:23:freechips.rocketchip.system.DefaultRV32Config.fir@72307.4]
  assign _T_158_1_tl_state_size = QueueCompatibility_5_io_deq_bits_tl_state_size; // @[UserYanker.scala 75:23:freechips.rocketchip.system.DefaultRV32Config.fir@72305.4 UserYanker.scala 75:23:freechips.rocketchip.system.DefaultRV32Config.fir@72308.4]
  assign _GEN_98 = 4'h1 == auto_out_b_bits_id ? _T_158_1_tl_state_size : _T_158_0_tl_state_size; // @[BundleMap.scala 248:19:freechips.rocketchip.system.DefaultRV32Config.fir@72338.4]
  assign _T_158_1_tl_state_source = QueueCompatibility_5_io_deq_bits_tl_state_source; // @[UserYanker.scala 75:23:freechips.rocketchip.system.DefaultRV32Config.fir@72305.4 UserYanker.scala 75:23:freechips.rocketchip.system.DefaultRV32Config.fir@72308.4]
  assign _GEN_99 = 4'h1 == auto_out_b_bits_id ? _T_158_1_tl_state_source : _T_158_0_tl_state_source; // @[BundleMap.scala 248:19:freechips.rocketchip.system.DefaultRV32Config.fir@72338.4]
  assign _T_158_2_tl_state_size = QueueCompatibility_6_io_deq_bits_tl_state_size; // @[UserYanker.scala 75:23:freechips.rocketchip.system.DefaultRV32Config.fir@72305.4 UserYanker.scala 75:23:freechips.rocketchip.system.DefaultRV32Config.fir@72309.4]
  assign _GEN_100 = 4'h2 == auto_out_b_bits_id ? _T_158_2_tl_state_size : _GEN_98; // @[BundleMap.scala 248:19:freechips.rocketchip.system.DefaultRV32Config.fir@72338.4]
  assign _T_158_2_tl_state_source = QueueCompatibility_6_io_deq_bits_tl_state_source; // @[UserYanker.scala 75:23:freechips.rocketchip.system.DefaultRV32Config.fir@72305.4 UserYanker.scala 75:23:freechips.rocketchip.system.DefaultRV32Config.fir@72309.4]
  assign _GEN_101 = 4'h2 == auto_out_b_bits_id ? _T_158_2_tl_state_source : _GEN_99; // @[BundleMap.scala 248:19:freechips.rocketchip.system.DefaultRV32Config.fir@72338.4]
  assign _T_158_3_tl_state_size = QueueCompatibility_7_io_deq_bits_tl_state_size; // @[UserYanker.scala 75:23:freechips.rocketchip.system.DefaultRV32Config.fir@72305.4 UserYanker.scala 75:23:freechips.rocketchip.system.DefaultRV32Config.fir@72310.4]
  assign _GEN_102 = 4'h3 == auto_out_b_bits_id ? _T_158_3_tl_state_size : _GEN_100; // @[BundleMap.scala 248:19:freechips.rocketchip.system.DefaultRV32Config.fir@72338.4]
  assign _T_158_3_tl_state_source = QueueCompatibility_7_io_deq_bits_tl_state_source; // @[UserYanker.scala 75:23:freechips.rocketchip.system.DefaultRV32Config.fir@72305.4 UserYanker.scala 75:23:freechips.rocketchip.system.DefaultRV32Config.fir@72310.4]
  assign _GEN_103 = 4'h3 == auto_out_b_bits_id ? _T_158_3_tl_state_source : _GEN_101; // @[BundleMap.scala 248:19:freechips.rocketchip.system.DefaultRV32Config.fir@72338.4]
  assign _GEN_104 = 4'h4 == auto_out_b_bits_id ? 4'h0 : _GEN_102; // @[BundleMap.scala 248:19:freechips.rocketchip.system.DefaultRV32Config.fir@72338.4]
  assign _GEN_105 = 4'h4 == auto_out_b_bits_id ? 2'h0 : _GEN_103; // @[BundleMap.scala 248:19:freechips.rocketchip.system.DefaultRV32Config.fir@72338.4]
  assign _GEN_106 = 4'h5 == auto_out_b_bits_id ? 4'h0 : _GEN_104; // @[BundleMap.scala 248:19:freechips.rocketchip.system.DefaultRV32Config.fir@72338.4]
  assign _GEN_107 = 4'h5 == auto_out_b_bits_id ? 2'h0 : _GEN_105; // @[BundleMap.scala 248:19:freechips.rocketchip.system.DefaultRV32Config.fir@72338.4]
  assign _GEN_108 = 4'h6 == auto_out_b_bits_id ? 4'h0 : _GEN_106; // @[BundleMap.scala 248:19:freechips.rocketchip.system.DefaultRV32Config.fir@72338.4]
  assign _GEN_109 = 4'h6 == auto_out_b_bits_id ? 2'h0 : _GEN_107; // @[BundleMap.scala 248:19:freechips.rocketchip.system.DefaultRV32Config.fir@72338.4]
  assign _GEN_110 = 4'h7 == auto_out_b_bits_id ? 4'h0 : _GEN_108; // @[BundleMap.scala 248:19:freechips.rocketchip.system.DefaultRV32Config.fir@72338.4]
  assign _GEN_111 = 4'h7 == auto_out_b_bits_id ? 2'h0 : _GEN_109; // @[BundleMap.scala 248:19:freechips.rocketchip.system.DefaultRV32Config.fir@72338.4]
  assign _GEN_112 = 4'h8 == auto_out_b_bits_id ? 4'h0 : _GEN_110; // @[BundleMap.scala 248:19:freechips.rocketchip.system.DefaultRV32Config.fir@72338.4]
  assign _GEN_113 = 4'h8 == auto_out_b_bits_id ? 2'h0 : _GEN_111; // @[BundleMap.scala 248:19:freechips.rocketchip.system.DefaultRV32Config.fir@72338.4]
  assign _GEN_114 = 4'h9 == auto_out_b_bits_id ? 4'h0 : _GEN_112; // @[BundleMap.scala 248:19:freechips.rocketchip.system.DefaultRV32Config.fir@72338.4]
  assign _GEN_115 = 4'h9 == auto_out_b_bits_id ? 2'h0 : _GEN_113; // @[BundleMap.scala 248:19:freechips.rocketchip.system.DefaultRV32Config.fir@72338.4]
  assign _GEN_116 = 4'ha == auto_out_b_bits_id ? 4'h0 : _GEN_114; // @[BundleMap.scala 248:19:freechips.rocketchip.system.DefaultRV32Config.fir@72338.4]
  assign _GEN_117 = 4'ha == auto_out_b_bits_id ? 2'h0 : _GEN_115; // @[BundleMap.scala 248:19:freechips.rocketchip.system.DefaultRV32Config.fir@72338.4]
  assign _GEN_118 = 4'hb == auto_out_b_bits_id ? 4'h0 : _GEN_116; // @[BundleMap.scala 248:19:freechips.rocketchip.system.DefaultRV32Config.fir@72338.4]
  assign _GEN_119 = 4'hb == auto_out_b_bits_id ? 2'h0 : _GEN_117; // @[BundleMap.scala 248:19:freechips.rocketchip.system.DefaultRV32Config.fir@72338.4]
  assign _GEN_120 = 4'hc == auto_out_b_bits_id ? 4'h0 : _GEN_118; // @[BundleMap.scala 248:19:freechips.rocketchip.system.DefaultRV32Config.fir@72338.4]
  assign _GEN_121 = 4'hc == auto_out_b_bits_id ? 2'h0 : _GEN_119; // @[BundleMap.scala 248:19:freechips.rocketchip.system.DefaultRV32Config.fir@72338.4]
  assign _GEN_122 = 4'hd == auto_out_b_bits_id ? 4'h0 : _GEN_120; // @[BundleMap.scala 248:19:freechips.rocketchip.system.DefaultRV32Config.fir@72338.4]
  assign _GEN_123 = 4'hd == auto_out_b_bits_id ? 2'h0 : _GEN_121; // @[BundleMap.scala 248:19:freechips.rocketchip.system.DefaultRV32Config.fir@72338.4]
  assign _GEN_124 = 4'he == auto_out_b_bits_id ? 4'h0 : _GEN_122; // @[BundleMap.scala 248:19:freechips.rocketchip.system.DefaultRV32Config.fir@72338.4]
  assign _GEN_125 = 4'he == auto_out_b_bits_id ? 2'h0 : _GEN_123; // @[BundleMap.scala 248:19:freechips.rocketchip.system.DefaultRV32Config.fir@72338.4]
  assign _T_165 = 16'h1 << auto_in_aw_bits_id; // @[OneHot.scala 65:12:freechips.rocketchip.system.DefaultRV32Config.fir@72341.4]
  assign _T_184 = 16'h1 << auto_out_b_bits_id; // @[OneHot.scala 65:12:freechips.rocketchip.system.DefaultRV32Config.fir@72360.4]
  assign _T_202 = auto_out_b_valid & auto_in_b_ready; // @[UserYanker.scala 83:37:freechips.rocketchip.system.DefaultRV32Config.fir@72378.4]
  assign _T_204 = auto_in_aw_valid & auto_out_aw_ready; // @[UserYanker.scala 84:37:freechips.rocketchip.system.DefaultRV32Config.fir@72381.4]
  assign auto_in_aw_ready = auto_out_aw_ready & _GEN_79; // @[LazyModule.scala 303:16:freechips.rocketchip.system.DefaultRV32Config.fir@71907.4]
  assign auto_in_w_ready = auto_out_w_ready; // @[LazyModule.scala 303:16:freechips.rocketchip.system.DefaultRV32Config.fir@71907.4]
  assign auto_in_b_valid = auto_out_b_valid; // @[LazyModule.scala 303:16:freechips.rocketchip.system.DefaultRV32Config.fir@71907.4]
  assign auto_in_b_bits_id = auto_out_b_bits_id; // @[LazyModule.scala 303:16:freechips.rocketchip.system.DefaultRV32Config.fir@71907.4]
  assign auto_in_b_bits_resp = auto_out_b_bits_resp; // @[LazyModule.scala 303:16:freechips.rocketchip.system.DefaultRV32Config.fir@71907.4]
  assign auto_in_b_bits_echo_tl_state_size = 4'hf == auto_out_b_bits_id ? 4'h0 : _GEN_124; // @[LazyModule.scala 303:16:freechips.rocketchip.system.DefaultRV32Config.fir@71907.4]
  assign auto_in_b_bits_echo_tl_state_source = 4'hf == auto_out_b_bits_id ? 2'h0 : _GEN_125; // @[LazyModule.scala 303:16:freechips.rocketchip.system.DefaultRV32Config.fir@71907.4]
  assign auto_in_ar_ready = auto_out_ar_ready & _GEN_15; // @[LazyModule.scala 303:16:freechips.rocketchip.system.DefaultRV32Config.fir@71907.4]
  assign auto_in_r_valid = auto_out_r_valid; // @[LazyModule.scala 303:16:freechips.rocketchip.system.DefaultRV32Config.fir@71907.4]
  assign auto_in_r_bits_id = auto_out_r_bits_id; // @[LazyModule.scala 303:16:freechips.rocketchip.system.DefaultRV32Config.fir@71907.4]
  assign auto_in_r_bits_data = auto_out_r_bits_data; // @[LazyModule.scala 303:16:freechips.rocketchip.system.DefaultRV32Config.fir@71907.4]
  assign auto_in_r_bits_resp = auto_out_r_bits_resp; // @[LazyModule.scala 303:16:freechips.rocketchip.system.DefaultRV32Config.fir@71907.4]
  assign auto_in_r_bits_echo_tl_state_size = 4'hf == auto_out_r_bits_id ? 4'h0 : _GEN_60; // @[LazyModule.scala 303:16:freechips.rocketchip.system.DefaultRV32Config.fir@71907.4]
  assign auto_in_r_bits_echo_tl_state_source = 4'hf == auto_out_r_bits_id ? 2'h0 : _GEN_61; // @[LazyModule.scala 303:16:freechips.rocketchip.system.DefaultRV32Config.fir@71907.4]
  assign auto_in_r_bits_last = auto_out_r_bits_last; // @[LazyModule.scala 303:16:freechips.rocketchip.system.DefaultRV32Config.fir@71907.4]
  assign auto_out_aw_valid = auto_in_aw_valid & _GEN_79; // @[LazyModule.scala 305:12:freechips.rocketchip.system.DefaultRV32Config.fir@71906.4]
  assign auto_out_aw_bits_id = auto_in_aw_bits_id; // @[LazyModule.scala 305:12:freechips.rocketchip.system.DefaultRV32Config.fir@71906.4]
  assign auto_out_aw_bits_addr = auto_in_aw_bits_addr; // @[LazyModule.scala 305:12:freechips.rocketchip.system.DefaultRV32Config.fir@71906.4]
  assign auto_out_aw_bits_len = auto_in_aw_bits_len; // @[LazyModule.scala 305:12:freechips.rocketchip.system.DefaultRV32Config.fir@71906.4]
  assign auto_out_aw_bits_size = auto_in_aw_bits_size; // @[LazyModule.scala 305:12:freechips.rocketchip.system.DefaultRV32Config.fir@71906.4]
  assign auto_out_aw_bits_burst = auto_in_aw_bits_burst; // @[LazyModule.scala 305:12:freechips.rocketchip.system.DefaultRV32Config.fir@71906.4]
  assign auto_out_aw_bits_lock = auto_in_aw_bits_lock; // @[LazyModule.scala 305:12:freechips.rocketchip.system.DefaultRV32Config.fir@71906.4]
  assign auto_out_aw_bits_cache = auto_in_aw_bits_cache; // @[LazyModule.scala 305:12:freechips.rocketchip.system.DefaultRV32Config.fir@71906.4]
  assign auto_out_aw_bits_prot = auto_in_aw_bits_prot; // @[LazyModule.scala 305:12:freechips.rocketchip.system.DefaultRV32Config.fir@71906.4]
  assign auto_out_aw_bits_qos = auto_in_aw_bits_qos; // @[LazyModule.scala 305:12:freechips.rocketchip.system.DefaultRV32Config.fir@71906.4]
  assign auto_out_w_valid = auto_in_w_valid; // @[LazyModule.scala 305:12:freechips.rocketchip.system.DefaultRV32Config.fir@71906.4]
  assign auto_out_w_bits_data = auto_in_w_bits_data; // @[LazyModule.scala 305:12:freechips.rocketchip.system.DefaultRV32Config.fir@71906.4]
  assign auto_out_w_bits_strb = auto_in_w_bits_strb; // @[LazyModule.scala 305:12:freechips.rocketchip.system.DefaultRV32Config.fir@71906.4]
  assign auto_out_w_bits_last = auto_in_w_bits_last; // @[LazyModule.scala 305:12:freechips.rocketchip.system.DefaultRV32Config.fir@71906.4]
  assign auto_out_b_ready = auto_in_b_ready; // @[LazyModule.scala 305:12:freechips.rocketchip.system.DefaultRV32Config.fir@71906.4]
  assign auto_out_ar_valid = auto_in_ar_valid & _GEN_15; // @[LazyModule.scala 305:12:freechips.rocketchip.system.DefaultRV32Config.fir@71906.4]
  assign auto_out_ar_bits_id = auto_in_ar_bits_id; // @[LazyModule.scala 305:12:freechips.rocketchip.system.DefaultRV32Config.fir@71906.4]
  assign auto_out_ar_bits_addr = auto_in_ar_bits_addr; // @[LazyModule.scala 305:12:freechips.rocketchip.system.DefaultRV32Config.fir@71906.4]
  assign auto_out_ar_bits_len = auto_in_ar_bits_len; // @[LazyModule.scala 305:12:freechips.rocketchip.system.DefaultRV32Config.fir@71906.4]
  assign auto_out_ar_bits_size = auto_in_ar_bits_size; // @[LazyModule.scala 305:12:freechips.rocketchip.system.DefaultRV32Config.fir@71906.4]
  assign auto_out_ar_bits_burst = auto_in_ar_bits_burst; // @[LazyModule.scala 305:12:freechips.rocketchip.system.DefaultRV32Config.fir@71906.4]
  assign auto_out_ar_bits_lock = auto_in_ar_bits_lock; // @[LazyModule.scala 305:12:freechips.rocketchip.system.DefaultRV32Config.fir@71906.4]
  assign auto_out_ar_bits_cache = auto_in_ar_bits_cache; // @[LazyModule.scala 305:12:freechips.rocketchip.system.DefaultRV32Config.fir@71906.4]
  assign auto_out_ar_bits_prot = auto_in_ar_bits_prot; // @[LazyModule.scala 305:12:freechips.rocketchip.system.DefaultRV32Config.fir@71906.4]
  assign auto_out_ar_bits_qos = auto_in_ar_bits_qos; // @[LazyModule.scala 305:12:freechips.rocketchip.system.DefaultRV32Config.fir@71906.4]
  assign auto_out_r_ready = auto_in_r_ready; // @[LazyModule.scala 305:12:freechips.rocketchip.system.DefaultRV32Config.fir@71906.4]
  assign QueueCompatibility_clock = clock; // @[:freechips.rocketchip.system.DefaultRV32Config.fir@71910.4]
  assign QueueCompatibility_reset = reset; // @[:freechips.rocketchip.system.DefaultRV32Config.fir@71911.4]
  assign QueueCompatibility_io_enq_valid = _T_77 & _T_37[0]; // @[UserYanker.scala 63:21:freechips.rocketchip.system.DefaultRV32Config.fir@72118.4]
  assign QueueCompatibility_io_enq_bits_tl_state_size = auto_in_ar_bits_echo_tl_state_size; // @[BundleMap.scala 248:19:freechips.rocketchip.system.DefaultRV32Config.fir@72120.4]
  assign QueueCompatibility_io_enq_bits_tl_state_source = auto_in_ar_bits_echo_tl_state_source; // @[BundleMap.scala 248:19:freechips.rocketchip.system.DefaultRV32Config.fir@72119.4]
  assign QueueCompatibility_io_deq_ready = _T_75 & auto_out_r_bits_last; // @[UserYanker.scala 62:21:freechips.rocketchip.system.DefaultRV32Config.fir@72115.4]
  assign QueueCompatibility_1_clock = clock; // @[:freechips.rocketchip.system.DefaultRV32Config.fir@71914.4]
  assign QueueCompatibility_1_reset = reset; // @[:freechips.rocketchip.system.DefaultRV32Config.fir@71915.4]
  assign QueueCompatibility_1_io_enq_valid = _T_77 & _T_37[1]; // @[UserYanker.scala 63:21:freechips.rocketchip.system.DefaultRV32Config.fir@72127.4]
  assign QueueCompatibility_1_io_enq_bits_tl_state_size = auto_in_ar_bits_echo_tl_state_size; // @[BundleMap.scala 248:19:freechips.rocketchip.system.DefaultRV32Config.fir@72129.4]
  assign QueueCompatibility_1_io_enq_bits_tl_state_source = auto_in_ar_bits_echo_tl_state_source; // @[BundleMap.scala 248:19:freechips.rocketchip.system.DefaultRV32Config.fir@72128.4]
  assign QueueCompatibility_1_io_deq_ready = _T_80 & auto_out_r_bits_last; // @[UserYanker.scala 62:21:freechips.rocketchip.system.DefaultRV32Config.fir@72124.4]
  assign QueueCompatibility_2_clock = clock; // @[:freechips.rocketchip.system.DefaultRV32Config.fir@71918.4]
  assign QueueCompatibility_2_reset = reset; // @[:freechips.rocketchip.system.DefaultRV32Config.fir@71919.4]
  assign QueueCompatibility_2_io_enq_valid = _T_77 & _T_37[2]; // @[UserYanker.scala 63:21:freechips.rocketchip.system.DefaultRV32Config.fir@72136.4]
  assign QueueCompatibility_2_io_enq_bits_tl_state_size = auto_in_ar_bits_echo_tl_state_size; // @[BundleMap.scala 248:19:freechips.rocketchip.system.DefaultRV32Config.fir@72138.4]
  assign QueueCompatibility_2_io_enq_bits_tl_state_source = auto_in_ar_bits_echo_tl_state_source; // @[BundleMap.scala 248:19:freechips.rocketchip.system.DefaultRV32Config.fir@72137.4]
  assign QueueCompatibility_2_io_deq_ready = _T_85 & auto_out_r_bits_last; // @[UserYanker.scala 62:21:freechips.rocketchip.system.DefaultRV32Config.fir@72133.4]
  assign QueueCompatibility_3_clock = clock; // @[:freechips.rocketchip.system.DefaultRV32Config.fir@71922.4]
  assign QueueCompatibility_3_reset = reset; // @[:freechips.rocketchip.system.DefaultRV32Config.fir@71923.4]
  assign QueueCompatibility_3_io_enq_valid = _T_77 & _T_37[3]; // @[UserYanker.scala 63:21:freechips.rocketchip.system.DefaultRV32Config.fir@72145.4]
  assign QueueCompatibility_3_io_enq_bits_tl_state_size = auto_in_ar_bits_echo_tl_state_size; // @[BundleMap.scala 248:19:freechips.rocketchip.system.DefaultRV32Config.fir@72147.4]
  assign QueueCompatibility_3_io_enq_bits_tl_state_source = auto_in_ar_bits_echo_tl_state_source; // @[BundleMap.scala 248:19:freechips.rocketchip.system.DefaultRV32Config.fir@72146.4]
  assign QueueCompatibility_3_io_deq_ready = _T_90 & auto_out_r_bits_last; // @[UserYanker.scala 62:21:freechips.rocketchip.system.DefaultRV32Config.fir@72142.4]
  assign QueueCompatibility_4_clock = clock; // @[:freechips.rocketchip.system.DefaultRV32Config.fir@71950.4]
  assign QueueCompatibility_4_reset = reset; // @[:freechips.rocketchip.system.DefaultRV32Config.fir@71951.4]
  assign QueueCompatibility_4_io_enq_valid = _T_204 & _T_165[0]; // @[UserYanker.scala 84:21:freechips.rocketchip.system.DefaultRV32Config.fir@72383.4]
  assign QueueCompatibility_4_io_enq_bits_tl_state_size = auto_in_aw_bits_echo_tl_state_size; // @[BundleMap.scala 248:19:freechips.rocketchip.system.DefaultRV32Config.fir@72385.4]
  assign QueueCompatibility_4_io_enq_bits_tl_state_source = auto_in_aw_bits_echo_tl_state_source; // @[BundleMap.scala 248:19:freechips.rocketchip.system.DefaultRV32Config.fir@72384.4]
  assign QueueCompatibility_4_io_deq_ready = _T_202 & _T_184[0]; // @[UserYanker.scala 83:21:freechips.rocketchip.system.DefaultRV32Config.fir@72380.4]
  assign QueueCompatibility_5_clock = clock; // @[:freechips.rocketchip.system.DefaultRV32Config.fir@71954.4]
  assign QueueCompatibility_5_reset = reset; // @[:freechips.rocketchip.system.DefaultRV32Config.fir@71955.4]
  assign QueueCompatibility_5_io_enq_valid = _T_204 & _T_165[1]; // @[UserYanker.scala 84:21:freechips.rocketchip.system.DefaultRV32Config.fir@72391.4]
  assign QueueCompatibility_5_io_enq_bits_tl_state_size = auto_in_aw_bits_echo_tl_state_size; // @[BundleMap.scala 248:19:freechips.rocketchip.system.DefaultRV32Config.fir@72393.4]
  assign QueueCompatibility_5_io_enq_bits_tl_state_source = auto_in_aw_bits_echo_tl_state_source; // @[BundleMap.scala 248:19:freechips.rocketchip.system.DefaultRV32Config.fir@72392.4]
  assign QueueCompatibility_5_io_deq_ready = _T_202 & _T_184[1]; // @[UserYanker.scala 83:21:freechips.rocketchip.system.DefaultRV32Config.fir@72388.4]
  assign QueueCompatibility_6_clock = clock; // @[:freechips.rocketchip.system.DefaultRV32Config.fir@71958.4]
  assign QueueCompatibility_6_reset = reset; // @[:freechips.rocketchip.system.DefaultRV32Config.fir@71959.4]
  assign QueueCompatibility_6_io_enq_valid = _T_204 & _T_165[2]; // @[UserYanker.scala 84:21:freechips.rocketchip.system.DefaultRV32Config.fir@72399.4]
  assign QueueCompatibility_6_io_enq_bits_tl_state_size = auto_in_aw_bits_echo_tl_state_size; // @[BundleMap.scala 248:19:freechips.rocketchip.system.DefaultRV32Config.fir@72401.4]
  assign QueueCompatibility_6_io_enq_bits_tl_state_source = auto_in_aw_bits_echo_tl_state_source; // @[BundleMap.scala 248:19:freechips.rocketchip.system.DefaultRV32Config.fir@72400.4]
  assign QueueCompatibility_6_io_deq_ready = _T_202 & _T_184[2]; // @[UserYanker.scala 83:21:freechips.rocketchip.system.DefaultRV32Config.fir@72396.4]
  assign QueueCompatibility_7_clock = clock; // @[:freechips.rocketchip.system.DefaultRV32Config.fir@71962.4]
  assign QueueCompatibility_7_reset = reset; // @[:freechips.rocketchip.system.DefaultRV32Config.fir@71963.4]
  assign QueueCompatibility_7_io_enq_valid = _T_204 & _T_165[3]; // @[UserYanker.scala 84:21:freechips.rocketchip.system.DefaultRV32Config.fir@72407.4]
  assign QueueCompatibility_7_io_enq_bits_tl_state_size = auto_in_aw_bits_echo_tl_state_size; // @[BundleMap.scala 248:19:freechips.rocketchip.system.DefaultRV32Config.fir@72409.4]
  assign QueueCompatibility_7_io_enq_bits_tl_state_source = auto_in_aw_bits_echo_tl_state_source; // @[BundleMap.scala 248:19:freechips.rocketchip.system.DefaultRV32Config.fir@72408.4]
  assign QueueCompatibility_7_io_deq_ready = _T_202 & _T_184[3]; // @[UserYanker.scala 83:21:freechips.rocketchip.system.DefaultRV32Config.fir@72404.4]
  always @(posedge clock) begin
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_35) begin
          $fwrite(32'h80000002,"Assertion failed\n    at UserYanker.scala:55 assert (!out.r.valid || r_valid) // Q must be ready faster than the response\n"); // @[UserYanker.scala 55:14:freechips.rocketchip.system.DefaultRV32Config.fir@72061.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_35) begin
          $fatal; // @[UserYanker.scala 55:14:freechips.rocketchip.system.DefaultRV32Config.fir@72062.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_163) begin
          $fwrite(32'h80000002,"Assertion failed\n    at UserYanker.scala:76 assert (!out.b.valid || b_valid) // Q must be ready faster than the response\n"); // @[UserYanker.scala 76:14:freechips.rocketchip.system.DefaultRV32Config.fir@72329.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_163) begin
          $fatal; // @[UserYanker.scala 76:14:freechips.rocketchip.system.DefaultRV32Config.fir@72330.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
  end
endmodule
