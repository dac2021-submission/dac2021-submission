module BroadcastFilter( // @[:freechips.rocketchip.system.DefaultRV32Config.fir@78834.2]
  output        io_request_ready, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@78837.4]
  input         io_request_valid, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@78837.4]
  input  [1:0]  io_request_bits_mshr, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@78837.4]
  input  [25:0] io_request_bits_address, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@78837.4]
  input         io_request_bits_allocOH, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@78837.4]
  input         io_request_bits_needT, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@78837.4]
  input         io_response_ready, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@78837.4]
  output        io_response_valid, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@78837.4]
  output [1:0]  io_response_bits_mshr, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@78837.4]
  output [25:0] io_response_bits_address, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@78837.4]
  output        io_response_bits_allocOH, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@78837.4]
  output        io_response_bits_needT // @[:freechips.rocketchip.system.DefaultRV32Config.fir@78837.4]
);
  assign io_request_ready = io_response_ready; // @[Broadcast.scala 339:20:freechips.rocketchip.system.DefaultRV32Config.fir@78843.4]
  assign io_response_valid = io_request_valid; // @[Broadcast.scala 340:21:freechips.rocketchip.system.DefaultRV32Config.fir@78844.4]
  assign io_response_bits_mshr = io_request_bits_mshr; // @[Broadcast.scala 342:28:freechips.rocketchip.system.DefaultRV32Config.fir@78845.4]
  assign io_response_bits_address = io_request_bits_address; // @[Broadcast.scala 343:28:freechips.rocketchip.system.DefaultRV32Config.fir@78846.4]
  assign io_response_bits_allocOH = io_request_bits_allocOH; // @[Broadcast.scala 345:28:freechips.rocketchip.system.DefaultRV32Config.fir@78848.4]
  assign io_response_bits_needT = io_request_bits_needT; // @[Broadcast.scala 344:28:freechips.rocketchip.system.DefaultRV32Config.fir@78847.4]
endmodule
