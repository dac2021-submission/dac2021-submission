module IntSyncCrossingSource( // @[:freechips.rocketchip.system.DefaultRV32Config.fir@99766.2]
  input   auto_in_0, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@99769.4]
  output  auto_out_sync_0 // @[:freechips.rocketchip.system.DefaultRV32Config.fir@99769.4]
);
  assign auto_out_sync_0 = auto_in_0; // @[LazyModule.scala 305:12:freechips.rocketchip.system.DefaultRV32Config.fir@99778.4]
endmodule
