module TLB_1( // @[:freechips.rocketchip.system.DefaultRV32Config.fir@198349.2]
  input         clock, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@198350.4]
  input         reset, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@198351.4]
  output        io_req_ready, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@198352.4]
  input         io_req_valid, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@198352.4]
  input  [31:0] io_req_bits_vaddr, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@198352.4]
  output        io_resp_miss, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@198352.4]
  output [31:0] io_resp_paddr, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@198352.4]
  output        io_resp_pf_inst, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@198352.4]
  output        io_resp_ae_inst, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@198352.4]
  output        io_resp_cacheable, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@198352.4]
  input         io_sfence_valid, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@198352.4]
  input         io_sfence_bits_rs1, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@198352.4]
  input         io_sfence_bits_rs2, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@198352.4]
  input  [31:0] io_sfence_bits_addr, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@198352.4]
  input         io_ptw_req_ready, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@198352.4]
  output        io_ptw_req_valid, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@198352.4]
  output        io_ptw_req_bits_valid, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@198352.4]
  output [19:0] io_ptw_req_bits_bits_addr, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@198352.4]
  input         io_ptw_resp_valid, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@198352.4]
  input         io_ptw_resp_bits_ae, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@198352.4]
  input  [53:0] io_ptw_resp_bits_pte_ppn, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@198352.4]
  input         io_ptw_resp_bits_pte_d, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@198352.4]
  input         io_ptw_resp_bits_pte_a, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@198352.4]
  input         io_ptw_resp_bits_pte_g, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@198352.4]
  input         io_ptw_resp_bits_pte_u, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@198352.4]
  input         io_ptw_resp_bits_pte_x, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@198352.4]
  input         io_ptw_resp_bits_pte_w, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@198352.4]
  input         io_ptw_resp_bits_pte_r, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@198352.4]
  input         io_ptw_resp_bits_pte_v, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@198352.4]
  input         io_ptw_resp_bits_level, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@198352.4]
  input         io_ptw_resp_bits_homogeneous, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@198352.4]
  input         io_ptw_ptbr_mode, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@198352.4]
  input         io_ptw_status_debug, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@198352.4]
  input  [1:0]  io_ptw_status_prv, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@198352.4]
  input         io_ptw_pmp_0_cfg_l, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@198352.4]
  input  [1:0]  io_ptw_pmp_0_cfg_a, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@198352.4]
  input         io_ptw_pmp_0_cfg_x, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@198352.4]
  input         io_ptw_pmp_0_cfg_w, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@198352.4]
  input         io_ptw_pmp_0_cfg_r, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@198352.4]
  input  [29:0] io_ptw_pmp_0_addr, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@198352.4]
  input  [31:0] io_ptw_pmp_0_mask, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@198352.4]
  input         io_ptw_pmp_1_cfg_l, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@198352.4]
  input  [1:0]  io_ptw_pmp_1_cfg_a, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@198352.4]
  input         io_ptw_pmp_1_cfg_x, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@198352.4]
  input         io_ptw_pmp_1_cfg_w, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@198352.4]
  input         io_ptw_pmp_1_cfg_r, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@198352.4]
  input  [29:0] io_ptw_pmp_1_addr, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@198352.4]
  input  [31:0] io_ptw_pmp_1_mask, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@198352.4]
  input         io_ptw_pmp_2_cfg_l, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@198352.4]
  input  [1:0]  io_ptw_pmp_2_cfg_a, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@198352.4]
  input         io_ptw_pmp_2_cfg_x, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@198352.4]
  input         io_ptw_pmp_2_cfg_w, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@198352.4]
  input         io_ptw_pmp_2_cfg_r, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@198352.4]
  input  [29:0] io_ptw_pmp_2_addr, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@198352.4]
  input  [31:0] io_ptw_pmp_2_mask, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@198352.4]
  input         io_ptw_pmp_3_cfg_l, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@198352.4]
  input  [1:0]  io_ptw_pmp_3_cfg_a, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@198352.4]
  input         io_ptw_pmp_3_cfg_x, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@198352.4]
  input         io_ptw_pmp_3_cfg_w, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@198352.4]
  input         io_ptw_pmp_3_cfg_r, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@198352.4]
  input  [29:0] io_ptw_pmp_3_addr, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@198352.4]
  input  [31:0] io_ptw_pmp_3_mask, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@198352.4]
  input         io_ptw_pmp_4_cfg_l, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@198352.4]
  input  [1:0]  io_ptw_pmp_4_cfg_a, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@198352.4]
  input         io_ptw_pmp_4_cfg_x, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@198352.4]
  input         io_ptw_pmp_4_cfg_w, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@198352.4]
  input         io_ptw_pmp_4_cfg_r, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@198352.4]
  input  [29:0] io_ptw_pmp_4_addr, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@198352.4]
  input  [31:0] io_ptw_pmp_4_mask, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@198352.4]
  input         io_ptw_pmp_5_cfg_l, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@198352.4]
  input  [1:0]  io_ptw_pmp_5_cfg_a, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@198352.4]
  input         io_ptw_pmp_5_cfg_x, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@198352.4]
  input         io_ptw_pmp_5_cfg_w, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@198352.4]
  input         io_ptw_pmp_5_cfg_r, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@198352.4]
  input  [29:0] io_ptw_pmp_5_addr, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@198352.4]
  input  [31:0] io_ptw_pmp_5_mask, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@198352.4]
  input         io_ptw_pmp_6_cfg_l, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@198352.4]
  input  [1:0]  io_ptw_pmp_6_cfg_a, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@198352.4]
  input         io_ptw_pmp_6_cfg_x, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@198352.4]
  input         io_ptw_pmp_6_cfg_w, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@198352.4]
  input         io_ptw_pmp_6_cfg_r, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@198352.4]
  input  [29:0] io_ptw_pmp_6_addr, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@198352.4]
  input  [31:0] io_ptw_pmp_6_mask, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@198352.4]
  input         io_ptw_pmp_7_cfg_l, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@198352.4]
  input  [1:0]  io_ptw_pmp_7_cfg_a, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@198352.4]
  input         io_ptw_pmp_7_cfg_x, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@198352.4]
  input         io_ptw_pmp_7_cfg_w, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@198352.4]
  input         io_ptw_pmp_7_cfg_r, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@198352.4]
  input  [29:0] io_ptw_pmp_7_addr, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@198352.4]
  input  [31:0] io_ptw_pmp_7_mask, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@198352.4]
  input         io_kill // @[:freechips.rocketchip.system.DefaultRV32Config.fir@198352.4]
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [63:0] _RAND_1;
  reg [63:0] _RAND_2;
  reg [63:0] _RAND_3;
  reg [63:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [63:0] _RAND_10;
  reg [63:0] _RAND_11;
  reg [63:0] _RAND_12;
  reg [63:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [63:0] _RAND_19;
  reg [63:0] _RAND_20;
  reg [63:0] _RAND_21;
  reg [63:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [63:0] _RAND_28;
  reg [63:0] _RAND_29;
  reg [63:0] _RAND_30;
  reg [63:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [31:0] _RAND_34;
  reg [31:0] _RAND_35;
  reg [31:0] _RAND_36;
  reg [63:0] _RAND_37;
  reg [63:0] _RAND_38;
  reg [63:0] _RAND_39;
  reg [63:0] _RAND_40;
  reg [31:0] _RAND_41;
  reg [31:0] _RAND_42;
  reg [31:0] _RAND_43;
  reg [31:0] _RAND_44;
  reg [31:0] _RAND_45;
  reg [63:0] _RAND_46;
  reg [63:0] _RAND_47;
  reg [63:0] _RAND_48;
  reg [63:0] _RAND_49;
  reg [31:0] _RAND_50;
  reg [31:0] _RAND_51;
  reg [31:0] _RAND_52;
  reg [31:0] _RAND_53;
  reg [31:0] _RAND_54;
  reg [63:0] _RAND_55;
  reg [63:0] _RAND_56;
  reg [63:0] _RAND_57;
  reg [63:0] _RAND_58;
  reg [31:0] _RAND_59;
  reg [31:0] _RAND_60;
  reg [31:0] _RAND_61;
  reg [31:0] _RAND_62;
  reg [31:0] _RAND_63;
  reg [63:0] _RAND_64;
  reg [63:0] _RAND_65;
  reg [63:0] _RAND_66;
  reg [63:0] _RAND_67;
  reg [31:0] _RAND_68;
  reg [31:0] _RAND_69;
  reg [31:0] _RAND_70;
  reg [31:0] _RAND_71;
  reg [31:0] _RAND_72;
  reg [63:0] _RAND_73;
  reg [31:0] _RAND_74;
  reg [31:0] _RAND_75;
  reg [63:0] _RAND_76;
  reg [31:0] _RAND_77;
  reg [31:0] _RAND_78;
  reg [63:0] _RAND_79;
  reg [31:0] _RAND_80;
  reg [31:0] _RAND_81;
  reg [63:0] _RAND_82;
  reg [31:0] _RAND_83;
  reg [31:0] _RAND_84;
  reg [31:0] _RAND_85;
  reg [63:0] _RAND_86;
  reg [31:0] _RAND_87;
  reg [31:0] _RAND_88;
  reg [31:0] _RAND_89;
  reg [31:0] _RAND_90;
  reg [31:0] _RAND_91;
  reg [31:0] _RAND_92;
  reg [31:0] _RAND_93;
  reg [31:0] _RAND_94;
  reg [31:0] _RAND_95;
`endif // RANDOMIZE_REG_INIT
  wire [19:0] OptimizationBarrier_io_x_ppn; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@198417.4]
  wire  OptimizationBarrier_io_x_u; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@198417.4]
  wire  OptimizationBarrier_io_x_ae; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@198417.4]
  wire  OptimizationBarrier_io_x_sw; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@198417.4]
  wire  OptimizationBarrier_io_x_sx; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@198417.4]
  wire  OptimizationBarrier_io_x_sr; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@198417.4]
  wire  OptimizationBarrier_io_x_pw; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@198417.4]
  wire  OptimizationBarrier_io_x_px; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@198417.4]
  wire  OptimizationBarrier_io_x_pr; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@198417.4]
  wire  OptimizationBarrier_io_x_ppp; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@198417.4]
  wire  OptimizationBarrier_io_x_pal; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@198417.4]
  wire  OptimizationBarrier_io_x_paa; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@198417.4]
  wire  OptimizationBarrier_io_x_eff; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@198417.4]
  wire  OptimizationBarrier_io_x_c; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@198417.4]
  wire [19:0] OptimizationBarrier_io_y_ppn; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@198417.4]
  wire  OptimizationBarrier_io_y_u; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@198417.4]
  wire  OptimizationBarrier_io_y_ae; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@198417.4]
  wire  OptimizationBarrier_io_y_sw; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@198417.4]
  wire  OptimizationBarrier_io_y_sx; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@198417.4]
  wire  OptimizationBarrier_io_y_sr; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@198417.4]
  wire  OptimizationBarrier_io_y_pw; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@198417.4]
  wire  OptimizationBarrier_io_y_px; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@198417.4]
  wire  OptimizationBarrier_io_y_pr; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@198417.4]
  wire  OptimizationBarrier_io_y_ppp; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@198417.4]
  wire  OptimizationBarrier_io_y_pal; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@198417.4]
  wire  OptimizationBarrier_io_y_paa; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@198417.4]
  wire  OptimizationBarrier_io_y_eff; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@198417.4]
  wire  OptimizationBarrier_io_y_c; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@198417.4]
  wire [1:0] pmp_io_prv; // @[TLB.scala 190:19:freechips.rocketchip.system.DefaultRV32Config.fir@198438.4]
  wire  pmp_io_pmp_0_cfg_l; // @[TLB.scala 190:19:freechips.rocketchip.system.DefaultRV32Config.fir@198438.4]
  wire [1:0] pmp_io_pmp_0_cfg_a; // @[TLB.scala 190:19:freechips.rocketchip.system.DefaultRV32Config.fir@198438.4]
  wire  pmp_io_pmp_0_cfg_x; // @[TLB.scala 190:19:freechips.rocketchip.system.DefaultRV32Config.fir@198438.4]
  wire  pmp_io_pmp_0_cfg_w; // @[TLB.scala 190:19:freechips.rocketchip.system.DefaultRV32Config.fir@198438.4]
  wire  pmp_io_pmp_0_cfg_r; // @[TLB.scala 190:19:freechips.rocketchip.system.DefaultRV32Config.fir@198438.4]
  wire [29:0] pmp_io_pmp_0_addr; // @[TLB.scala 190:19:freechips.rocketchip.system.DefaultRV32Config.fir@198438.4]
  wire [31:0] pmp_io_pmp_0_mask; // @[TLB.scala 190:19:freechips.rocketchip.system.DefaultRV32Config.fir@198438.4]
  wire  pmp_io_pmp_1_cfg_l; // @[TLB.scala 190:19:freechips.rocketchip.system.DefaultRV32Config.fir@198438.4]
  wire [1:0] pmp_io_pmp_1_cfg_a; // @[TLB.scala 190:19:freechips.rocketchip.system.DefaultRV32Config.fir@198438.4]
  wire  pmp_io_pmp_1_cfg_x; // @[TLB.scala 190:19:freechips.rocketchip.system.DefaultRV32Config.fir@198438.4]
  wire  pmp_io_pmp_1_cfg_w; // @[TLB.scala 190:19:freechips.rocketchip.system.DefaultRV32Config.fir@198438.4]
  wire  pmp_io_pmp_1_cfg_r; // @[TLB.scala 190:19:freechips.rocketchip.system.DefaultRV32Config.fir@198438.4]
  wire [29:0] pmp_io_pmp_1_addr; // @[TLB.scala 190:19:freechips.rocketchip.system.DefaultRV32Config.fir@198438.4]
  wire [31:0] pmp_io_pmp_1_mask; // @[TLB.scala 190:19:freechips.rocketchip.system.DefaultRV32Config.fir@198438.4]
  wire  pmp_io_pmp_2_cfg_l; // @[TLB.scala 190:19:freechips.rocketchip.system.DefaultRV32Config.fir@198438.4]
  wire [1:0] pmp_io_pmp_2_cfg_a; // @[TLB.scala 190:19:freechips.rocketchip.system.DefaultRV32Config.fir@198438.4]
  wire  pmp_io_pmp_2_cfg_x; // @[TLB.scala 190:19:freechips.rocketchip.system.DefaultRV32Config.fir@198438.4]
  wire  pmp_io_pmp_2_cfg_w; // @[TLB.scala 190:19:freechips.rocketchip.system.DefaultRV32Config.fir@198438.4]
  wire  pmp_io_pmp_2_cfg_r; // @[TLB.scala 190:19:freechips.rocketchip.system.DefaultRV32Config.fir@198438.4]
  wire [29:0] pmp_io_pmp_2_addr; // @[TLB.scala 190:19:freechips.rocketchip.system.DefaultRV32Config.fir@198438.4]
  wire [31:0] pmp_io_pmp_2_mask; // @[TLB.scala 190:19:freechips.rocketchip.system.DefaultRV32Config.fir@198438.4]
  wire  pmp_io_pmp_3_cfg_l; // @[TLB.scala 190:19:freechips.rocketchip.system.DefaultRV32Config.fir@198438.4]
  wire [1:0] pmp_io_pmp_3_cfg_a; // @[TLB.scala 190:19:freechips.rocketchip.system.DefaultRV32Config.fir@198438.4]
  wire  pmp_io_pmp_3_cfg_x; // @[TLB.scala 190:19:freechips.rocketchip.system.DefaultRV32Config.fir@198438.4]
  wire  pmp_io_pmp_3_cfg_w; // @[TLB.scala 190:19:freechips.rocketchip.system.DefaultRV32Config.fir@198438.4]
  wire  pmp_io_pmp_3_cfg_r; // @[TLB.scala 190:19:freechips.rocketchip.system.DefaultRV32Config.fir@198438.4]
  wire [29:0] pmp_io_pmp_3_addr; // @[TLB.scala 190:19:freechips.rocketchip.system.DefaultRV32Config.fir@198438.4]
  wire [31:0] pmp_io_pmp_3_mask; // @[TLB.scala 190:19:freechips.rocketchip.system.DefaultRV32Config.fir@198438.4]
  wire  pmp_io_pmp_4_cfg_l; // @[TLB.scala 190:19:freechips.rocketchip.system.DefaultRV32Config.fir@198438.4]
  wire [1:0] pmp_io_pmp_4_cfg_a; // @[TLB.scala 190:19:freechips.rocketchip.system.DefaultRV32Config.fir@198438.4]
  wire  pmp_io_pmp_4_cfg_x; // @[TLB.scala 190:19:freechips.rocketchip.system.DefaultRV32Config.fir@198438.4]
  wire  pmp_io_pmp_4_cfg_w; // @[TLB.scala 190:19:freechips.rocketchip.system.DefaultRV32Config.fir@198438.4]
  wire  pmp_io_pmp_4_cfg_r; // @[TLB.scala 190:19:freechips.rocketchip.system.DefaultRV32Config.fir@198438.4]
  wire [29:0] pmp_io_pmp_4_addr; // @[TLB.scala 190:19:freechips.rocketchip.system.DefaultRV32Config.fir@198438.4]
  wire [31:0] pmp_io_pmp_4_mask; // @[TLB.scala 190:19:freechips.rocketchip.system.DefaultRV32Config.fir@198438.4]
  wire  pmp_io_pmp_5_cfg_l; // @[TLB.scala 190:19:freechips.rocketchip.system.DefaultRV32Config.fir@198438.4]
  wire [1:0] pmp_io_pmp_5_cfg_a; // @[TLB.scala 190:19:freechips.rocketchip.system.DefaultRV32Config.fir@198438.4]
  wire  pmp_io_pmp_5_cfg_x; // @[TLB.scala 190:19:freechips.rocketchip.system.DefaultRV32Config.fir@198438.4]
  wire  pmp_io_pmp_5_cfg_w; // @[TLB.scala 190:19:freechips.rocketchip.system.DefaultRV32Config.fir@198438.4]
  wire  pmp_io_pmp_5_cfg_r; // @[TLB.scala 190:19:freechips.rocketchip.system.DefaultRV32Config.fir@198438.4]
  wire [29:0] pmp_io_pmp_5_addr; // @[TLB.scala 190:19:freechips.rocketchip.system.DefaultRV32Config.fir@198438.4]
  wire [31:0] pmp_io_pmp_5_mask; // @[TLB.scala 190:19:freechips.rocketchip.system.DefaultRV32Config.fir@198438.4]
  wire  pmp_io_pmp_6_cfg_l; // @[TLB.scala 190:19:freechips.rocketchip.system.DefaultRV32Config.fir@198438.4]
  wire [1:0] pmp_io_pmp_6_cfg_a; // @[TLB.scala 190:19:freechips.rocketchip.system.DefaultRV32Config.fir@198438.4]
  wire  pmp_io_pmp_6_cfg_x; // @[TLB.scala 190:19:freechips.rocketchip.system.DefaultRV32Config.fir@198438.4]
  wire  pmp_io_pmp_6_cfg_w; // @[TLB.scala 190:19:freechips.rocketchip.system.DefaultRV32Config.fir@198438.4]
  wire  pmp_io_pmp_6_cfg_r; // @[TLB.scala 190:19:freechips.rocketchip.system.DefaultRV32Config.fir@198438.4]
  wire [29:0] pmp_io_pmp_6_addr; // @[TLB.scala 190:19:freechips.rocketchip.system.DefaultRV32Config.fir@198438.4]
  wire [31:0] pmp_io_pmp_6_mask; // @[TLB.scala 190:19:freechips.rocketchip.system.DefaultRV32Config.fir@198438.4]
  wire  pmp_io_pmp_7_cfg_l; // @[TLB.scala 190:19:freechips.rocketchip.system.DefaultRV32Config.fir@198438.4]
  wire [1:0] pmp_io_pmp_7_cfg_a; // @[TLB.scala 190:19:freechips.rocketchip.system.DefaultRV32Config.fir@198438.4]
  wire  pmp_io_pmp_7_cfg_x; // @[TLB.scala 190:19:freechips.rocketchip.system.DefaultRV32Config.fir@198438.4]
  wire  pmp_io_pmp_7_cfg_w; // @[TLB.scala 190:19:freechips.rocketchip.system.DefaultRV32Config.fir@198438.4]
  wire  pmp_io_pmp_7_cfg_r; // @[TLB.scala 190:19:freechips.rocketchip.system.DefaultRV32Config.fir@198438.4]
  wire [29:0] pmp_io_pmp_7_addr; // @[TLB.scala 190:19:freechips.rocketchip.system.DefaultRV32Config.fir@198438.4]
  wire [31:0] pmp_io_pmp_7_mask; // @[TLB.scala 190:19:freechips.rocketchip.system.DefaultRV32Config.fir@198438.4]
  wire [31:0] pmp_io_addr; // @[TLB.scala 190:19:freechips.rocketchip.system.DefaultRV32Config.fir@198438.4]
  wire  pmp_io_r; // @[TLB.scala 190:19:freechips.rocketchip.system.DefaultRV32Config.fir@198438.4]
  wire  pmp_io_w; // @[TLB.scala 190:19:freechips.rocketchip.system.DefaultRV32Config.fir@198438.4]
  wire  pmp_io_x; // @[TLB.scala 190:19:freechips.rocketchip.system.DefaultRV32Config.fir@198438.4]
  wire [19:0] OptimizationBarrier_1_io_x_ppn; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@199139.4]
  wire  OptimizationBarrier_1_io_x_u; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@199139.4]
  wire  OptimizationBarrier_1_io_x_ae; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@199139.4]
  wire  OptimizationBarrier_1_io_x_sw; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@199139.4]
  wire  OptimizationBarrier_1_io_x_sx; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@199139.4]
  wire  OptimizationBarrier_1_io_x_sr; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@199139.4]
  wire  OptimizationBarrier_1_io_x_pw; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@199139.4]
  wire  OptimizationBarrier_1_io_x_px; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@199139.4]
  wire  OptimizationBarrier_1_io_x_pr; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@199139.4]
  wire  OptimizationBarrier_1_io_x_ppp; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@199139.4]
  wire  OptimizationBarrier_1_io_x_pal; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@199139.4]
  wire  OptimizationBarrier_1_io_x_paa; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@199139.4]
  wire  OptimizationBarrier_1_io_x_eff; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@199139.4]
  wire  OptimizationBarrier_1_io_x_c; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@199139.4]
  wire [19:0] OptimizationBarrier_1_io_y_ppn; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@199139.4]
  wire  OptimizationBarrier_1_io_y_u; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@199139.4]
  wire  OptimizationBarrier_1_io_y_ae; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@199139.4]
  wire  OptimizationBarrier_1_io_y_sw; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@199139.4]
  wire  OptimizationBarrier_1_io_y_sx; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@199139.4]
  wire  OptimizationBarrier_1_io_y_sr; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@199139.4]
  wire  OptimizationBarrier_1_io_y_pw; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@199139.4]
  wire  OptimizationBarrier_1_io_y_px; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@199139.4]
  wire  OptimizationBarrier_1_io_y_pr; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@199139.4]
  wire  OptimizationBarrier_1_io_y_ppp; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@199139.4]
  wire  OptimizationBarrier_1_io_y_pal; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@199139.4]
  wire  OptimizationBarrier_1_io_y_paa; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@199139.4]
  wire  OptimizationBarrier_1_io_y_eff; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@199139.4]
  wire  OptimizationBarrier_1_io_y_c; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@199139.4]
  wire [19:0] OptimizationBarrier_2_io_x_ppn; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@199182.4]
  wire  OptimizationBarrier_2_io_x_u; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@199182.4]
  wire  OptimizationBarrier_2_io_x_ae; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@199182.4]
  wire  OptimizationBarrier_2_io_x_sw; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@199182.4]
  wire  OptimizationBarrier_2_io_x_sx; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@199182.4]
  wire  OptimizationBarrier_2_io_x_sr; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@199182.4]
  wire  OptimizationBarrier_2_io_x_pw; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@199182.4]
  wire  OptimizationBarrier_2_io_x_px; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@199182.4]
  wire  OptimizationBarrier_2_io_x_pr; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@199182.4]
  wire  OptimizationBarrier_2_io_x_ppp; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@199182.4]
  wire  OptimizationBarrier_2_io_x_pal; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@199182.4]
  wire  OptimizationBarrier_2_io_x_paa; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@199182.4]
  wire  OptimizationBarrier_2_io_x_eff; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@199182.4]
  wire  OptimizationBarrier_2_io_x_c; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@199182.4]
  wire [19:0] OptimizationBarrier_2_io_y_ppn; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@199182.4]
  wire  OptimizationBarrier_2_io_y_u; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@199182.4]
  wire  OptimizationBarrier_2_io_y_ae; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@199182.4]
  wire  OptimizationBarrier_2_io_y_sw; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@199182.4]
  wire  OptimizationBarrier_2_io_y_sx; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@199182.4]
  wire  OptimizationBarrier_2_io_y_sr; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@199182.4]
  wire  OptimizationBarrier_2_io_y_pw; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@199182.4]
  wire  OptimizationBarrier_2_io_y_px; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@199182.4]
  wire  OptimizationBarrier_2_io_y_pr; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@199182.4]
  wire  OptimizationBarrier_2_io_y_ppp; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@199182.4]
  wire  OptimizationBarrier_2_io_y_pal; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@199182.4]
  wire  OptimizationBarrier_2_io_y_paa; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@199182.4]
  wire  OptimizationBarrier_2_io_y_eff; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@199182.4]
  wire  OptimizationBarrier_2_io_y_c; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@199182.4]
  wire [19:0] OptimizationBarrier_3_io_x_ppn; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@199225.4]
  wire  OptimizationBarrier_3_io_x_u; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@199225.4]
  wire  OptimizationBarrier_3_io_x_ae; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@199225.4]
  wire  OptimizationBarrier_3_io_x_sw; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@199225.4]
  wire  OptimizationBarrier_3_io_x_sx; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@199225.4]
  wire  OptimizationBarrier_3_io_x_sr; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@199225.4]
  wire  OptimizationBarrier_3_io_x_pw; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@199225.4]
  wire  OptimizationBarrier_3_io_x_px; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@199225.4]
  wire  OptimizationBarrier_3_io_x_pr; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@199225.4]
  wire  OptimizationBarrier_3_io_x_ppp; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@199225.4]
  wire  OptimizationBarrier_3_io_x_pal; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@199225.4]
  wire  OptimizationBarrier_3_io_x_paa; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@199225.4]
  wire  OptimizationBarrier_3_io_x_eff; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@199225.4]
  wire  OptimizationBarrier_3_io_x_c; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@199225.4]
  wire [19:0] OptimizationBarrier_3_io_y_ppn; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@199225.4]
  wire  OptimizationBarrier_3_io_y_u; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@199225.4]
  wire  OptimizationBarrier_3_io_y_ae; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@199225.4]
  wire  OptimizationBarrier_3_io_y_sw; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@199225.4]
  wire  OptimizationBarrier_3_io_y_sx; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@199225.4]
  wire  OptimizationBarrier_3_io_y_sr; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@199225.4]
  wire  OptimizationBarrier_3_io_y_pw; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@199225.4]
  wire  OptimizationBarrier_3_io_y_px; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@199225.4]
  wire  OptimizationBarrier_3_io_y_pr; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@199225.4]
  wire  OptimizationBarrier_3_io_y_ppp; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@199225.4]
  wire  OptimizationBarrier_3_io_y_pal; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@199225.4]
  wire  OptimizationBarrier_3_io_y_paa; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@199225.4]
  wire  OptimizationBarrier_3_io_y_eff; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@199225.4]
  wire  OptimizationBarrier_3_io_y_c; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@199225.4]
  wire [19:0] OptimizationBarrier_4_io_x_ppn; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@199268.4]
  wire  OptimizationBarrier_4_io_x_u; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@199268.4]
  wire  OptimizationBarrier_4_io_x_ae; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@199268.4]
  wire  OptimizationBarrier_4_io_x_sw; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@199268.4]
  wire  OptimizationBarrier_4_io_x_sx; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@199268.4]
  wire  OptimizationBarrier_4_io_x_sr; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@199268.4]
  wire  OptimizationBarrier_4_io_x_pw; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@199268.4]
  wire  OptimizationBarrier_4_io_x_px; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@199268.4]
  wire  OptimizationBarrier_4_io_x_pr; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@199268.4]
  wire  OptimizationBarrier_4_io_x_ppp; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@199268.4]
  wire  OptimizationBarrier_4_io_x_pal; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@199268.4]
  wire  OptimizationBarrier_4_io_x_paa; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@199268.4]
  wire  OptimizationBarrier_4_io_x_eff; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@199268.4]
  wire  OptimizationBarrier_4_io_x_c; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@199268.4]
  wire [19:0] OptimizationBarrier_4_io_y_ppn; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@199268.4]
  wire  OptimizationBarrier_4_io_y_u; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@199268.4]
  wire  OptimizationBarrier_4_io_y_ae; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@199268.4]
  wire  OptimizationBarrier_4_io_y_sw; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@199268.4]
  wire  OptimizationBarrier_4_io_y_sx; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@199268.4]
  wire  OptimizationBarrier_4_io_y_sr; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@199268.4]
  wire  OptimizationBarrier_4_io_y_pw; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@199268.4]
  wire  OptimizationBarrier_4_io_y_px; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@199268.4]
  wire  OptimizationBarrier_4_io_y_pr; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@199268.4]
  wire  OptimizationBarrier_4_io_y_ppp; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@199268.4]
  wire  OptimizationBarrier_4_io_y_pal; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@199268.4]
  wire  OptimizationBarrier_4_io_y_paa; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@199268.4]
  wire  OptimizationBarrier_4_io_y_eff; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@199268.4]
  wire  OptimizationBarrier_4_io_y_c; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@199268.4]
  wire [19:0] OptimizationBarrier_5_io_x_ppn; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@199311.4]
  wire  OptimizationBarrier_5_io_x_u; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@199311.4]
  wire  OptimizationBarrier_5_io_x_ae; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@199311.4]
  wire  OptimizationBarrier_5_io_x_sw; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@199311.4]
  wire  OptimizationBarrier_5_io_x_sx; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@199311.4]
  wire  OptimizationBarrier_5_io_x_sr; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@199311.4]
  wire  OptimizationBarrier_5_io_x_pw; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@199311.4]
  wire  OptimizationBarrier_5_io_x_px; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@199311.4]
  wire  OptimizationBarrier_5_io_x_pr; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@199311.4]
  wire  OptimizationBarrier_5_io_x_ppp; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@199311.4]
  wire  OptimizationBarrier_5_io_x_pal; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@199311.4]
  wire  OptimizationBarrier_5_io_x_paa; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@199311.4]
  wire  OptimizationBarrier_5_io_x_eff; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@199311.4]
  wire  OptimizationBarrier_5_io_x_c; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@199311.4]
  wire [19:0] OptimizationBarrier_5_io_y_ppn; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@199311.4]
  wire  OptimizationBarrier_5_io_y_u; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@199311.4]
  wire  OptimizationBarrier_5_io_y_ae; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@199311.4]
  wire  OptimizationBarrier_5_io_y_sw; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@199311.4]
  wire  OptimizationBarrier_5_io_y_sx; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@199311.4]
  wire  OptimizationBarrier_5_io_y_sr; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@199311.4]
  wire  OptimizationBarrier_5_io_y_pw; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@199311.4]
  wire  OptimizationBarrier_5_io_y_px; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@199311.4]
  wire  OptimizationBarrier_5_io_y_pr; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@199311.4]
  wire  OptimizationBarrier_5_io_y_ppp; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@199311.4]
  wire  OptimizationBarrier_5_io_y_pal; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@199311.4]
  wire  OptimizationBarrier_5_io_y_paa; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@199311.4]
  wire  OptimizationBarrier_5_io_y_eff; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@199311.4]
  wire  OptimizationBarrier_5_io_y_c; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@199311.4]
  wire [19:0] OptimizationBarrier_6_io_x_ppn; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@199354.4]
  wire  OptimizationBarrier_6_io_x_u; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@199354.4]
  wire  OptimizationBarrier_6_io_x_ae; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@199354.4]
  wire  OptimizationBarrier_6_io_x_sw; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@199354.4]
  wire  OptimizationBarrier_6_io_x_sx; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@199354.4]
  wire  OptimizationBarrier_6_io_x_sr; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@199354.4]
  wire  OptimizationBarrier_6_io_x_pw; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@199354.4]
  wire  OptimizationBarrier_6_io_x_px; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@199354.4]
  wire  OptimizationBarrier_6_io_x_pr; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@199354.4]
  wire  OptimizationBarrier_6_io_x_ppp; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@199354.4]
  wire  OptimizationBarrier_6_io_x_pal; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@199354.4]
  wire  OptimizationBarrier_6_io_x_paa; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@199354.4]
  wire  OptimizationBarrier_6_io_x_eff; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@199354.4]
  wire  OptimizationBarrier_6_io_x_c; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@199354.4]
  wire [19:0] OptimizationBarrier_6_io_y_ppn; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@199354.4]
  wire  OptimizationBarrier_6_io_y_u; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@199354.4]
  wire  OptimizationBarrier_6_io_y_ae; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@199354.4]
  wire  OptimizationBarrier_6_io_y_sw; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@199354.4]
  wire  OptimizationBarrier_6_io_y_sx; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@199354.4]
  wire  OptimizationBarrier_6_io_y_sr; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@199354.4]
  wire  OptimizationBarrier_6_io_y_pw; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@199354.4]
  wire  OptimizationBarrier_6_io_y_px; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@199354.4]
  wire  OptimizationBarrier_6_io_y_pr; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@199354.4]
  wire  OptimizationBarrier_6_io_y_ppp; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@199354.4]
  wire  OptimizationBarrier_6_io_y_pal; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@199354.4]
  wire  OptimizationBarrier_6_io_y_paa; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@199354.4]
  wire  OptimizationBarrier_6_io_y_eff; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@199354.4]
  wire  OptimizationBarrier_6_io_y_c; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@199354.4]
  wire [19:0] OptimizationBarrier_7_io_x_ppn; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@199397.4]
  wire  OptimizationBarrier_7_io_x_u; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@199397.4]
  wire  OptimizationBarrier_7_io_x_ae; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@199397.4]
  wire  OptimizationBarrier_7_io_x_sw; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@199397.4]
  wire  OptimizationBarrier_7_io_x_sx; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@199397.4]
  wire  OptimizationBarrier_7_io_x_sr; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@199397.4]
  wire  OptimizationBarrier_7_io_x_pw; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@199397.4]
  wire  OptimizationBarrier_7_io_x_px; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@199397.4]
  wire  OptimizationBarrier_7_io_x_pr; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@199397.4]
  wire  OptimizationBarrier_7_io_x_ppp; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@199397.4]
  wire  OptimizationBarrier_7_io_x_pal; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@199397.4]
  wire  OptimizationBarrier_7_io_x_paa; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@199397.4]
  wire  OptimizationBarrier_7_io_x_eff; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@199397.4]
  wire  OptimizationBarrier_7_io_x_c; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@199397.4]
  wire [19:0] OptimizationBarrier_7_io_y_ppn; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@199397.4]
  wire  OptimizationBarrier_7_io_y_u; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@199397.4]
  wire  OptimizationBarrier_7_io_y_ae; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@199397.4]
  wire  OptimizationBarrier_7_io_y_sw; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@199397.4]
  wire  OptimizationBarrier_7_io_y_sx; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@199397.4]
  wire  OptimizationBarrier_7_io_y_sr; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@199397.4]
  wire  OptimizationBarrier_7_io_y_pw; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@199397.4]
  wire  OptimizationBarrier_7_io_y_px; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@199397.4]
  wire  OptimizationBarrier_7_io_y_pr; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@199397.4]
  wire  OptimizationBarrier_7_io_y_ppp; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@199397.4]
  wire  OptimizationBarrier_7_io_y_pal; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@199397.4]
  wire  OptimizationBarrier_7_io_y_paa; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@199397.4]
  wire  OptimizationBarrier_7_io_y_eff; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@199397.4]
  wire  OptimizationBarrier_7_io_y_c; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@199397.4]
  wire [19:0] OptimizationBarrier_8_io_x_ppn; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@199440.4]
  wire  OptimizationBarrier_8_io_x_u; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@199440.4]
  wire  OptimizationBarrier_8_io_x_ae; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@199440.4]
  wire  OptimizationBarrier_8_io_x_sw; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@199440.4]
  wire  OptimizationBarrier_8_io_x_sx; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@199440.4]
  wire  OptimizationBarrier_8_io_x_sr; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@199440.4]
  wire  OptimizationBarrier_8_io_x_pw; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@199440.4]
  wire  OptimizationBarrier_8_io_x_px; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@199440.4]
  wire  OptimizationBarrier_8_io_x_pr; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@199440.4]
  wire  OptimizationBarrier_8_io_x_ppp; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@199440.4]
  wire  OptimizationBarrier_8_io_x_pal; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@199440.4]
  wire  OptimizationBarrier_8_io_x_paa; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@199440.4]
  wire  OptimizationBarrier_8_io_x_eff; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@199440.4]
  wire  OptimizationBarrier_8_io_x_c; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@199440.4]
  wire [19:0] OptimizationBarrier_8_io_y_ppn; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@199440.4]
  wire  OptimizationBarrier_8_io_y_u; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@199440.4]
  wire  OptimizationBarrier_8_io_y_ae; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@199440.4]
  wire  OptimizationBarrier_8_io_y_sw; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@199440.4]
  wire  OptimizationBarrier_8_io_y_sx; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@199440.4]
  wire  OptimizationBarrier_8_io_y_sr; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@199440.4]
  wire  OptimizationBarrier_8_io_y_pw; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@199440.4]
  wire  OptimizationBarrier_8_io_y_px; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@199440.4]
  wire  OptimizationBarrier_8_io_y_pr; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@199440.4]
  wire  OptimizationBarrier_8_io_y_ppp; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@199440.4]
  wire  OptimizationBarrier_8_io_y_pal; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@199440.4]
  wire  OptimizationBarrier_8_io_y_paa; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@199440.4]
  wire  OptimizationBarrier_8_io_y_eff; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@199440.4]
  wire  OptimizationBarrier_8_io_y_c; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@199440.4]
  wire [19:0] OptimizationBarrier_9_io_x_ppn; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@199482.4]
  wire  OptimizationBarrier_9_io_x_u; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@199482.4]
  wire  OptimizationBarrier_9_io_x_ae; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@199482.4]
  wire  OptimizationBarrier_9_io_x_sw; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@199482.4]
  wire  OptimizationBarrier_9_io_x_sx; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@199482.4]
  wire  OptimizationBarrier_9_io_x_sr; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@199482.4]
  wire  OptimizationBarrier_9_io_x_pw; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@199482.4]
  wire  OptimizationBarrier_9_io_x_px; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@199482.4]
  wire  OptimizationBarrier_9_io_x_pr; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@199482.4]
  wire  OptimizationBarrier_9_io_x_ppp; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@199482.4]
  wire  OptimizationBarrier_9_io_x_pal; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@199482.4]
  wire  OptimizationBarrier_9_io_x_paa; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@199482.4]
  wire  OptimizationBarrier_9_io_x_eff; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@199482.4]
  wire  OptimizationBarrier_9_io_x_c; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@199482.4]
  wire [19:0] OptimizationBarrier_9_io_y_ppn; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@199482.4]
  wire  OptimizationBarrier_9_io_y_u; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@199482.4]
  wire  OptimizationBarrier_9_io_y_ae; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@199482.4]
  wire  OptimizationBarrier_9_io_y_sw; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@199482.4]
  wire  OptimizationBarrier_9_io_y_sx; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@199482.4]
  wire  OptimizationBarrier_9_io_y_sr; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@199482.4]
  wire  OptimizationBarrier_9_io_y_pw; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@199482.4]
  wire  OptimizationBarrier_9_io_y_px; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@199482.4]
  wire  OptimizationBarrier_9_io_y_pr; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@199482.4]
  wire  OptimizationBarrier_9_io_y_ppp; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@199482.4]
  wire  OptimizationBarrier_9_io_y_pal; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@199482.4]
  wire  OptimizationBarrier_9_io_y_paa; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@199482.4]
  wire  OptimizationBarrier_9_io_y_eff; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@199482.4]
  wire  OptimizationBarrier_9_io_y_c; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@199482.4]
  wire [19:0] OptimizationBarrier_10_io_x_ppn; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@199531.4]
  wire  OptimizationBarrier_10_io_x_u; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@199531.4]
  wire  OptimizationBarrier_10_io_x_ae; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@199531.4]
  wire  OptimizationBarrier_10_io_x_sw; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@199531.4]
  wire  OptimizationBarrier_10_io_x_sx; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@199531.4]
  wire  OptimizationBarrier_10_io_x_sr; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@199531.4]
  wire  OptimizationBarrier_10_io_x_pw; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@199531.4]
  wire  OptimizationBarrier_10_io_x_px; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@199531.4]
  wire  OptimizationBarrier_10_io_x_pr; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@199531.4]
  wire  OptimizationBarrier_10_io_x_ppp; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@199531.4]
  wire  OptimizationBarrier_10_io_x_pal; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@199531.4]
  wire  OptimizationBarrier_10_io_x_paa; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@199531.4]
  wire  OptimizationBarrier_10_io_x_eff; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@199531.4]
  wire  OptimizationBarrier_10_io_x_c; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@199531.4]
  wire [19:0] OptimizationBarrier_10_io_y_ppn; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@199531.4]
  wire  OptimizationBarrier_10_io_y_u; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@199531.4]
  wire  OptimizationBarrier_10_io_y_ae; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@199531.4]
  wire  OptimizationBarrier_10_io_y_sw; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@199531.4]
  wire  OptimizationBarrier_10_io_y_sx; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@199531.4]
  wire  OptimizationBarrier_10_io_y_sr; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@199531.4]
  wire  OptimizationBarrier_10_io_y_pw; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@199531.4]
  wire  OptimizationBarrier_10_io_y_px; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@199531.4]
  wire  OptimizationBarrier_10_io_y_pr; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@199531.4]
  wire  OptimizationBarrier_10_io_y_ppp; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@199531.4]
  wire  OptimizationBarrier_10_io_y_pal; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@199531.4]
  wire  OptimizationBarrier_10_io_y_paa; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@199531.4]
  wire  OptimizationBarrier_10_io_y_eff; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@199531.4]
  wire  OptimizationBarrier_10_io_y_c; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@199531.4]
  wire [19:0] OptimizationBarrier_11_io_x_ppn; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@199580.4]
  wire  OptimizationBarrier_11_io_x_u; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@199580.4]
  wire  OptimizationBarrier_11_io_x_ae; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@199580.4]
  wire  OptimizationBarrier_11_io_x_sw; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@199580.4]
  wire  OptimizationBarrier_11_io_x_sx; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@199580.4]
  wire  OptimizationBarrier_11_io_x_sr; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@199580.4]
  wire  OptimizationBarrier_11_io_x_pw; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@199580.4]
  wire  OptimizationBarrier_11_io_x_px; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@199580.4]
  wire  OptimizationBarrier_11_io_x_pr; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@199580.4]
  wire  OptimizationBarrier_11_io_x_ppp; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@199580.4]
  wire  OptimizationBarrier_11_io_x_pal; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@199580.4]
  wire  OptimizationBarrier_11_io_x_paa; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@199580.4]
  wire  OptimizationBarrier_11_io_x_eff; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@199580.4]
  wire  OptimizationBarrier_11_io_x_c; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@199580.4]
  wire [19:0] OptimizationBarrier_11_io_y_ppn; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@199580.4]
  wire  OptimizationBarrier_11_io_y_u; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@199580.4]
  wire  OptimizationBarrier_11_io_y_ae; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@199580.4]
  wire  OptimizationBarrier_11_io_y_sw; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@199580.4]
  wire  OptimizationBarrier_11_io_y_sx; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@199580.4]
  wire  OptimizationBarrier_11_io_y_sr; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@199580.4]
  wire  OptimizationBarrier_11_io_y_pw; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@199580.4]
  wire  OptimizationBarrier_11_io_y_px; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@199580.4]
  wire  OptimizationBarrier_11_io_y_pr; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@199580.4]
  wire  OptimizationBarrier_11_io_y_ppp; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@199580.4]
  wire  OptimizationBarrier_11_io_y_pal; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@199580.4]
  wire  OptimizationBarrier_11_io_y_paa; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@199580.4]
  wire  OptimizationBarrier_11_io_y_eff; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@199580.4]
  wire  OptimizationBarrier_11_io_y_c; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@199580.4]
  wire [19:0] OptimizationBarrier_12_io_x_ppn; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@199629.4]
  wire  OptimizationBarrier_12_io_x_u; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@199629.4]
  wire  OptimizationBarrier_12_io_x_ae; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@199629.4]
  wire  OptimizationBarrier_12_io_x_sw; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@199629.4]
  wire  OptimizationBarrier_12_io_x_sx; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@199629.4]
  wire  OptimizationBarrier_12_io_x_sr; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@199629.4]
  wire  OptimizationBarrier_12_io_x_pw; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@199629.4]
  wire  OptimizationBarrier_12_io_x_px; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@199629.4]
  wire  OptimizationBarrier_12_io_x_pr; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@199629.4]
  wire  OptimizationBarrier_12_io_x_ppp; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@199629.4]
  wire  OptimizationBarrier_12_io_x_pal; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@199629.4]
  wire  OptimizationBarrier_12_io_x_paa; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@199629.4]
  wire  OptimizationBarrier_12_io_x_eff; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@199629.4]
  wire  OptimizationBarrier_12_io_x_c; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@199629.4]
  wire [19:0] OptimizationBarrier_12_io_y_ppn; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@199629.4]
  wire  OptimizationBarrier_12_io_y_u; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@199629.4]
  wire  OptimizationBarrier_12_io_y_ae; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@199629.4]
  wire  OptimizationBarrier_12_io_y_sw; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@199629.4]
  wire  OptimizationBarrier_12_io_y_sx; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@199629.4]
  wire  OptimizationBarrier_12_io_y_sr; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@199629.4]
  wire  OptimizationBarrier_12_io_y_pw; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@199629.4]
  wire  OptimizationBarrier_12_io_y_px; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@199629.4]
  wire  OptimizationBarrier_12_io_y_pr; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@199629.4]
  wire  OptimizationBarrier_12_io_y_ppp; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@199629.4]
  wire  OptimizationBarrier_12_io_y_pal; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@199629.4]
  wire  OptimizationBarrier_12_io_y_paa; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@199629.4]
  wire  OptimizationBarrier_12_io_y_eff; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@199629.4]
  wire  OptimizationBarrier_12_io_y_c; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@199629.4]
  wire [19:0] OptimizationBarrier_13_io_x_ppn; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@199678.4]
  wire  OptimizationBarrier_13_io_x_u; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@199678.4]
  wire  OptimizationBarrier_13_io_x_ae; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@199678.4]
  wire  OptimizationBarrier_13_io_x_sw; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@199678.4]
  wire  OptimizationBarrier_13_io_x_sx; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@199678.4]
  wire  OptimizationBarrier_13_io_x_sr; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@199678.4]
  wire  OptimizationBarrier_13_io_x_pw; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@199678.4]
  wire  OptimizationBarrier_13_io_x_px; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@199678.4]
  wire  OptimizationBarrier_13_io_x_pr; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@199678.4]
  wire  OptimizationBarrier_13_io_x_ppp; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@199678.4]
  wire  OptimizationBarrier_13_io_x_pal; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@199678.4]
  wire  OptimizationBarrier_13_io_x_paa; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@199678.4]
  wire  OptimizationBarrier_13_io_x_eff; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@199678.4]
  wire  OptimizationBarrier_13_io_x_c; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@199678.4]
  wire [19:0] OptimizationBarrier_13_io_y_ppn; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@199678.4]
  wire  OptimizationBarrier_13_io_y_u; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@199678.4]
  wire  OptimizationBarrier_13_io_y_ae; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@199678.4]
  wire  OptimizationBarrier_13_io_y_sw; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@199678.4]
  wire  OptimizationBarrier_13_io_y_sx; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@199678.4]
  wire  OptimizationBarrier_13_io_y_sr; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@199678.4]
  wire  OptimizationBarrier_13_io_y_pw; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@199678.4]
  wire  OptimizationBarrier_13_io_y_px; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@199678.4]
  wire  OptimizationBarrier_13_io_y_pr; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@199678.4]
  wire  OptimizationBarrier_13_io_y_ppp; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@199678.4]
  wire  OptimizationBarrier_13_io_y_pal; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@199678.4]
  wire  OptimizationBarrier_13_io_y_paa; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@199678.4]
  wire  OptimizationBarrier_13_io_y_eff; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@199678.4]
  wire  OptimizationBarrier_13_io_y_c; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@199678.4]
  wire [19:0] OptimizationBarrier_14_io_x_ppn; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@200159.4]
  wire  OptimizationBarrier_14_io_x_u; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@200159.4]
  wire  OptimizationBarrier_14_io_x_ae; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@200159.4]
  wire  OptimizationBarrier_14_io_x_sw; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@200159.4]
  wire  OptimizationBarrier_14_io_x_sx; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@200159.4]
  wire  OptimizationBarrier_14_io_x_sr; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@200159.4]
  wire  OptimizationBarrier_14_io_x_pw; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@200159.4]
  wire  OptimizationBarrier_14_io_x_px; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@200159.4]
  wire  OptimizationBarrier_14_io_x_pr; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@200159.4]
  wire  OptimizationBarrier_14_io_x_ppp; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@200159.4]
  wire  OptimizationBarrier_14_io_x_pal; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@200159.4]
  wire  OptimizationBarrier_14_io_x_paa; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@200159.4]
  wire  OptimizationBarrier_14_io_x_eff; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@200159.4]
  wire  OptimizationBarrier_14_io_x_c; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@200159.4]
  wire [19:0] OptimizationBarrier_14_io_y_ppn; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@200159.4]
  wire  OptimizationBarrier_14_io_y_u; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@200159.4]
  wire  OptimizationBarrier_14_io_y_ae; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@200159.4]
  wire  OptimizationBarrier_14_io_y_sw; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@200159.4]
  wire  OptimizationBarrier_14_io_y_sx; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@200159.4]
  wire  OptimizationBarrier_14_io_y_sr; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@200159.4]
  wire  OptimizationBarrier_14_io_y_pw; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@200159.4]
  wire  OptimizationBarrier_14_io_y_px; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@200159.4]
  wire  OptimizationBarrier_14_io_y_pr; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@200159.4]
  wire  OptimizationBarrier_14_io_y_ppp; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@200159.4]
  wire  OptimizationBarrier_14_io_y_pal; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@200159.4]
  wire  OptimizationBarrier_14_io_y_paa; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@200159.4]
  wire  OptimizationBarrier_14_io_y_eff; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@200159.4]
  wire  OptimizationBarrier_14_io_y_c; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@200159.4]
  wire [19:0] OptimizationBarrier_15_io_x_ppn; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@200202.4]
  wire  OptimizationBarrier_15_io_x_u; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@200202.4]
  wire  OptimizationBarrier_15_io_x_ae; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@200202.4]
  wire  OptimizationBarrier_15_io_x_sw; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@200202.4]
  wire  OptimizationBarrier_15_io_x_sx; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@200202.4]
  wire  OptimizationBarrier_15_io_x_sr; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@200202.4]
  wire  OptimizationBarrier_15_io_x_pw; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@200202.4]
  wire  OptimizationBarrier_15_io_x_px; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@200202.4]
  wire  OptimizationBarrier_15_io_x_pr; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@200202.4]
  wire  OptimizationBarrier_15_io_x_ppp; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@200202.4]
  wire  OptimizationBarrier_15_io_x_pal; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@200202.4]
  wire  OptimizationBarrier_15_io_x_paa; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@200202.4]
  wire  OptimizationBarrier_15_io_x_eff; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@200202.4]
  wire  OptimizationBarrier_15_io_x_c; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@200202.4]
  wire [19:0] OptimizationBarrier_15_io_y_ppn; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@200202.4]
  wire  OptimizationBarrier_15_io_y_u; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@200202.4]
  wire  OptimizationBarrier_15_io_y_ae; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@200202.4]
  wire  OptimizationBarrier_15_io_y_sw; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@200202.4]
  wire  OptimizationBarrier_15_io_y_sx; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@200202.4]
  wire  OptimizationBarrier_15_io_y_sr; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@200202.4]
  wire  OptimizationBarrier_15_io_y_pw; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@200202.4]
  wire  OptimizationBarrier_15_io_y_px; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@200202.4]
  wire  OptimizationBarrier_15_io_y_pr; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@200202.4]
  wire  OptimizationBarrier_15_io_y_ppp; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@200202.4]
  wire  OptimizationBarrier_15_io_y_pal; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@200202.4]
  wire  OptimizationBarrier_15_io_y_paa; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@200202.4]
  wire  OptimizationBarrier_15_io_y_eff; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@200202.4]
  wire  OptimizationBarrier_15_io_y_c; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@200202.4]
  wire [19:0] OptimizationBarrier_16_io_x_ppn; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@200245.4]
  wire  OptimizationBarrier_16_io_x_u; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@200245.4]
  wire  OptimizationBarrier_16_io_x_ae; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@200245.4]
  wire  OptimizationBarrier_16_io_x_sw; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@200245.4]
  wire  OptimizationBarrier_16_io_x_sx; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@200245.4]
  wire  OptimizationBarrier_16_io_x_sr; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@200245.4]
  wire  OptimizationBarrier_16_io_x_pw; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@200245.4]
  wire  OptimizationBarrier_16_io_x_px; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@200245.4]
  wire  OptimizationBarrier_16_io_x_pr; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@200245.4]
  wire  OptimizationBarrier_16_io_x_ppp; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@200245.4]
  wire  OptimizationBarrier_16_io_x_pal; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@200245.4]
  wire  OptimizationBarrier_16_io_x_paa; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@200245.4]
  wire  OptimizationBarrier_16_io_x_eff; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@200245.4]
  wire  OptimizationBarrier_16_io_x_c; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@200245.4]
  wire [19:0] OptimizationBarrier_16_io_y_ppn; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@200245.4]
  wire  OptimizationBarrier_16_io_y_u; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@200245.4]
  wire  OptimizationBarrier_16_io_y_ae; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@200245.4]
  wire  OptimizationBarrier_16_io_y_sw; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@200245.4]
  wire  OptimizationBarrier_16_io_y_sx; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@200245.4]
  wire  OptimizationBarrier_16_io_y_sr; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@200245.4]
  wire  OptimizationBarrier_16_io_y_pw; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@200245.4]
  wire  OptimizationBarrier_16_io_y_px; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@200245.4]
  wire  OptimizationBarrier_16_io_y_pr; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@200245.4]
  wire  OptimizationBarrier_16_io_y_ppp; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@200245.4]
  wire  OptimizationBarrier_16_io_y_pal; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@200245.4]
  wire  OptimizationBarrier_16_io_y_paa; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@200245.4]
  wire  OptimizationBarrier_16_io_y_eff; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@200245.4]
  wire  OptimizationBarrier_16_io_y_c; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@200245.4]
  wire [19:0] OptimizationBarrier_17_io_x_ppn; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@200288.4]
  wire  OptimizationBarrier_17_io_x_u; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@200288.4]
  wire  OptimizationBarrier_17_io_x_ae; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@200288.4]
  wire  OptimizationBarrier_17_io_x_sw; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@200288.4]
  wire  OptimizationBarrier_17_io_x_sx; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@200288.4]
  wire  OptimizationBarrier_17_io_x_sr; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@200288.4]
  wire  OptimizationBarrier_17_io_x_pw; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@200288.4]
  wire  OptimizationBarrier_17_io_x_px; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@200288.4]
  wire  OptimizationBarrier_17_io_x_pr; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@200288.4]
  wire  OptimizationBarrier_17_io_x_ppp; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@200288.4]
  wire  OptimizationBarrier_17_io_x_pal; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@200288.4]
  wire  OptimizationBarrier_17_io_x_paa; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@200288.4]
  wire  OptimizationBarrier_17_io_x_eff; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@200288.4]
  wire  OptimizationBarrier_17_io_x_c; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@200288.4]
  wire [19:0] OptimizationBarrier_17_io_y_ppn; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@200288.4]
  wire  OptimizationBarrier_17_io_y_u; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@200288.4]
  wire  OptimizationBarrier_17_io_y_ae; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@200288.4]
  wire  OptimizationBarrier_17_io_y_sw; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@200288.4]
  wire  OptimizationBarrier_17_io_y_sx; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@200288.4]
  wire  OptimizationBarrier_17_io_y_sr; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@200288.4]
  wire  OptimizationBarrier_17_io_y_pw; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@200288.4]
  wire  OptimizationBarrier_17_io_y_px; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@200288.4]
  wire  OptimizationBarrier_17_io_y_pr; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@200288.4]
  wire  OptimizationBarrier_17_io_y_ppp; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@200288.4]
  wire  OptimizationBarrier_17_io_y_pal; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@200288.4]
  wire  OptimizationBarrier_17_io_y_paa; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@200288.4]
  wire  OptimizationBarrier_17_io_y_eff; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@200288.4]
  wire  OptimizationBarrier_17_io_y_c; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@200288.4]
  wire [19:0] OptimizationBarrier_18_io_x_ppn; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@200331.4]
  wire  OptimizationBarrier_18_io_x_u; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@200331.4]
  wire  OptimizationBarrier_18_io_x_ae; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@200331.4]
  wire  OptimizationBarrier_18_io_x_sw; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@200331.4]
  wire  OptimizationBarrier_18_io_x_sx; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@200331.4]
  wire  OptimizationBarrier_18_io_x_sr; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@200331.4]
  wire  OptimizationBarrier_18_io_x_pw; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@200331.4]
  wire  OptimizationBarrier_18_io_x_px; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@200331.4]
  wire  OptimizationBarrier_18_io_x_pr; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@200331.4]
  wire  OptimizationBarrier_18_io_x_ppp; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@200331.4]
  wire  OptimizationBarrier_18_io_x_pal; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@200331.4]
  wire  OptimizationBarrier_18_io_x_paa; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@200331.4]
  wire  OptimizationBarrier_18_io_x_eff; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@200331.4]
  wire  OptimizationBarrier_18_io_x_c; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@200331.4]
  wire [19:0] OptimizationBarrier_18_io_y_ppn; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@200331.4]
  wire  OptimizationBarrier_18_io_y_u; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@200331.4]
  wire  OptimizationBarrier_18_io_y_ae; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@200331.4]
  wire  OptimizationBarrier_18_io_y_sw; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@200331.4]
  wire  OptimizationBarrier_18_io_y_sx; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@200331.4]
  wire  OptimizationBarrier_18_io_y_sr; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@200331.4]
  wire  OptimizationBarrier_18_io_y_pw; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@200331.4]
  wire  OptimizationBarrier_18_io_y_px; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@200331.4]
  wire  OptimizationBarrier_18_io_y_pr; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@200331.4]
  wire  OptimizationBarrier_18_io_y_ppp; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@200331.4]
  wire  OptimizationBarrier_18_io_y_pal; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@200331.4]
  wire  OptimizationBarrier_18_io_y_paa; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@200331.4]
  wire  OptimizationBarrier_18_io_y_eff; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@200331.4]
  wire  OptimizationBarrier_18_io_y_c; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@200331.4]
  wire [19:0] OptimizationBarrier_19_io_x_ppn; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@200374.4]
  wire  OptimizationBarrier_19_io_x_u; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@200374.4]
  wire  OptimizationBarrier_19_io_x_ae; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@200374.4]
  wire  OptimizationBarrier_19_io_x_sw; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@200374.4]
  wire  OptimizationBarrier_19_io_x_sx; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@200374.4]
  wire  OptimizationBarrier_19_io_x_sr; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@200374.4]
  wire  OptimizationBarrier_19_io_x_pw; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@200374.4]
  wire  OptimizationBarrier_19_io_x_px; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@200374.4]
  wire  OptimizationBarrier_19_io_x_pr; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@200374.4]
  wire  OptimizationBarrier_19_io_x_ppp; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@200374.4]
  wire  OptimizationBarrier_19_io_x_pal; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@200374.4]
  wire  OptimizationBarrier_19_io_x_paa; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@200374.4]
  wire  OptimizationBarrier_19_io_x_eff; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@200374.4]
  wire  OptimizationBarrier_19_io_x_c; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@200374.4]
  wire [19:0] OptimizationBarrier_19_io_y_ppn; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@200374.4]
  wire  OptimizationBarrier_19_io_y_u; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@200374.4]
  wire  OptimizationBarrier_19_io_y_ae; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@200374.4]
  wire  OptimizationBarrier_19_io_y_sw; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@200374.4]
  wire  OptimizationBarrier_19_io_y_sx; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@200374.4]
  wire  OptimizationBarrier_19_io_y_sr; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@200374.4]
  wire  OptimizationBarrier_19_io_y_pw; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@200374.4]
  wire  OptimizationBarrier_19_io_y_px; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@200374.4]
  wire  OptimizationBarrier_19_io_y_pr; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@200374.4]
  wire  OptimizationBarrier_19_io_y_ppp; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@200374.4]
  wire  OptimizationBarrier_19_io_y_pal; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@200374.4]
  wire  OptimizationBarrier_19_io_y_paa; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@200374.4]
  wire  OptimizationBarrier_19_io_y_eff; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@200374.4]
  wire  OptimizationBarrier_19_io_y_c; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@200374.4]
  wire [19:0] OptimizationBarrier_20_io_x_ppn; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@200417.4]
  wire  OptimizationBarrier_20_io_x_u; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@200417.4]
  wire  OptimizationBarrier_20_io_x_ae; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@200417.4]
  wire  OptimizationBarrier_20_io_x_sw; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@200417.4]
  wire  OptimizationBarrier_20_io_x_sx; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@200417.4]
  wire  OptimizationBarrier_20_io_x_sr; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@200417.4]
  wire  OptimizationBarrier_20_io_x_pw; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@200417.4]
  wire  OptimizationBarrier_20_io_x_px; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@200417.4]
  wire  OptimizationBarrier_20_io_x_pr; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@200417.4]
  wire  OptimizationBarrier_20_io_x_ppp; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@200417.4]
  wire  OptimizationBarrier_20_io_x_pal; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@200417.4]
  wire  OptimizationBarrier_20_io_x_paa; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@200417.4]
  wire  OptimizationBarrier_20_io_x_eff; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@200417.4]
  wire  OptimizationBarrier_20_io_x_c; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@200417.4]
  wire [19:0] OptimizationBarrier_20_io_y_ppn; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@200417.4]
  wire  OptimizationBarrier_20_io_y_u; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@200417.4]
  wire  OptimizationBarrier_20_io_y_ae; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@200417.4]
  wire  OptimizationBarrier_20_io_y_sw; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@200417.4]
  wire  OptimizationBarrier_20_io_y_sx; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@200417.4]
  wire  OptimizationBarrier_20_io_y_sr; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@200417.4]
  wire  OptimizationBarrier_20_io_y_pw; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@200417.4]
  wire  OptimizationBarrier_20_io_y_px; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@200417.4]
  wire  OptimizationBarrier_20_io_y_pr; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@200417.4]
  wire  OptimizationBarrier_20_io_y_ppp; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@200417.4]
  wire  OptimizationBarrier_20_io_y_pal; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@200417.4]
  wire  OptimizationBarrier_20_io_y_paa; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@200417.4]
  wire  OptimizationBarrier_20_io_y_eff; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@200417.4]
  wire  OptimizationBarrier_20_io_y_c; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@200417.4]
  wire [19:0] OptimizationBarrier_21_io_x_ppn; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@200460.4]
  wire  OptimizationBarrier_21_io_x_u; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@200460.4]
  wire  OptimizationBarrier_21_io_x_ae; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@200460.4]
  wire  OptimizationBarrier_21_io_x_sw; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@200460.4]
  wire  OptimizationBarrier_21_io_x_sx; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@200460.4]
  wire  OptimizationBarrier_21_io_x_sr; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@200460.4]
  wire  OptimizationBarrier_21_io_x_pw; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@200460.4]
  wire  OptimizationBarrier_21_io_x_px; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@200460.4]
  wire  OptimizationBarrier_21_io_x_pr; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@200460.4]
  wire  OptimizationBarrier_21_io_x_ppp; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@200460.4]
  wire  OptimizationBarrier_21_io_x_pal; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@200460.4]
  wire  OptimizationBarrier_21_io_x_paa; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@200460.4]
  wire  OptimizationBarrier_21_io_x_eff; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@200460.4]
  wire  OptimizationBarrier_21_io_x_c; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@200460.4]
  wire [19:0] OptimizationBarrier_21_io_y_ppn; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@200460.4]
  wire  OptimizationBarrier_21_io_y_u; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@200460.4]
  wire  OptimizationBarrier_21_io_y_ae; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@200460.4]
  wire  OptimizationBarrier_21_io_y_sw; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@200460.4]
  wire  OptimizationBarrier_21_io_y_sx; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@200460.4]
  wire  OptimizationBarrier_21_io_y_sr; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@200460.4]
  wire  OptimizationBarrier_21_io_y_pw; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@200460.4]
  wire  OptimizationBarrier_21_io_y_px; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@200460.4]
  wire  OptimizationBarrier_21_io_y_pr; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@200460.4]
  wire  OptimizationBarrier_21_io_y_ppp; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@200460.4]
  wire  OptimizationBarrier_21_io_y_pal; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@200460.4]
  wire  OptimizationBarrier_21_io_y_paa; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@200460.4]
  wire  OptimizationBarrier_21_io_y_eff; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@200460.4]
  wire  OptimizationBarrier_21_io_y_c; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@200460.4]
  wire [19:0] OptimizationBarrier_22_io_x_ppn; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@200502.4]
  wire  OptimizationBarrier_22_io_x_u; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@200502.4]
  wire  OptimizationBarrier_22_io_x_ae; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@200502.4]
  wire  OptimizationBarrier_22_io_x_sw; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@200502.4]
  wire  OptimizationBarrier_22_io_x_sx; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@200502.4]
  wire  OptimizationBarrier_22_io_x_sr; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@200502.4]
  wire  OptimizationBarrier_22_io_x_pw; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@200502.4]
  wire  OptimizationBarrier_22_io_x_px; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@200502.4]
  wire  OptimizationBarrier_22_io_x_pr; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@200502.4]
  wire  OptimizationBarrier_22_io_x_ppp; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@200502.4]
  wire  OptimizationBarrier_22_io_x_pal; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@200502.4]
  wire  OptimizationBarrier_22_io_x_paa; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@200502.4]
  wire  OptimizationBarrier_22_io_x_eff; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@200502.4]
  wire  OptimizationBarrier_22_io_x_c; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@200502.4]
  wire [19:0] OptimizationBarrier_22_io_y_ppn; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@200502.4]
  wire  OptimizationBarrier_22_io_y_u; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@200502.4]
  wire  OptimizationBarrier_22_io_y_ae; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@200502.4]
  wire  OptimizationBarrier_22_io_y_sw; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@200502.4]
  wire  OptimizationBarrier_22_io_y_sx; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@200502.4]
  wire  OptimizationBarrier_22_io_y_sr; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@200502.4]
  wire  OptimizationBarrier_22_io_y_pw; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@200502.4]
  wire  OptimizationBarrier_22_io_y_px; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@200502.4]
  wire  OptimizationBarrier_22_io_y_pr; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@200502.4]
  wire  OptimizationBarrier_22_io_y_ppp; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@200502.4]
  wire  OptimizationBarrier_22_io_y_pal; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@200502.4]
  wire  OptimizationBarrier_22_io_y_paa; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@200502.4]
  wire  OptimizationBarrier_22_io_y_eff; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@200502.4]
  wire  OptimizationBarrier_22_io_y_c; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@200502.4]
  wire [19:0] OptimizationBarrier_23_io_x_ppn; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@200544.4]
  wire  OptimizationBarrier_23_io_x_u; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@200544.4]
  wire  OptimizationBarrier_23_io_x_ae; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@200544.4]
  wire  OptimizationBarrier_23_io_x_sw; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@200544.4]
  wire  OptimizationBarrier_23_io_x_sx; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@200544.4]
  wire  OptimizationBarrier_23_io_x_sr; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@200544.4]
  wire  OptimizationBarrier_23_io_x_pw; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@200544.4]
  wire  OptimizationBarrier_23_io_x_px; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@200544.4]
  wire  OptimizationBarrier_23_io_x_pr; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@200544.4]
  wire  OptimizationBarrier_23_io_x_ppp; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@200544.4]
  wire  OptimizationBarrier_23_io_x_pal; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@200544.4]
  wire  OptimizationBarrier_23_io_x_paa; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@200544.4]
  wire  OptimizationBarrier_23_io_x_eff; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@200544.4]
  wire  OptimizationBarrier_23_io_x_c; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@200544.4]
  wire [19:0] OptimizationBarrier_23_io_y_ppn; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@200544.4]
  wire  OptimizationBarrier_23_io_y_u; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@200544.4]
  wire  OptimizationBarrier_23_io_y_ae; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@200544.4]
  wire  OptimizationBarrier_23_io_y_sw; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@200544.4]
  wire  OptimizationBarrier_23_io_y_sx; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@200544.4]
  wire  OptimizationBarrier_23_io_y_sr; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@200544.4]
  wire  OptimizationBarrier_23_io_y_pw; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@200544.4]
  wire  OptimizationBarrier_23_io_y_px; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@200544.4]
  wire  OptimizationBarrier_23_io_y_pr; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@200544.4]
  wire  OptimizationBarrier_23_io_y_ppp; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@200544.4]
  wire  OptimizationBarrier_23_io_y_pal; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@200544.4]
  wire  OptimizationBarrier_23_io_y_paa; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@200544.4]
  wire  OptimizationBarrier_23_io_y_eff; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@200544.4]
  wire  OptimizationBarrier_23_io_y_c; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@200544.4]
  wire [19:0] OptimizationBarrier_24_io_x_ppn; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@200586.4]
  wire  OptimizationBarrier_24_io_x_u; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@200586.4]
  wire  OptimizationBarrier_24_io_x_ae; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@200586.4]
  wire  OptimizationBarrier_24_io_x_sw; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@200586.4]
  wire  OptimizationBarrier_24_io_x_sx; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@200586.4]
  wire  OptimizationBarrier_24_io_x_sr; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@200586.4]
  wire  OptimizationBarrier_24_io_x_pw; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@200586.4]
  wire  OptimizationBarrier_24_io_x_px; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@200586.4]
  wire  OptimizationBarrier_24_io_x_pr; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@200586.4]
  wire  OptimizationBarrier_24_io_x_ppp; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@200586.4]
  wire  OptimizationBarrier_24_io_x_pal; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@200586.4]
  wire  OptimizationBarrier_24_io_x_paa; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@200586.4]
  wire  OptimizationBarrier_24_io_x_eff; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@200586.4]
  wire  OptimizationBarrier_24_io_x_c; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@200586.4]
  wire [19:0] OptimizationBarrier_24_io_y_ppn; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@200586.4]
  wire  OptimizationBarrier_24_io_y_u; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@200586.4]
  wire  OptimizationBarrier_24_io_y_ae; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@200586.4]
  wire  OptimizationBarrier_24_io_y_sw; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@200586.4]
  wire  OptimizationBarrier_24_io_y_sx; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@200586.4]
  wire  OptimizationBarrier_24_io_y_sr; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@200586.4]
  wire  OptimizationBarrier_24_io_y_pw; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@200586.4]
  wire  OptimizationBarrier_24_io_y_px; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@200586.4]
  wire  OptimizationBarrier_24_io_y_pr; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@200586.4]
  wire  OptimizationBarrier_24_io_y_ppp; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@200586.4]
  wire  OptimizationBarrier_24_io_y_pal; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@200586.4]
  wire  OptimizationBarrier_24_io_y_paa; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@200586.4]
  wire  OptimizationBarrier_24_io_y_eff; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@200586.4]
  wire  OptimizationBarrier_24_io_y_c; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@200586.4]
  wire [19:0] OptimizationBarrier_25_io_x_ppn; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@200628.4]
  wire  OptimizationBarrier_25_io_x_u; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@200628.4]
  wire  OptimizationBarrier_25_io_x_ae; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@200628.4]
  wire  OptimizationBarrier_25_io_x_sw; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@200628.4]
  wire  OptimizationBarrier_25_io_x_sx; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@200628.4]
  wire  OptimizationBarrier_25_io_x_sr; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@200628.4]
  wire  OptimizationBarrier_25_io_x_pw; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@200628.4]
  wire  OptimizationBarrier_25_io_x_px; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@200628.4]
  wire  OptimizationBarrier_25_io_x_pr; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@200628.4]
  wire  OptimizationBarrier_25_io_x_ppp; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@200628.4]
  wire  OptimizationBarrier_25_io_x_pal; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@200628.4]
  wire  OptimizationBarrier_25_io_x_paa; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@200628.4]
  wire  OptimizationBarrier_25_io_x_eff; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@200628.4]
  wire  OptimizationBarrier_25_io_x_c; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@200628.4]
  wire [19:0] OptimizationBarrier_25_io_y_ppn; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@200628.4]
  wire  OptimizationBarrier_25_io_y_u; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@200628.4]
  wire  OptimizationBarrier_25_io_y_ae; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@200628.4]
  wire  OptimizationBarrier_25_io_y_sw; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@200628.4]
  wire  OptimizationBarrier_25_io_y_sx; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@200628.4]
  wire  OptimizationBarrier_25_io_y_sr; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@200628.4]
  wire  OptimizationBarrier_25_io_y_pw; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@200628.4]
  wire  OptimizationBarrier_25_io_y_px; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@200628.4]
  wire  OptimizationBarrier_25_io_y_pr; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@200628.4]
  wire  OptimizationBarrier_25_io_y_ppp; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@200628.4]
  wire  OptimizationBarrier_25_io_y_pal; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@200628.4]
  wire  OptimizationBarrier_25_io_y_paa; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@200628.4]
  wire  OptimizationBarrier_25_io_y_eff; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@200628.4]
  wire  OptimizationBarrier_25_io_y_c; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@200628.4]
  wire [19:0] OptimizationBarrier_26_io_x_ppn; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@200670.4]
  wire  OptimizationBarrier_26_io_x_u; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@200670.4]
  wire  OptimizationBarrier_26_io_x_ae; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@200670.4]
  wire  OptimizationBarrier_26_io_x_sw; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@200670.4]
  wire  OptimizationBarrier_26_io_x_sx; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@200670.4]
  wire  OptimizationBarrier_26_io_x_sr; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@200670.4]
  wire  OptimizationBarrier_26_io_x_pw; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@200670.4]
  wire  OptimizationBarrier_26_io_x_px; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@200670.4]
  wire  OptimizationBarrier_26_io_x_pr; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@200670.4]
  wire  OptimizationBarrier_26_io_x_ppp; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@200670.4]
  wire  OptimizationBarrier_26_io_x_pal; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@200670.4]
  wire  OptimizationBarrier_26_io_x_paa; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@200670.4]
  wire  OptimizationBarrier_26_io_x_eff; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@200670.4]
  wire  OptimizationBarrier_26_io_x_c; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@200670.4]
  wire [19:0] OptimizationBarrier_26_io_y_ppn; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@200670.4]
  wire  OptimizationBarrier_26_io_y_u; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@200670.4]
  wire  OptimizationBarrier_26_io_y_ae; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@200670.4]
  wire  OptimizationBarrier_26_io_y_sw; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@200670.4]
  wire  OptimizationBarrier_26_io_y_sx; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@200670.4]
  wire  OptimizationBarrier_26_io_y_sr; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@200670.4]
  wire  OptimizationBarrier_26_io_y_pw; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@200670.4]
  wire  OptimizationBarrier_26_io_y_px; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@200670.4]
  wire  OptimizationBarrier_26_io_y_pr; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@200670.4]
  wire  OptimizationBarrier_26_io_y_ppp; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@200670.4]
  wire  OptimizationBarrier_26_io_y_pal; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@200670.4]
  wire  OptimizationBarrier_26_io_y_paa; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@200670.4]
  wire  OptimizationBarrier_26_io_y_eff; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@200670.4]
  wire  OptimizationBarrier_26_io_y_c; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@200670.4]
  wire [19:0] OptimizationBarrier_27_io_x_ppn; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@200713.4]
  wire  OptimizationBarrier_27_io_x_u; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@200713.4]
  wire  OptimizationBarrier_27_io_x_ae; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@200713.4]
  wire  OptimizationBarrier_27_io_x_sw; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@200713.4]
  wire  OptimizationBarrier_27_io_x_sx; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@200713.4]
  wire  OptimizationBarrier_27_io_x_sr; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@200713.4]
  wire  OptimizationBarrier_27_io_x_pw; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@200713.4]
  wire  OptimizationBarrier_27_io_x_px; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@200713.4]
  wire  OptimizationBarrier_27_io_x_pr; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@200713.4]
  wire  OptimizationBarrier_27_io_x_ppp; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@200713.4]
  wire  OptimizationBarrier_27_io_x_pal; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@200713.4]
  wire  OptimizationBarrier_27_io_x_paa; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@200713.4]
  wire  OptimizationBarrier_27_io_x_eff; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@200713.4]
  wire  OptimizationBarrier_27_io_x_c; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@200713.4]
  wire [19:0] OptimizationBarrier_27_io_y_ppn; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@200713.4]
  wire  OptimizationBarrier_27_io_y_u; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@200713.4]
  wire  OptimizationBarrier_27_io_y_ae; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@200713.4]
  wire  OptimizationBarrier_27_io_y_sw; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@200713.4]
  wire  OptimizationBarrier_27_io_y_sx; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@200713.4]
  wire  OptimizationBarrier_27_io_y_sr; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@200713.4]
  wire  OptimizationBarrier_27_io_y_pw; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@200713.4]
  wire  OptimizationBarrier_27_io_y_px; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@200713.4]
  wire  OptimizationBarrier_27_io_y_pr; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@200713.4]
  wire  OptimizationBarrier_27_io_y_ppp; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@200713.4]
  wire  OptimizationBarrier_27_io_y_pal; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@200713.4]
  wire  OptimizationBarrier_27_io_y_paa; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@200713.4]
  wire  OptimizationBarrier_27_io_y_eff; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@200713.4]
  wire  OptimizationBarrier_27_io_y_c; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@200713.4]
  wire [19:0] OptimizationBarrier_28_io_x_ppn; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@200756.4]
  wire  OptimizationBarrier_28_io_x_u; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@200756.4]
  wire  OptimizationBarrier_28_io_x_ae; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@200756.4]
  wire  OptimizationBarrier_28_io_x_sw; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@200756.4]
  wire  OptimizationBarrier_28_io_x_sx; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@200756.4]
  wire  OptimizationBarrier_28_io_x_sr; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@200756.4]
  wire  OptimizationBarrier_28_io_x_pw; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@200756.4]
  wire  OptimizationBarrier_28_io_x_px; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@200756.4]
  wire  OptimizationBarrier_28_io_x_pr; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@200756.4]
  wire  OptimizationBarrier_28_io_x_ppp; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@200756.4]
  wire  OptimizationBarrier_28_io_x_pal; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@200756.4]
  wire  OptimizationBarrier_28_io_x_paa; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@200756.4]
  wire  OptimizationBarrier_28_io_x_eff; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@200756.4]
  wire  OptimizationBarrier_28_io_x_c; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@200756.4]
  wire [19:0] OptimizationBarrier_28_io_y_ppn; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@200756.4]
  wire  OptimizationBarrier_28_io_y_u; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@200756.4]
  wire  OptimizationBarrier_28_io_y_ae; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@200756.4]
  wire  OptimizationBarrier_28_io_y_sw; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@200756.4]
  wire  OptimizationBarrier_28_io_y_sx; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@200756.4]
  wire  OptimizationBarrier_28_io_y_sr; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@200756.4]
  wire  OptimizationBarrier_28_io_y_pw; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@200756.4]
  wire  OptimizationBarrier_28_io_y_px; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@200756.4]
  wire  OptimizationBarrier_28_io_y_pr; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@200756.4]
  wire  OptimizationBarrier_28_io_y_ppp; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@200756.4]
  wire  OptimizationBarrier_28_io_y_pal; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@200756.4]
  wire  OptimizationBarrier_28_io_y_paa; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@200756.4]
  wire  OptimizationBarrier_28_io_y_eff; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@200756.4]
  wire  OptimizationBarrier_28_io_y_c; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@200756.4]
  wire [19:0] OptimizationBarrier_29_io_x_ppn; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@200799.4]
  wire  OptimizationBarrier_29_io_x_u; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@200799.4]
  wire  OptimizationBarrier_29_io_x_ae; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@200799.4]
  wire  OptimizationBarrier_29_io_x_sw; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@200799.4]
  wire  OptimizationBarrier_29_io_x_sx; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@200799.4]
  wire  OptimizationBarrier_29_io_x_sr; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@200799.4]
  wire  OptimizationBarrier_29_io_x_pw; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@200799.4]
  wire  OptimizationBarrier_29_io_x_px; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@200799.4]
  wire  OptimizationBarrier_29_io_x_pr; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@200799.4]
  wire  OptimizationBarrier_29_io_x_ppp; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@200799.4]
  wire  OptimizationBarrier_29_io_x_pal; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@200799.4]
  wire  OptimizationBarrier_29_io_x_paa; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@200799.4]
  wire  OptimizationBarrier_29_io_x_eff; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@200799.4]
  wire  OptimizationBarrier_29_io_x_c; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@200799.4]
  wire [19:0] OptimizationBarrier_29_io_y_ppn; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@200799.4]
  wire  OptimizationBarrier_29_io_y_u; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@200799.4]
  wire  OptimizationBarrier_29_io_y_ae; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@200799.4]
  wire  OptimizationBarrier_29_io_y_sw; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@200799.4]
  wire  OptimizationBarrier_29_io_y_sx; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@200799.4]
  wire  OptimizationBarrier_29_io_y_sr; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@200799.4]
  wire  OptimizationBarrier_29_io_y_pw; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@200799.4]
  wire  OptimizationBarrier_29_io_y_px; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@200799.4]
  wire  OptimizationBarrier_29_io_y_pr; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@200799.4]
  wire  OptimizationBarrier_29_io_y_ppp; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@200799.4]
  wire  OptimizationBarrier_29_io_y_pal; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@200799.4]
  wire  OptimizationBarrier_29_io_y_paa; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@200799.4]
  wire  OptimizationBarrier_29_io_y_eff; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@200799.4]
  wire  OptimizationBarrier_29_io_y_c; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@200799.4]
  wire [19:0] OptimizationBarrier_30_io_x_ppn; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@200842.4]
  wire  OptimizationBarrier_30_io_x_u; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@200842.4]
  wire  OptimizationBarrier_30_io_x_ae; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@200842.4]
  wire  OptimizationBarrier_30_io_x_sw; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@200842.4]
  wire  OptimizationBarrier_30_io_x_sx; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@200842.4]
  wire  OptimizationBarrier_30_io_x_sr; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@200842.4]
  wire  OptimizationBarrier_30_io_x_pw; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@200842.4]
  wire  OptimizationBarrier_30_io_x_px; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@200842.4]
  wire  OptimizationBarrier_30_io_x_pr; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@200842.4]
  wire  OptimizationBarrier_30_io_x_ppp; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@200842.4]
  wire  OptimizationBarrier_30_io_x_pal; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@200842.4]
  wire  OptimizationBarrier_30_io_x_paa; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@200842.4]
  wire  OptimizationBarrier_30_io_x_eff; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@200842.4]
  wire  OptimizationBarrier_30_io_x_c; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@200842.4]
  wire [19:0] OptimizationBarrier_30_io_y_ppn; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@200842.4]
  wire  OptimizationBarrier_30_io_y_u; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@200842.4]
  wire  OptimizationBarrier_30_io_y_ae; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@200842.4]
  wire  OptimizationBarrier_30_io_y_sw; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@200842.4]
  wire  OptimizationBarrier_30_io_y_sx; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@200842.4]
  wire  OptimizationBarrier_30_io_y_sr; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@200842.4]
  wire  OptimizationBarrier_30_io_y_pw; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@200842.4]
  wire  OptimizationBarrier_30_io_y_px; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@200842.4]
  wire  OptimizationBarrier_30_io_y_pr; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@200842.4]
  wire  OptimizationBarrier_30_io_y_ppp; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@200842.4]
  wire  OptimizationBarrier_30_io_y_pal; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@200842.4]
  wire  OptimizationBarrier_30_io_y_paa; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@200842.4]
  wire  OptimizationBarrier_30_io_y_eff; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@200842.4]
  wire  OptimizationBarrier_30_io_y_c; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@200842.4]
  wire [19:0] OptimizationBarrier_31_io_x_ppn; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@200885.4]
  wire  OptimizationBarrier_31_io_x_u; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@200885.4]
  wire  OptimizationBarrier_31_io_x_ae; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@200885.4]
  wire  OptimizationBarrier_31_io_x_sw; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@200885.4]
  wire  OptimizationBarrier_31_io_x_sx; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@200885.4]
  wire  OptimizationBarrier_31_io_x_sr; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@200885.4]
  wire  OptimizationBarrier_31_io_x_pw; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@200885.4]
  wire  OptimizationBarrier_31_io_x_px; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@200885.4]
  wire  OptimizationBarrier_31_io_x_pr; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@200885.4]
  wire  OptimizationBarrier_31_io_x_ppp; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@200885.4]
  wire  OptimizationBarrier_31_io_x_pal; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@200885.4]
  wire  OptimizationBarrier_31_io_x_paa; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@200885.4]
  wire  OptimizationBarrier_31_io_x_eff; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@200885.4]
  wire  OptimizationBarrier_31_io_x_c; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@200885.4]
  wire [19:0] OptimizationBarrier_31_io_y_ppn; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@200885.4]
  wire  OptimizationBarrier_31_io_y_u; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@200885.4]
  wire  OptimizationBarrier_31_io_y_ae; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@200885.4]
  wire  OptimizationBarrier_31_io_y_sw; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@200885.4]
  wire  OptimizationBarrier_31_io_y_sx; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@200885.4]
  wire  OptimizationBarrier_31_io_y_sr; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@200885.4]
  wire  OptimizationBarrier_31_io_y_pw; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@200885.4]
  wire  OptimizationBarrier_31_io_y_px; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@200885.4]
  wire  OptimizationBarrier_31_io_y_pr; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@200885.4]
  wire  OptimizationBarrier_31_io_y_ppp; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@200885.4]
  wire  OptimizationBarrier_31_io_y_pal; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@200885.4]
  wire  OptimizationBarrier_31_io_y_paa; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@200885.4]
  wire  OptimizationBarrier_31_io_y_eff; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@200885.4]
  wire  OptimizationBarrier_31_io_y_c; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@200885.4]
  wire [19:0] OptimizationBarrier_32_io_x_ppn; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@200928.4]
  wire  OptimizationBarrier_32_io_x_u; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@200928.4]
  wire  OptimizationBarrier_32_io_x_ae; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@200928.4]
  wire  OptimizationBarrier_32_io_x_sw; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@200928.4]
  wire  OptimizationBarrier_32_io_x_sx; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@200928.4]
  wire  OptimizationBarrier_32_io_x_sr; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@200928.4]
  wire  OptimizationBarrier_32_io_x_pw; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@200928.4]
  wire  OptimizationBarrier_32_io_x_px; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@200928.4]
  wire  OptimizationBarrier_32_io_x_pr; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@200928.4]
  wire  OptimizationBarrier_32_io_x_ppp; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@200928.4]
  wire  OptimizationBarrier_32_io_x_pal; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@200928.4]
  wire  OptimizationBarrier_32_io_x_paa; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@200928.4]
  wire  OptimizationBarrier_32_io_x_eff; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@200928.4]
  wire  OptimizationBarrier_32_io_x_c; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@200928.4]
  wire [19:0] OptimizationBarrier_32_io_y_ppn; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@200928.4]
  wire  OptimizationBarrier_32_io_y_u; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@200928.4]
  wire  OptimizationBarrier_32_io_y_ae; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@200928.4]
  wire  OptimizationBarrier_32_io_y_sw; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@200928.4]
  wire  OptimizationBarrier_32_io_y_sx; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@200928.4]
  wire  OptimizationBarrier_32_io_y_sr; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@200928.4]
  wire  OptimizationBarrier_32_io_y_pw; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@200928.4]
  wire  OptimizationBarrier_32_io_y_px; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@200928.4]
  wire  OptimizationBarrier_32_io_y_pr; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@200928.4]
  wire  OptimizationBarrier_32_io_y_ppp; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@200928.4]
  wire  OptimizationBarrier_32_io_y_pal; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@200928.4]
  wire  OptimizationBarrier_32_io_y_paa; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@200928.4]
  wire  OptimizationBarrier_32_io_y_eff; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@200928.4]
  wire  OptimizationBarrier_32_io_y_c; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@200928.4]
  wire [19:0] OptimizationBarrier_33_io_x_ppn; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@200971.4]
  wire  OptimizationBarrier_33_io_x_u; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@200971.4]
  wire  OptimizationBarrier_33_io_x_ae; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@200971.4]
  wire  OptimizationBarrier_33_io_x_sw; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@200971.4]
  wire  OptimizationBarrier_33_io_x_sx; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@200971.4]
  wire  OptimizationBarrier_33_io_x_sr; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@200971.4]
  wire  OptimizationBarrier_33_io_x_pw; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@200971.4]
  wire  OptimizationBarrier_33_io_x_px; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@200971.4]
  wire  OptimizationBarrier_33_io_x_pr; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@200971.4]
  wire  OptimizationBarrier_33_io_x_ppp; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@200971.4]
  wire  OptimizationBarrier_33_io_x_pal; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@200971.4]
  wire  OptimizationBarrier_33_io_x_paa; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@200971.4]
  wire  OptimizationBarrier_33_io_x_eff; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@200971.4]
  wire  OptimizationBarrier_33_io_x_c; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@200971.4]
  wire [19:0] OptimizationBarrier_33_io_y_ppn; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@200971.4]
  wire  OptimizationBarrier_33_io_y_u; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@200971.4]
  wire  OptimizationBarrier_33_io_y_ae; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@200971.4]
  wire  OptimizationBarrier_33_io_y_sw; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@200971.4]
  wire  OptimizationBarrier_33_io_y_sx; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@200971.4]
  wire  OptimizationBarrier_33_io_y_sr; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@200971.4]
  wire  OptimizationBarrier_33_io_y_pw; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@200971.4]
  wire  OptimizationBarrier_33_io_y_px; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@200971.4]
  wire  OptimizationBarrier_33_io_y_pr; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@200971.4]
  wire  OptimizationBarrier_33_io_y_ppp; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@200971.4]
  wire  OptimizationBarrier_33_io_y_pal; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@200971.4]
  wire  OptimizationBarrier_33_io_y_paa; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@200971.4]
  wire  OptimizationBarrier_33_io_y_eff; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@200971.4]
  wire  OptimizationBarrier_33_io_y_c; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@200971.4]
  wire [19:0] OptimizationBarrier_34_io_x_ppn; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@201014.4]
  wire  OptimizationBarrier_34_io_x_u; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@201014.4]
  wire  OptimizationBarrier_34_io_x_ae; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@201014.4]
  wire  OptimizationBarrier_34_io_x_sw; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@201014.4]
  wire  OptimizationBarrier_34_io_x_sx; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@201014.4]
  wire  OptimizationBarrier_34_io_x_sr; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@201014.4]
  wire  OptimizationBarrier_34_io_x_pw; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@201014.4]
  wire  OptimizationBarrier_34_io_x_px; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@201014.4]
  wire  OptimizationBarrier_34_io_x_pr; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@201014.4]
  wire  OptimizationBarrier_34_io_x_ppp; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@201014.4]
  wire  OptimizationBarrier_34_io_x_pal; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@201014.4]
  wire  OptimizationBarrier_34_io_x_paa; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@201014.4]
  wire  OptimizationBarrier_34_io_x_eff; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@201014.4]
  wire  OptimizationBarrier_34_io_x_c; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@201014.4]
  wire [19:0] OptimizationBarrier_34_io_y_ppn; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@201014.4]
  wire  OptimizationBarrier_34_io_y_u; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@201014.4]
  wire  OptimizationBarrier_34_io_y_ae; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@201014.4]
  wire  OptimizationBarrier_34_io_y_sw; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@201014.4]
  wire  OptimizationBarrier_34_io_y_sx; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@201014.4]
  wire  OptimizationBarrier_34_io_y_sr; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@201014.4]
  wire  OptimizationBarrier_34_io_y_pw; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@201014.4]
  wire  OptimizationBarrier_34_io_y_px; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@201014.4]
  wire  OptimizationBarrier_34_io_y_pr; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@201014.4]
  wire  OptimizationBarrier_34_io_y_ppp; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@201014.4]
  wire  OptimizationBarrier_34_io_y_pal; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@201014.4]
  wire  OptimizationBarrier_34_io_y_paa; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@201014.4]
  wire  OptimizationBarrier_34_io_y_eff; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@201014.4]
  wire  OptimizationBarrier_34_io_y_c; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@201014.4]
  wire [19:0] OptimizationBarrier_35_io_x_ppn; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@201056.4]
  wire  OptimizationBarrier_35_io_x_u; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@201056.4]
  wire  OptimizationBarrier_35_io_x_ae; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@201056.4]
  wire  OptimizationBarrier_35_io_x_sw; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@201056.4]
  wire  OptimizationBarrier_35_io_x_sx; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@201056.4]
  wire  OptimizationBarrier_35_io_x_sr; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@201056.4]
  wire  OptimizationBarrier_35_io_x_pw; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@201056.4]
  wire  OptimizationBarrier_35_io_x_px; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@201056.4]
  wire  OptimizationBarrier_35_io_x_pr; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@201056.4]
  wire  OptimizationBarrier_35_io_x_ppp; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@201056.4]
  wire  OptimizationBarrier_35_io_x_pal; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@201056.4]
  wire  OptimizationBarrier_35_io_x_paa; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@201056.4]
  wire  OptimizationBarrier_35_io_x_eff; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@201056.4]
  wire  OptimizationBarrier_35_io_x_c; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@201056.4]
  wire [19:0] OptimizationBarrier_35_io_y_ppn; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@201056.4]
  wire  OptimizationBarrier_35_io_y_u; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@201056.4]
  wire  OptimizationBarrier_35_io_y_ae; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@201056.4]
  wire  OptimizationBarrier_35_io_y_sw; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@201056.4]
  wire  OptimizationBarrier_35_io_y_sx; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@201056.4]
  wire  OptimizationBarrier_35_io_y_sr; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@201056.4]
  wire  OptimizationBarrier_35_io_y_pw; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@201056.4]
  wire  OptimizationBarrier_35_io_y_px; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@201056.4]
  wire  OptimizationBarrier_35_io_y_pr; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@201056.4]
  wire  OptimizationBarrier_35_io_y_ppp; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@201056.4]
  wire  OptimizationBarrier_35_io_y_pal; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@201056.4]
  wire  OptimizationBarrier_35_io_y_paa; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@201056.4]
  wire  OptimizationBarrier_35_io_y_eff; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@201056.4]
  wire  OptimizationBarrier_35_io_y_c; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@201056.4]
  wire [19:0] OptimizationBarrier_36_io_x_ppn; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@201098.4]
  wire  OptimizationBarrier_36_io_x_u; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@201098.4]
  wire  OptimizationBarrier_36_io_x_ae; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@201098.4]
  wire  OptimizationBarrier_36_io_x_sw; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@201098.4]
  wire  OptimizationBarrier_36_io_x_sx; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@201098.4]
  wire  OptimizationBarrier_36_io_x_sr; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@201098.4]
  wire  OptimizationBarrier_36_io_x_pw; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@201098.4]
  wire  OptimizationBarrier_36_io_x_px; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@201098.4]
  wire  OptimizationBarrier_36_io_x_pr; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@201098.4]
  wire  OptimizationBarrier_36_io_x_ppp; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@201098.4]
  wire  OptimizationBarrier_36_io_x_pal; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@201098.4]
  wire  OptimizationBarrier_36_io_x_paa; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@201098.4]
  wire  OptimizationBarrier_36_io_x_eff; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@201098.4]
  wire  OptimizationBarrier_36_io_x_c; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@201098.4]
  wire [19:0] OptimizationBarrier_36_io_y_ppn; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@201098.4]
  wire  OptimizationBarrier_36_io_y_u; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@201098.4]
  wire  OptimizationBarrier_36_io_y_ae; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@201098.4]
  wire  OptimizationBarrier_36_io_y_sw; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@201098.4]
  wire  OptimizationBarrier_36_io_y_sx; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@201098.4]
  wire  OptimizationBarrier_36_io_y_sr; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@201098.4]
  wire  OptimizationBarrier_36_io_y_pw; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@201098.4]
  wire  OptimizationBarrier_36_io_y_px; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@201098.4]
  wire  OptimizationBarrier_36_io_y_pr; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@201098.4]
  wire  OptimizationBarrier_36_io_y_ppp; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@201098.4]
  wire  OptimizationBarrier_36_io_y_pal; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@201098.4]
  wire  OptimizationBarrier_36_io_y_paa; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@201098.4]
  wire  OptimizationBarrier_36_io_y_eff; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@201098.4]
  wire  OptimizationBarrier_36_io_y_c; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@201098.4]
  wire [19:0] OptimizationBarrier_37_io_x_ppn; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@201140.4]
  wire  OptimizationBarrier_37_io_x_u; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@201140.4]
  wire  OptimizationBarrier_37_io_x_ae; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@201140.4]
  wire  OptimizationBarrier_37_io_x_sw; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@201140.4]
  wire  OptimizationBarrier_37_io_x_sx; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@201140.4]
  wire  OptimizationBarrier_37_io_x_sr; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@201140.4]
  wire  OptimizationBarrier_37_io_x_pw; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@201140.4]
  wire  OptimizationBarrier_37_io_x_px; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@201140.4]
  wire  OptimizationBarrier_37_io_x_pr; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@201140.4]
  wire  OptimizationBarrier_37_io_x_ppp; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@201140.4]
  wire  OptimizationBarrier_37_io_x_pal; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@201140.4]
  wire  OptimizationBarrier_37_io_x_paa; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@201140.4]
  wire  OptimizationBarrier_37_io_x_eff; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@201140.4]
  wire  OptimizationBarrier_37_io_x_c; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@201140.4]
  wire [19:0] OptimizationBarrier_37_io_y_ppn; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@201140.4]
  wire  OptimizationBarrier_37_io_y_u; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@201140.4]
  wire  OptimizationBarrier_37_io_y_ae; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@201140.4]
  wire  OptimizationBarrier_37_io_y_sw; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@201140.4]
  wire  OptimizationBarrier_37_io_y_sx; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@201140.4]
  wire  OptimizationBarrier_37_io_y_sr; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@201140.4]
  wire  OptimizationBarrier_37_io_y_pw; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@201140.4]
  wire  OptimizationBarrier_37_io_y_px; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@201140.4]
  wire  OptimizationBarrier_37_io_y_pr; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@201140.4]
  wire  OptimizationBarrier_37_io_y_ppp; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@201140.4]
  wire  OptimizationBarrier_37_io_y_pal; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@201140.4]
  wire  OptimizationBarrier_37_io_y_paa; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@201140.4]
  wire  OptimizationBarrier_37_io_y_eff; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@201140.4]
  wire  OptimizationBarrier_37_io_y_c; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@201140.4]
  wire [19:0] OptimizationBarrier_38_io_x_ppn; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@201182.4]
  wire  OptimizationBarrier_38_io_x_u; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@201182.4]
  wire  OptimizationBarrier_38_io_x_ae; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@201182.4]
  wire  OptimizationBarrier_38_io_x_sw; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@201182.4]
  wire  OptimizationBarrier_38_io_x_sx; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@201182.4]
  wire  OptimizationBarrier_38_io_x_sr; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@201182.4]
  wire  OptimizationBarrier_38_io_x_pw; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@201182.4]
  wire  OptimizationBarrier_38_io_x_px; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@201182.4]
  wire  OptimizationBarrier_38_io_x_pr; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@201182.4]
  wire  OptimizationBarrier_38_io_x_ppp; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@201182.4]
  wire  OptimizationBarrier_38_io_x_pal; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@201182.4]
  wire  OptimizationBarrier_38_io_x_paa; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@201182.4]
  wire  OptimizationBarrier_38_io_x_eff; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@201182.4]
  wire  OptimizationBarrier_38_io_x_c; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@201182.4]
  wire [19:0] OptimizationBarrier_38_io_y_ppn; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@201182.4]
  wire  OptimizationBarrier_38_io_y_u; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@201182.4]
  wire  OptimizationBarrier_38_io_y_ae; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@201182.4]
  wire  OptimizationBarrier_38_io_y_sw; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@201182.4]
  wire  OptimizationBarrier_38_io_y_sx; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@201182.4]
  wire  OptimizationBarrier_38_io_y_sr; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@201182.4]
  wire  OptimizationBarrier_38_io_y_pw; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@201182.4]
  wire  OptimizationBarrier_38_io_y_px; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@201182.4]
  wire  OptimizationBarrier_38_io_y_pr; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@201182.4]
  wire  OptimizationBarrier_38_io_y_ppp; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@201182.4]
  wire  OptimizationBarrier_38_io_y_pal; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@201182.4]
  wire  OptimizationBarrier_38_io_y_paa; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@201182.4]
  wire  OptimizationBarrier_38_io_y_eff; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@201182.4]
  wire  OptimizationBarrier_38_io_y_c; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@201182.4]
  reg [19:0] sectored_entries_0_tag; // @[TLB.scala 162:29:freechips.rocketchip.system.DefaultRV32Config.fir@198357.4]
  reg [34:0] sectored_entries_0_data_0; // @[TLB.scala 162:29:freechips.rocketchip.system.DefaultRV32Config.fir@198357.4]
  reg [34:0] sectored_entries_0_data_1; // @[TLB.scala 162:29:freechips.rocketchip.system.DefaultRV32Config.fir@198357.4]
  reg [34:0] sectored_entries_0_data_2; // @[TLB.scala 162:29:freechips.rocketchip.system.DefaultRV32Config.fir@198357.4]
  reg [34:0] sectored_entries_0_data_3; // @[TLB.scala 162:29:freechips.rocketchip.system.DefaultRV32Config.fir@198357.4]
  reg  sectored_entries_0_valid_0; // @[TLB.scala 162:29:freechips.rocketchip.system.DefaultRV32Config.fir@198357.4]
  reg  sectored_entries_0_valid_1; // @[TLB.scala 162:29:freechips.rocketchip.system.DefaultRV32Config.fir@198357.4]
  reg  sectored_entries_0_valid_2; // @[TLB.scala 162:29:freechips.rocketchip.system.DefaultRV32Config.fir@198357.4]
  reg  sectored_entries_0_valid_3; // @[TLB.scala 162:29:freechips.rocketchip.system.DefaultRV32Config.fir@198357.4]
  reg [19:0] sectored_entries_1_tag; // @[TLB.scala 162:29:freechips.rocketchip.system.DefaultRV32Config.fir@198357.4]
  reg [34:0] sectored_entries_1_data_0; // @[TLB.scala 162:29:freechips.rocketchip.system.DefaultRV32Config.fir@198357.4]
  reg [34:0] sectored_entries_1_data_1; // @[TLB.scala 162:29:freechips.rocketchip.system.DefaultRV32Config.fir@198357.4]
  reg [34:0] sectored_entries_1_data_2; // @[TLB.scala 162:29:freechips.rocketchip.system.DefaultRV32Config.fir@198357.4]
  reg [34:0] sectored_entries_1_data_3; // @[TLB.scala 162:29:freechips.rocketchip.system.DefaultRV32Config.fir@198357.4]
  reg  sectored_entries_1_valid_0; // @[TLB.scala 162:29:freechips.rocketchip.system.DefaultRV32Config.fir@198357.4]
  reg  sectored_entries_1_valid_1; // @[TLB.scala 162:29:freechips.rocketchip.system.DefaultRV32Config.fir@198357.4]
  reg  sectored_entries_1_valid_2; // @[TLB.scala 162:29:freechips.rocketchip.system.DefaultRV32Config.fir@198357.4]
  reg  sectored_entries_1_valid_3; // @[TLB.scala 162:29:freechips.rocketchip.system.DefaultRV32Config.fir@198357.4]
  reg [19:0] sectored_entries_2_tag; // @[TLB.scala 162:29:freechips.rocketchip.system.DefaultRV32Config.fir@198357.4]
  reg [34:0] sectored_entries_2_data_0; // @[TLB.scala 162:29:freechips.rocketchip.system.DefaultRV32Config.fir@198357.4]
  reg [34:0] sectored_entries_2_data_1; // @[TLB.scala 162:29:freechips.rocketchip.system.DefaultRV32Config.fir@198357.4]
  reg [34:0] sectored_entries_2_data_2; // @[TLB.scala 162:29:freechips.rocketchip.system.DefaultRV32Config.fir@198357.4]
  reg [34:0] sectored_entries_2_data_3; // @[TLB.scala 162:29:freechips.rocketchip.system.DefaultRV32Config.fir@198357.4]
  reg  sectored_entries_2_valid_0; // @[TLB.scala 162:29:freechips.rocketchip.system.DefaultRV32Config.fir@198357.4]
  reg  sectored_entries_2_valid_1; // @[TLB.scala 162:29:freechips.rocketchip.system.DefaultRV32Config.fir@198357.4]
  reg  sectored_entries_2_valid_2; // @[TLB.scala 162:29:freechips.rocketchip.system.DefaultRV32Config.fir@198357.4]
  reg  sectored_entries_2_valid_3; // @[TLB.scala 162:29:freechips.rocketchip.system.DefaultRV32Config.fir@198357.4]
  reg [19:0] sectored_entries_3_tag; // @[TLB.scala 162:29:freechips.rocketchip.system.DefaultRV32Config.fir@198357.4]
  reg [34:0] sectored_entries_3_data_0; // @[TLB.scala 162:29:freechips.rocketchip.system.DefaultRV32Config.fir@198357.4]
  reg [34:0] sectored_entries_3_data_1; // @[TLB.scala 162:29:freechips.rocketchip.system.DefaultRV32Config.fir@198357.4]
  reg [34:0] sectored_entries_3_data_2; // @[TLB.scala 162:29:freechips.rocketchip.system.DefaultRV32Config.fir@198357.4]
  reg [34:0] sectored_entries_3_data_3; // @[TLB.scala 162:29:freechips.rocketchip.system.DefaultRV32Config.fir@198357.4]
  reg  sectored_entries_3_valid_0; // @[TLB.scala 162:29:freechips.rocketchip.system.DefaultRV32Config.fir@198357.4]
  reg  sectored_entries_3_valid_1; // @[TLB.scala 162:29:freechips.rocketchip.system.DefaultRV32Config.fir@198357.4]
  reg  sectored_entries_3_valid_2; // @[TLB.scala 162:29:freechips.rocketchip.system.DefaultRV32Config.fir@198357.4]
  reg  sectored_entries_3_valid_3; // @[TLB.scala 162:29:freechips.rocketchip.system.DefaultRV32Config.fir@198357.4]
  reg [19:0] sectored_entries_4_tag; // @[TLB.scala 162:29:freechips.rocketchip.system.DefaultRV32Config.fir@198357.4]
  reg [34:0] sectored_entries_4_data_0; // @[TLB.scala 162:29:freechips.rocketchip.system.DefaultRV32Config.fir@198357.4]
  reg [34:0] sectored_entries_4_data_1; // @[TLB.scala 162:29:freechips.rocketchip.system.DefaultRV32Config.fir@198357.4]
  reg [34:0] sectored_entries_4_data_2; // @[TLB.scala 162:29:freechips.rocketchip.system.DefaultRV32Config.fir@198357.4]
  reg [34:0] sectored_entries_4_data_3; // @[TLB.scala 162:29:freechips.rocketchip.system.DefaultRV32Config.fir@198357.4]
  reg  sectored_entries_4_valid_0; // @[TLB.scala 162:29:freechips.rocketchip.system.DefaultRV32Config.fir@198357.4]
  reg  sectored_entries_4_valid_1; // @[TLB.scala 162:29:freechips.rocketchip.system.DefaultRV32Config.fir@198357.4]
  reg  sectored_entries_4_valid_2; // @[TLB.scala 162:29:freechips.rocketchip.system.DefaultRV32Config.fir@198357.4]
  reg  sectored_entries_4_valid_3; // @[TLB.scala 162:29:freechips.rocketchip.system.DefaultRV32Config.fir@198357.4]
  reg [19:0] sectored_entries_5_tag; // @[TLB.scala 162:29:freechips.rocketchip.system.DefaultRV32Config.fir@198357.4]
  reg [34:0] sectored_entries_5_data_0; // @[TLB.scala 162:29:freechips.rocketchip.system.DefaultRV32Config.fir@198357.4]
  reg [34:0] sectored_entries_5_data_1; // @[TLB.scala 162:29:freechips.rocketchip.system.DefaultRV32Config.fir@198357.4]
  reg [34:0] sectored_entries_5_data_2; // @[TLB.scala 162:29:freechips.rocketchip.system.DefaultRV32Config.fir@198357.4]
  reg [34:0] sectored_entries_5_data_3; // @[TLB.scala 162:29:freechips.rocketchip.system.DefaultRV32Config.fir@198357.4]
  reg  sectored_entries_5_valid_0; // @[TLB.scala 162:29:freechips.rocketchip.system.DefaultRV32Config.fir@198357.4]
  reg  sectored_entries_5_valid_1; // @[TLB.scala 162:29:freechips.rocketchip.system.DefaultRV32Config.fir@198357.4]
  reg  sectored_entries_5_valid_2; // @[TLB.scala 162:29:freechips.rocketchip.system.DefaultRV32Config.fir@198357.4]
  reg  sectored_entries_5_valid_3; // @[TLB.scala 162:29:freechips.rocketchip.system.DefaultRV32Config.fir@198357.4]
  reg [19:0] sectored_entries_6_tag; // @[TLB.scala 162:29:freechips.rocketchip.system.DefaultRV32Config.fir@198357.4]
  reg [34:0] sectored_entries_6_data_0; // @[TLB.scala 162:29:freechips.rocketchip.system.DefaultRV32Config.fir@198357.4]
  reg [34:0] sectored_entries_6_data_1; // @[TLB.scala 162:29:freechips.rocketchip.system.DefaultRV32Config.fir@198357.4]
  reg [34:0] sectored_entries_6_data_2; // @[TLB.scala 162:29:freechips.rocketchip.system.DefaultRV32Config.fir@198357.4]
  reg [34:0] sectored_entries_6_data_3; // @[TLB.scala 162:29:freechips.rocketchip.system.DefaultRV32Config.fir@198357.4]
  reg  sectored_entries_6_valid_0; // @[TLB.scala 162:29:freechips.rocketchip.system.DefaultRV32Config.fir@198357.4]
  reg  sectored_entries_6_valid_1; // @[TLB.scala 162:29:freechips.rocketchip.system.DefaultRV32Config.fir@198357.4]
  reg  sectored_entries_6_valid_2; // @[TLB.scala 162:29:freechips.rocketchip.system.DefaultRV32Config.fir@198357.4]
  reg  sectored_entries_6_valid_3; // @[TLB.scala 162:29:freechips.rocketchip.system.DefaultRV32Config.fir@198357.4]
  reg [19:0] sectored_entries_7_tag; // @[TLB.scala 162:29:freechips.rocketchip.system.DefaultRV32Config.fir@198357.4]
  reg [34:0] sectored_entries_7_data_0; // @[TLB.scala 162:29:freechips.rocketchip.system.DefaultRV32Config.fir@198357.4]
  reg [34:0] sectored_entries_7_data_1; // @[TLB.scala 162:29:freechips.rocketchip.system.DefaultRV32Config.fir@198357.4]
  reg [34:0] sectored_entries_7_data_2; // @[TLB.scala 162:29:freechips.rocketchip.system.DefaultRV32Config.fir@198357.4]
  reg [34:0] sectored_entries_7_data_3; // @[TLB.scala 162:29:freechips.rocketchip.system.DefaultRV32Config.fir@198357.4]
  reg  sectored_entries_7_valid_0; // @[TLB.scala 162:29:freechips.rocketchip.system.DefaultRV32Config.fir@198357.4]
  reg  sectored_entries_7_valid_1; // @[TLB.scala 162:29:freechips.rocketchip.system.DefaultRV32Config.fir@198357.4]
  reg  sectored_entries_7_valid_2; // @[TLB.scala 162:29:freechips.rocketchip.system.DefaultRV32Config.fir@198357.4]
  reg  sectored_entries_7_valid_3; // @[TLB.scala 162:29:freechips.rocketchip.system.DefaultRV32Config.fir@198357.4]
  reg [19:0] superpage_entries_0_tag; // @[TLB.scala 163:30:freechips.rocketchip.system.DefaultRV32Config.fir@198358.4]
  reg [34:0] superpage_entries_0_data_0; // @[TLB.scala 163:30:freechips.rocketchip.system.DefaultRV32Config.fir@198358.4]
  reg  superpage_entries_0_valid_0; // @[TLB.scala 163:30:freechips.rocketchip.system.DefaultRV32Config.fir@198358.4]
  reg [19:0] superpage_entries_1_tag; // @[TLB.scala 163:30:freechips.rocketchip.system.DefaultRV32Config.fir@198358.4]
  reg [34:0] superpage_entries_1_data_0; // @[TLB.scala 163:30:freechips.rocketchip.system.DefaultRV32Config.fir@198358.4]
  reg  superpage_entries_1_valid_0; // @[TLB.scala 163:30:freechips.rocketchip.system.DefaultRV32Config.fir@198358.4]
  reg [19:0] superpage_entries_2_tag; // @[TLB.scala 163:30:freechips.rocketchip.system.DefaultRV32Config.fir@198358.4]
  reg [34:0] superpage_entries_2_data_0; // @[TLB.scala 163:30:freechips.rocketchip.system.DefaultRV32Config.fir@198358.4]
  reg  superpage_entries_2_valid_0; // @[TLB.scala 163:30:freechips.rocketchip.system.DefaultRV32Config.fir@198358.4]
  reg [19:0] superpage_entries_3_tag; // @[TLB.scala 163:30:freechips.rocketchip.system.DefaultRV32Config.fir@198358.4]
  reg [34:0] superpage_entries_3_data_0; // @[TLB.scala 163:30:freechips.rocketchip.system.DefaultRV32Config.fir@198358.4]
  reg  superpage_entries_3_valid_0; // @[TLB.scala 163:30:freechips.rocketchip.system.DefaultRV32Config.fir@198358.4]
  reg  special_entry_level; // @[TLB.scala 164:56:freechips.rocketchip.system.DefaultRV32Config.fir@198359.4]
  reg [19:0] special_entry_tag; // @[TLB.scala 164:56:freechips.rocketchip.system.DefaultRV32Config.fir@198359.4]
  reg [34:0] special_entry_data_0; // @[TLB.scala 164:56:freechips.rocketchip.system.DefaultRV32Config.fir@198359.4]
  reg  special_entry_valid_0; // @[TLB.scala 164:56:freechips.rocketchip.system.DefaultRV32Config.fir@198359.4]
  reg [1:0] state; // @[TLB.scala 169:18:freechips.rocketchip.system.DefaultRV32Config.fir@198360.4]
  reg [19:0] r_refill_tag; // @[TLB.scala 170:25:freechips.rocketchip.system.DefaultRV32Config.fir@198361.4]
  reg [1:0] r_superpage_repl_addr; // @[TLB.scala 171:34:freechips.rocketchip.system.DefaultRV32Config.fir@198362.4]
  reg [2:0] r_sectored_repl_addr; // @[TLB.scala 172:33:freechips.rocketchip.system.DefaultRV32Config.fir@198363.4]
  reg [2:0] r_sectored_hit_addr; // @[TLB.scala 173:32:freechips.rocketchip.system.DefaultRV32Config.fir@198364.4]
  reg  r_sectored_hit; // @[TLB.scala 174:27:freechips.rocketchip.system.DefaultRV32Config.fir@198365.4]
  wire  priv_s; // @[TLB.scala 177:20:freechips.rocketchip.system.DefaultRV32Config.fir@198366.4]
  wire  priv_uses_vm; // @[TLB.scala 178:27:freechips.rocketchip.system.DefaultRV32Config.fir@198367.4]
  wire  vm_enabled; // @[TLB.scala 179:83:freechips.rocketchip.system.DefaultRV32Config.fir@198370.4]
  wire [19:0] vpn; // @[TLB.scala 182:30:freechips.rocketchip.system.DefaultRV32Config.fir@198373.4]
  wire [19:0] refill_ppn; // @[TLB.scala 183:44:freechips.rocketchip.system.DefaultRV32Config.fir@198374.4]
  wire  _T_4; // @[package.scala 15:47:freechips.rocketchip.system.DefaultRV32Config.fir@198376.4]
  wire  _T_5; // @[package.scala 15:47:freechips.rocketchip.system.DefaultRV32Config.fir@198377.4]
  wire  invalidate_refill; // @[package.scala 64:59:freechips.rocketchip.system.DefaultRV32Config.fir@198378.4]
  wire  _T_26; // @[TLB.scala 108:28:freechips.rocketchip.system.DefaultRV32Config.fir@198423.4]
  wire [19:0] _T_28; // @[TLB.scala 109:28:freechips.rocketchip.system.DefaultRV32Config.fir@198425.4]
  wire [19:0] _T_29; // @[TLB.scala 109:47:freechips.rocketchip.system.DefaultRV32Config.fir@198426.4]
  wire [19:0] _T_31; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@198428.4]
  wire [19:0] _T_33; // @[TLB.scala 187:20:freechips.rocketchip.system.DefaultRV32Config.fir@198430.4]
  wire [19:0] mpu_ppn; // @[TLB.scala 186:20:freechips.rocketchip.system.DefaultRV32Config.fir@198431.4]
  wire [31:0] mpu_physaddr; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@198433.4]
  wire [2:0] _T_37; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@198436.4]
  wire [2:0] mpu_priv; // @[TLB.scala 189:27:freechips.rocketchip.system.DefaultRV32Config.fir@198437.4]
  wire [31:0] _T_38; // @[Parameters.scala 137:31:freechips.rocketchip.system.DefaultRV32Config.fir@198453.4]
  wire [32:0] _T_39; // @[Parameters.scala 137:49:freechips.rocketchip.system.DefaultRV32Config.fir@198454.4]
  wire [32:0] _T_41; // @[Parameters.scala 137:52:freechips.rocketchip.system.DefaultRV32Config.fir@198456.4]
  wire  _T_42; // @[Parameters.scala 137:67:freechips.rocketchip.system.DefaultRV32Config.fir@198457.4]
  wire [31:0] _T_43; // @[Parameters.scala 137:31:freechips.rocketchip.system.DefaultRV32Config.fir@198458.4]
  wire [32:0] _T_44; // @[Parameters.scala 137:49:freechips.rocketchip.system.DefaultRV32Config.fir@198459.4]
  wire [32:0] _T_46; // @[Parameters.scala 137:52:freechips.rocketchip.system.DefaultRV32Config.fir@198461.4]
  wire  _T_47; // @[Parameters.scala 137:67:freechips.rocketchip.system.DefaultRV32Config.fir@198462.4]
  wire [31:0] _T_48; // @[Parameters.scala 137:31:freechips.rocketchip.system.DefaultRV32Config.fir@198463.4]
  wire [32:0] _T_49; // @[Parameters.scala 137:49:freechips.rocketchip.system.DefaultRV32Config.fir@198464.4]
  wire [32:0] _T_51; // @[Parameters.scala 137:52:freechips.rocketchip.system.DefaultRV32Config.fir@198466.4]
  wire  _T_52; // @[Parameters.scala 137:67:freechips.rocketchip.system.DefaultRV32Config.fir@198467.4]
  wire [32:0] _T_54; // @[Parameters.scala 137:49:freechips.rocketchip.system.DefaultRV32Config.fir@198469.4]
  wire [32:0] _T_56; // @[Parameters.scala 137:52:freechips.rocketchip.system.DefaultRV32Config.fir@198471.4]
  wire  _T_57; // @[Parameters.scala 137:67:freechips.rocketchip.system.DefaultRV32Config.fir@198472.4]
  wire [31:0] _T_58; // @[Parameters.scala 137:31:freechips.rocketchip.system.DefaultRV32Config.fir@198473.4]
  wire [32:0] _T_59; // @[Parameters.scala 137:49:freechips.rocketchip.system.DefaultRV32Config.fir@198474.4]
  wire [32:0] _T_61; // @[Parameters.scala 137:52:freechips.rocketchip.system.DefaultRV32Config.fir@198476.4]
  wire  _T_62; // @[Parameters.scala 137:67:freechips.rocketchip.system.DefaultRV32Config.fir@198477.4]
  wire [31:0] _T_63; // @[Parameters.scala 137:31:freechips.rocketchip.system.DefaultRV32Config.fir@198478.4]
  wire [32:0] _T_64; // @[Parameters.scala 137:49:freechips.rocketchip.system.DefaultRV32Config.fir@198479.4]
  wire [32:0] _T_66; // @[Parameters.scala 137:52:freechips.rocketchip.system.DefaultRV32Config.fir@198481.4]
  wire  _T_67; // @[Parameters.scala 137:67:freechips.rocketchip.system.DefaultRV32Config.fir@198482.4]
  wire [31:0] _T_68; // @[Parameters.scala 137:31:freechips.rocketchip.system.DefaultRV32Config.fir@198483.4]
  wire [32:0] _T_69; // @[Parameters.scala 137:49:freechips.rocketchip.system.DefaultRV32Config.fir@198484.4]
  wire [32:0] _T_71; // @[Parameters.scala 137:52:freechips.rocketchip.system.DefaultRV32Config.fir@198486.4]
  wire  _T_72; // @[Parameters.scala 137:67:freechips.rocketchip.system.DefaultRV32Config.fir@198487.4]
  wire  _T_74; // @[TLB.scala 195:67:freechips.rocketchip.system.DefaultRV32Config.fir@198497.4]
  wire  _T_75; // @[TLB.scala 195:67:freechips.rocketchip.system.DefaultRV32Config.fir@198498.4]
  wire  _T_76; // @[TLB.scala 195:67:freechips.rocketchip.system.DefaultRV32Config.fir@198499.4]
  wire  _T_77; // @[TLB.scala 195:67:freechips.rocketchip.system.DefaultRV32Config.fir@198500.4]
  wire  _T_78; // @[TLB.scala 195:67:freechips.rocketchip.system.DefaultRV32Config.fir@198501.4]
  wire  legal_address; // @[TLB.scala 195:67:freechips.rocketchip.system.DefaultRV32Config.fir@198502.4]
  wire [32:0] _T_87; // @[Parameters.scala 137:52:freechips.rocketchip.system.DefaultRV32Config.fir@198511.4]
  wire  _T_88; // @[Parameters.scala 137:67:freechips.rocketchip.system.DefaultRV32Config.fir@198512.4]
  wire  cacheable; // @[TLB.scala 197:19:freechips.rocketchip.system.DefaultRV32Config.fir@198518.4]
  wire [31:0] _T_148; // @[Parameters.scala 137:31:freechips.rocketchip.system.DefaultRV32Config.fir@198575.4]
  wire [32:0] _T_149; // @[Parameters.scala 137:49:freechips.rocketchip.system.DefaultRV32Config.fir@198576.4]
  wire [32:0] _T_151; // @[Parameters.scala 137:52:freechips.rocketchip.system.DefaultRV32Config.fir@198578.4]
  wire  _T_152; // @[Parameters.scala 137:67:freechips.rocketchip.system.DefaultRV32Config.fir@198579.4]
  wire [32:0] _T_165; // @[Parameters.scala 137:52:freechips.rocketchip.system.DefaultRV32Config.fir@198592.4]
  wire  _T_166; // @[Parameters.scala 137:67:freechips.rocketchip.system.DefaultRV32Config.fir@198593.4]
  wire  _T_173; // @[TLBPermissions.scala 82:66:freechips.rocketchip.system.DefaultRV32Config.fir@198600.4]
  wire  _T_186; // @[TLB.scala 200:39:freechips.rocketchip.system.DefaultRV32Config.fir@198613.4]
  wire  deny_access_to_debug; // @[TLB.scala 200:48:freechips.rocketchip.system.DefaultRV32Config.fir@198619.4]
  wire  _T_198; // @[TLB.scala 201:44:freechips.rocketchip.system.DefaultRV32Config.fir@198626.4]
  wire  _T_199; // @[TLB.scala 201:41:freechips.rocketchip.system.DefaultRV32Config.fir@198627.4]
  wire  prot_r; // @[TLB.scala 201:66:freechips.rocketchip.system.DefaultRV32Config.fir@198628.4]
  wire [31:0] _T_210; // @[Parameters.scala 137:31:freechips.rocketchip.system.DefaultRV32Config.fir@198639.4]
  wire [32:0] _T_211; // @[Parameters.scala 137:49:freechips.rocketchip.system.DefaultRV32Config.fir@198640.4]
  wire [32:0] _T_213; // @[Parameters.scala 137:52:freechips.rocketchip.system.DefaultRV32Config.fir@198642.4]
  wire  _T_214; // @[Parameters.scala 137:67:freechips.rocketchip.system.DefaultRV32Config.fir@198643.4]
  wire [32:0] _T_218; // @[Parameters.scala 137:52:freechips.rocketchip.system.DefaultRV32Config.fir@198647.4]
  wire  _T_219; // @[Parameters.scala 137:67:freechips.rocketchip.system.DefaultRV32Config.fir@198648.4]
  wire  _T_221; // @[Parameters.scala 528:89:freechips.rocketchip.system.DefaultRV32Config.fir@198650.4]
  wire  _T_222; // @[Parameters.scala 528:89:freechips.rocketchip.system.DefaultRV32Config.fir@198651.4]
  wire  _T_232; // @[TLB.scala 197:19:freechips.rocketchip.system.DefaultRV32Config.fir@198662.4]
  wire  _T_234; // @[TLB.scala 202:45:freechips.rocketchip.system.DefaultRV32Config.fir@198664.4]
  wire  prot_w; // @[TLB.scala 202:70:freechips.rocketchip.system.DefaultRV32Config.fir@198665.4]
  wire  prot_al; // @[TLB.scala 197:19:freechips.rocketchip.system.DefaultRV32Config.fir@198733.4]
  wire [32:0] _T_334; // @[Parameters.scala 137:52:freechips.rocketchip.system.DefaultRV32Config.fir@198771.4]
  wire  _T_335; // @[Parameters.scala 137:67:freechips.rocketchip.system.DefaultRV32Config.fir@198772.4]
  wire  _T_346; // @[Parameters.scala 528:89:freechips.rocketchip.system.DefaultRV32Config.fir@198783.4]
  wire  _T_347; // @[Parameters.scala 528:89:freechips.rocketchip.system.DefaultRV32Config.fir@198784.4]
  wire  _T_363; // @[TLB.scala 197:19:freechips.rocketchip.system.DefaultRV32Config.fir@198801.4]
  wire  _T_365; // @[TLB.scala 206:40:freechips.rocketchip.system.DefaultRV32Config.fir@198803.4]
  wire  prot_x; // @[TLB.scala 206:65:freechips.rocketchip.system.DefaultRV32Config.fir@198804.4]
  wire [32:0] _T_386; // @[Parameters.scala 137:52:freechips.rocketchip.system.DefaultRV32Config.fir@198825.4]
  wire  _T_387; // @[Parameters.scala 137:67:freechips.rocketchip.system.DefaultRV32Config.fir@198826.4]
  wire [32:0] _T_391; // @[Parameters.scala 137:52:freechips.rocketchip.system.DefaultRV32Config.fir@198830.4]
  wire  _T_392; // @[Parameters.scala 137:67:freechips.rocketchip.system.DefaultRV32Config.fir@198831.4]
  wire  _T_403; // @[Parameters.scala 528:89:freechips.rocketchip.system.DefaultRV32Config.fir@198842.4]
  wire  _T_404; // @[Parameters.scala 528:89:freechips.rocketchip.system.DefaultRV32Config.fir@198843.4]
  wire  _T_405; // @[Parameters.scala 528:89:freechips.rocketchip.system.DefaultRV32Config.fir@198844.4]
  wire  prot_eff; // @[TLB.scala 197:19:freechips.rocketchip.system.DefaultRV32Config.fir@198850.4]
  wire  _T_410; // @[package.scala 64:59:freechips.rocketchip.system.DefaultRV32Config.fir@198851.4]
  wire  _T_411; // @[package.scala 64:59:freechips.rocketchip.system.DefaultRV32Config.fir@198852.4]
  wire  _T_412; // @[package.scala 64:59:freechips.rocketchip.system.DefaultRV32Config.fir@198853.4]
  wire [19:0] _T_413; // @[TLB.scala 88:41:freechips.rocketchip.system.DefaultRV32Config.fir@198854.4]
  wire  _T_415; // @[TLB.scala 88:66:freechips.rocketchip.system.DefaultRV32Config.fir@198856.4]
  wire  sector_hits_0; // @[TLB.scala 87:40:freechips.rocketchip.system.DefaultRV32Config.fir@198857.4]
  wire  _T_416; // @[package.scala 64:59:freechips.rocketchip.system.DefaultRV32Config.fir@198858.4]
  wire  _T_417; // @[package.scala 64:59:freechips.rocketchip.system.DefaultRV32Config.fir@198859.4]
  wire  _T_418; // @[package.scala 64:59:freechips.rocketchip.system.DefaultRV32Config.fir@198860.4]
  wire [19:0] _T_419; // @[TLB.scala 88:41:freechips.rocketchip.system.DefaultRV32Config.fir@198861.4]
  wire  _T_421; // @[TLB.scala 88:66:freechips.rocketchip.system.DefaultRV32Config.fir@198863.4]
  wire  sector_hits_1; // @[TLB.scala 87:40:freechips.rocketchip.system.DefaultRV32Config.fir@198864.4]
  wire  _T_422; // @[package.scala 64:59:freechips.rocketchip.system.DefaultRV32Config.fir@198865.4]
  wire  _T_423; // @[package.scala 64:59:freechips.rocketchip.system.DefaultRV32Config.fir@198866.4]
  wire  _T_424; // @[package.scala 64:59:freechips.rocketchip.system.DefaultRV32Config.fir@198867.4]
  wire [19:0] _T_425; // @[TLB.scala 88:41:freechips.rocketchip.system.DefaultRV32Config.fir@198868.4]
  wire  _T_427; // @[TLB.scala 88:66:freechips.rocketchip.system.DefaultRV32Config.fir@198870.4]
  wire  sector_hits_2; // @[TLB.scala 87:40:freechips.rocketchip.system.DefaultRV32Config.fir@198871.4]
  wire  _T_428; // @[package.scala 64:59:freechips.rocketchip.system.DefaultRV32Config.fir@198872.4]
  wire  _T_429; // @[package.scala 64:59:freechips.rocketchip.system.DefaultRV32Config.fir@198873.4]
  wire  _T_430; // @[package.scala 64:59:freechips.rocketchip.system.DefaultRV32Config.fir@198874.4]
  wire [19:0] _T_431; // @[TLB.scala 88:41:freechips.rocketchip.system.DefaultRV32Config.fir@198875.4]
  wire  _T_433; // @[TLB.scala 88:66:freechips.rocketchip.system.DefaultRV32Config.fir@198877.4]
  wire  sector_hits_3; // @[TLB.scala 87:40:freechips.rocketchip.system.DefaultRV32Config.fir@198878.4]
  wire  _T_434; // @[package.scala 64:59:freechips.rocketchip.system.DefaultRV32Config.fir@198879.4]
  wire  _T_435; // @[package.scala 64:59:freechips.rocketchip.system.DefaultRV32Config.fir@198880.4]
  wire  _T_436; // @[package.scala 64:59:freechips.rocketchip.system.DefaultRV32Config.fir@198881.4]
  wire [19:0] _T_437; // @[TLB.scala 88:41:freechips.rocketchip.system.DefaultRV32Config.fir@198882.4]
  wire  _T_439; // @[TLB.scala 88:66:freechips.rocketchip.system.DefaultRV32Config.fir@198884.4]
  wire  sector_hits_4; // @[TLB.scala 87:40:freechips.rocketchip.system.DefaultRV32Config.fir@198885.4]
  wire  _T_440; // @[package.scala 64:59:freechips.rocketchip.system.DefaultRV32Config.fir@198886.4]
  wire  _T_441; // @[package.scala 64:59:freechips.rocketchip.system.DefaultRV32Config.fir@198887.4]
  wire  _T_442; // @[package.scala 64:59:freechips.rocketchip.system.DefaultRV32Config.fir@198888.4]
  wire [19:0] _T_443; // @[TLB.scala 88:41:freechips.rocketchip.system.DefaultRV32Config.fir@198889.4]
  wire  _T_445; // @[TLB.scala 88:66:freechips.rocketchip.system.DefaultRV32Config.fir@198891.4]
  wire  sector_hits_5; // @[TLB.scala 87:40:freechips.rocketchip.system.DefaultRV32Config.fir@198892.4]
  wire  _T_446; // @[package.scala 64:59:freechips.rocketchip.system.DefaultRV32Config.fir@198893.4]
  wire  _T_447; // @[package.scala 64:59:freechips.rocketchip.system.DefaultRV32Config.fir@198894.4]
  wire  _T_448; // @[package.scala 64:59:freechips.rocketchip.system.DefaultRV32Config.fir@198895.4]
  wire [19:0] _T_449; // @[TLB.scala 88:41:freechips.rocketchip.system.DefaultRV32Config.fir@198896.4]
  wire  _T_451; // @[TLB.scala 88:66:freechips.rocketchip.system.DefaultRV32Config.fir@198898.4]
  wire  sector_hits_6; // @[TLB.scala 87:40:freechips.rocketchip.system.DefaultRV32Config.fir@198899.4]
  wire  _T_452; // @[package.scala 64:59:freechips.rocketchip.system.DefaultRV32Config.fir@198900.4]
  wire  _T_453; // @[package.scala 64:59:freechips.rocketchip.system.DefaultRV32Config.fir@198901.4]
  wire  _T_454; // @[package.scala 64:59:freechips.rocketchip.system.DefaultRV32Config.fir@198902.4]
  wire [19:0] _T_455; // @[TLB.scala 88:41:freechips.rocketchip.system.DefaultRV32Config.fir@198903.4]
  wire  _T_457; // @[TLB.scala 88:66:freechips.rocketchip.system.DefaultRV32Config.fir@198905.4]
  wire  sector_hits_7; // @[TLB.scala 87:40:freechips.rocketchip.system.DefaultRV32Config.fir@198906.4]
  wire  _T_462; // @[TLB.scala 95:77:freechips.rocketchip.system.DefaultRV32Config.fir@198911.4]
  wire  superpage_hits_0; // @[TLB.scala 95:29:freechips.rocketchip.system.DefaultRV32Config.fir@198913.4]
  wire  _T_475; // @[TLB.scala 95:77:freechips.rocketchip.system.DefaultRV32Config.fir@198925.4]
  wire  superpage_hits_1; // @[TLB.scala 95:29:freechips.rocketchip.system.DefaultRV32Config.fir@198927.4]
  wire  _T_488; // @[TLB.scala 95:77:freechips.rocketchip.system.DefaultRV32Config.fir@198939.4]
  wire  superpage_hits_2; // @[TLB.scala 95:29:freechips.rocketchip.system.DefaultRV32Config.fir@198941.4]
  wire  _T_501; // @[TLB.scala 95:77:freechips.rocketchip.system.DefaultRV32Config.fir@198953.4]
  wire  superpage_hits_3; // @[TLB.scala 95:29:freechips.rocketchip.system.DefaultRV32Config.fir@198955.4]
  wire  _GEN_1; // @[TLB.scala 100:18:freechips.rocketchip.system.DefaultRV32Config.fir@198967.4]
  wire  _GEN_2; // @[TLB.scala 100:18:freechips.rocketchip.system.DefaultRV32Config.fir@198967.4]
  wire  _GEN_3; // @[TLB.scala 100:18:freechips.rocketchip.system.DefaultRV32Config.fir@198967.4]
  wire  _T_514; // @[TLB.scala 100:18:freechips.rocketchip.system.DefaultRV32Config.fir@198967.4]
  wire  hitsVec_0; // @[TLB.scala 211:44:freechips.rocketchip.system.DefaultRV32Config.fir@198968.4]
  wire  _GEN_5; // @[TLB.scala 100:18:freechips.rocketchip.system.DefaultRV32Config.fir@198973.4]
  wire  _GEN_6; // @[TLB.scala 100:18:freechips.rocketchip.system.DefaultRV32Config.fir@198973.4]
  wire  _GEN_7; // @[TLB.scala 100:18:freechips.rocketchip.system.DefaultRV32Config.fir@198973.4]
  wire  _T_519; // @[TLB.scala 100:18:freechips.rocketchip.system.DefaultRV32Config.fir@198973.4]
  wire  hitsVec_1; // @[TLB.scala 211:44:freechips.rocketchip.system.DefaultRV32Config.fir@198974.4]
  wire  _GEN_9; // @[TLB.scala 100:18:freechips.rocketchip.system.DefaultRV32Config.fir@198979.4]
  wire  _GEN_10; // @[TLB.scala 100:18:freechips.rocketchip.system.DefaultRV32Config.fir@198979.4]
  wire  _GEN_11; // @[TLB.scala 100:18:freechips.rocketchip.system.DefaultRV32Config.fir@198979.4]
  wire  _T_524; // @[TLB.scala 100:18:freechips.rocketchip.system.DefaultRV32Config.fir@198979.4]
  wire  hitsVec_2; // @[TLB.scala 211:44:freechips.rocketchip.system.DefaultRV32Config.fir@198980.4]
  wire  _GEN_13; // @[TLB.scala 100:18:freechips.rocketchip.system.DefaultRV32Config.fir@198985.4]
  wire  _GEN_14; // @[TLB.scala 100:18:freechips.rocketchip.system.DefaultRV32Config.fir@198985.4]
  wire  _GEN_15; // @[TLB.scala 100:18:freechips.rocketchip.system.DefaultRV32Config.fir@198985.4]
  wire  _T_529; // @[TLB.scala 100:18:freechips.rocketchip.system.DefaultRV32Config.fir@198985.4]
  wire  hitsVec_3; // @[TLB.scala 211:44:freechips.rocketchip.system.DefaultRV32Config.fir@198986.4]
  wire  _GEN_17; // @[TLB.scala 100:18:freechips.rocketchip.system.DefaultRV32Config.fir@198991.4]
  wire  _GEN_18; // @[TLB.scala 100:18:freechips.rocketchip.system.DefaultRV32Config.fir@198991.4]
  wire  _GEN_19; // @[TLB.scala 100:18:freechips.rocketchip.system.DefaultRV32Config.fir@198991.4]
  wire  _T_534; // @[TLB.scala 100:18:freechips.rocketchip.system.DefaultRV32Config.fir@198991.4]
  wire  hitsVec_4; // @[TLB.scala 211:44:freechips.rocketchip.system.DefaultRV32Config.fir@198992.4]
  wire  _GEN_21; // @[TLB.scala 100:18:freechips.rocketchip.system.DefaultRV32Config.fir@198997.4]
  wire  _GEN_22; // @[TLB.scala 100:18:freechips.rocketchip.system.DefaultRV32Config.fir@198997.4]
  wire  _GEN_23; // @[TLB.scala 100:18:freechips.rocketchip.system.DefaultRV32Config.fir@198997.4]
  wire  _T_539; // @[TLB.scala 100:18:freechips.rocketchip.system.DefaultRV32Config.fir@198997.4]
  wire  hitsVec_5; // @[TLB.scala 211:44:freechips.rocketchip.system.DefaultRV32Config.fir@198998.4]
  wire  _GEN_25; // @[TLB.scala 100:18:freechips.rocketchip.system.DefaultRV32Config.fir@199003.4]
  wire  _GEN_26; // @[TLB.scala 100:18:freechips.rocketchip.system.DefaultRV32Config.fir@199003.4]
  wire  _GEN_27; // @[TLB.scala 100:18:freechips.rocketchip.system.DefaultRV32Config.fir@199003.4]
  wire  _T_544; // @[TLB.scala 100:18:freechips.rocketchip.system.DefaultRV32Config.fir@199003.4]
  wire  hitsVec_6; // @[TLB.scala 211:44:freechips.rocketchip.system.DefaultRV32Config.fir@199004.4]
  wire  _GEN_29; // @[TLB.scala 100:18:freechips.rocketchip.system.DefaultRV32Config.fir@199009.4]
  wire  _GEN_30; // @[TLB.scala 100:18:freechips.rocketchip.system.DefaultRV32Config.fir@199009.4]
  wire  _GEN_31; // @[TLB.scala 100:18:freechips.rocketchip.system.DefaultRV32Config.fir@199009.4]
  wire  _T_549; // @[TLB.scala 100:18:freechips.rocketchip.system.DefaultRV32Config.fir@199009.4]
  wire  hitsVec_7; // @[TLB.scala 211:44:freechips.rocketchip.system.DefaultRV32Config.fir@199010.4]
  wire  hitsVec_8; // @[TLB.scala 211:44:freechips.rocketchip.system.DefaultRV32Config.fir@199025.4]
  wire  hitsVec_9; // @[TLB.scala 211:44:freechips.rocketchip.system.DefaultRV32Config.fir@199040.4]
  wire  hitsVec_10; // @[TLB.scala 211:44:freechips.rocketchip.system.DefaultRV32Config.fir@199055.4]
  wire  hitsVec_11; // @[TLB.scala 211:44:freechips.rocketchip.system.DefaultRV32Config.fir@199070.4]
  wire  _T_610; // @[TLB.scala 95:77:freechips.rocketchip.system.DefaultRV32Config.fir@199075.4]
  wire  _T_612; // @[TLB.scala 95:29:freechips.rocketchip.system.DefaultRV32Config.fir@199077.4]
  wire  _T_617; // @[TLB.scala 95:77:freechips.rocketchip.system.DefaultRV32Config.fir@199082.4]
  wire  _T_618; // @[TLB.scala 95:40:freechips.rocketchip.system.DefaultRV32Config.fir@199083.4]
  wire  _T_619; // @[TLB.scala 95:29:freechips.rocketchip.system.DefaultRV32Config.fir@199084.4]
  wire  hitsVec_12; // @[TLB.scala 211:44:freechips.rocketchip.system.DefaultRV32Config.fir@199085.4]
  wire [5:0] _T_624; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@199090.4]
  wire [12:0] real_hits; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@199097.4]
  wire  _T_631; // @[TLB.scala 213:18:freechips.rocketchip.system.DefaultRV32Config.fir@199098.4]
  wire [13:0] hits; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@199099.4]
  wire [34:0] _GEN_33; // @[:freechips.rocketchip.system.DefaultRV32Config.fir@199106.4]
  wire [34:0] _GEN_34; // @[:freechips.rocketchip.system.DefaultRV32Config.fir@199106.4]
  wire [34:0] _GEN_35; // @[:freechips.rocketchip.system.DefaultRV32Config.fir@199106.4]
  wire [34:0] _GEN_37; // @[:freechips.rocketchip.system.DefaultRV32Config.fir@199149.4]
  wire [34:0] _GEN_38; // @[:freechips.rocketchip.system.DefaultRV32Config.fir@199149.4]
  wire [34:0] _GEN_39; // @[:freechips.rocketchip.system.DefaultRV32Config.fir@199149.4]
  wire [34:0] _GEN_41; // @[:freechips.rocketchip.system.DefaultRV32Config.fir@199192.4]
  wire [34:0] _GEN_42; // @[:freechips.rocketchip.system.DefaultRV32Config.fir@199192.4]
  wire [34:0] _GEN_43; // @[:freechips.rocketchip.system.DefaultRV32Config.fir@199192.4]
  wire [34:0] _GEN_45; // @[:freechips.rocketchip.system.DefaultRV32Config.fir@199235.4]
  wire [34:0] _GEN_46; // @[:freechips.rocketchip.system.DefaultRV32Config.fir@199235.4]
  wire [34:0] _GEN_47; // @[:freechips.rocketchip.system.DefaultRV32Config.fir@199235.4]
  wire [34:0] _GEN_49; // @[:freechips.rocketchip.system.DefaultRV32Config.fir@199278.4]
  wire [34:0] _GEN_50; // @[:freechips.rocketchip.system.DefaultRV32Config.fir@199278.4]
  wire [34:0] _GEN_51; // @[:freechips.rocketchip.system.DefaultRV32Config.fir@199278.4]
  wire [34:0] _GEN_53; // @[:freechips.rocketchip.system.DefaultRV32Config.fir@199321.4]
  wire [34:0] _GEN_54; // @[:freechips.rocketchip.system.DefaultRV32Config.fir@199321.4]
  wire [34:0] _GEN_55; // @[:freechips.rocketchip.system.DefaultRV32Config.fir@199321.4]
  wire [34:0] _GEN_57; // @[:freechips.rocketchip.system.DefaultRV32Config.fir@199364.4]
  wire [34:0] _GEN_58; // @[:freechips.rocketchip.system.DefaultRV32Config.fir@199364.4]
  wire [34:0] _GEN_59; // @[:freechips.rocketchip.system.DefaultRV32Config.fir@199364.4]
  wire [34:0] _GEN_61; // @[:freechips.rocketchip.system.DefaultRV32Config.fir@199407.4]
  wire [34:0] _GEN_62; // @[:freechips.rocketchip.system.DefaultRV32Config.fir@199407.4]
  wire [34:0] _GEN_63; // @[:freechips.rocketchip.system.DefaultRV32Config.fir@199407.4]
  wire [19:0] _T_807; // @[TLB.scala 109:47:freechips.rocketchip.system.DefaultRV32Config.fir@199491.4]
  wire [19:0] _T_809; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@199493.4]
  wire [19:0] _T_832; // @[TLB.scala 109:47:freechips.rocketchip.system.DefaultRV32Config.fir@199540.4]
  wire [19:0] _T_834; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@199542.4]
  wire [19:0] _T_857; // @[TLB.scala 109:47:freechips.rocketchip.system.DefaultRV32Config.fir@199589.4]
  wire [19:0] _T_859; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@199591.4]
  wire [19:0] _T_882; // @[TLB.scala 109:47:freechips.rocketchip.system.DefaultRV32Config.fir@199638.4]
  wire [19:0] _T_884; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@199640.4]
  wire [19:0] _T_907; // @[TLB.scala 109:47:freechips.rocketchip.system.DefaultRV32Config.fir@199687.4]
  wire [19:0] _T_909; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@199689.4]
  wire [19:0] _T_911; // @[Mux.scala 27:72:freechips.rocketchip.system.DefaultRV32Config.fir@199691.4]
  wire [19:0] _T_912; // @[Mux.scala 27:72:freechips.rocketchip.system.DefaultRV32Config.fir@199692.4]
  wire [19:0] _T_913; // @[Mux.scala 27:72:freechips.rocketchip.system.DefaultRV32Config.fir@199693.4]
  wire [19:0] _T_914; // @[Mux.scala 27:72:freechips.rocketchip.system.DefaultRV32Config.fir@199694.4]
  wire [19:0] _T_915; // @[Mux.scala 27:72:freechips.rocketchip.system.DefaultRV32Config.fir@199695.4]
  wire [19:0] _T_916; // @[Mux.scala 27:72:freechips.rocketchip.system.DefaultRV32Config.fir@199696.4]
  wire [19:0] _T_917; // @[Mux.scala 27:72:freechips.rocketchip.system.DefaultRV32Config.fir@199697.4]
  wire [19:0] _T_918; // @[Mux.scala 27:72:freechips.rocketchip.system.DefaultRV32Config.fir@199698.4]
  wire [19:0] _T_919; // @[Mux.scala 27:72:freechips.rocketchip.system.DefaultRV32Config.fir@199699.4]
  wire [19:0] _T_920; // @[Mux.scala 27:72:freechips.rocketchip.system.DefaultRV32Config.fir@199700.4]
  wire [19:0] _T_921; // @[Mux.scala 27:72:freechips.rocketchip.system.DefaultRV32Config.fir@199701.4]
  wire [19:0] _T_922; // @[Mux.scala 27:72:freechips.rocketchip.system.DefaultRV32Config.fir@199702.4]
  wire [19:0] _T_923; // @[Mux.scala 27:72:freechips.rocketchip.system.DefaultRV32Config.fir@199703.4]
  wire [19:0] _T_924; // @[Mux.scala 27:72:freechips.rocketchip.system.DefaultRV32Config.fir@199704.4]
  wire [19:0] _T_925; // @[Mux.scala 27:72:freechips.rocketchip.system.DefaultRV32Config.fir@199705.4]
  wire [19:0] _T_926; // @[Mux.scala 27:72:freechips.rocketchip.system.DefaultRV32Config.fir@199706.4]
  wire [19:0] _T_927; // @[Mux.scala 27:72:freechips.rocketchip.system.DefaultRV32Config.fir@199707.4]
  wire [19:0] _T_928; // @[Mux.scala 27:72:freechips.rocketchip.system.DefaultRV32Config.fir@199708.4]
  wire [19:0] _T_929; // @[Mux.scala 27:72:freechips.rocketchip.system.DefaultRV32Config.fir@199709.4]
  wire [19:0] _T_930; // @[Mux.scala 27:72:freechips.rocketchip.system.DefaultRV32Config.fir@199710.4]
  wire [19:0] _T_931; // @[Mux.scala 27:72:freechips.rocketchip.system.DefaultRV32Config.fir@199711.4]
  wire [19:0] _T_932; // @[Mux.scala 27:72:freechips.rocketchip.system.DefaultRV32Config.fir@199712.4]
  wire [19:0] _T_933; // @[Mux.scala 27:72:freechips.rocketchip.system.DefaultRV32Config.fir@199713.4]
  wire [19:0] _T_934; // @[Mux.scala 27:72:freechips.rocketchip.system.DefaultRV32Config.fir@199714.4]
  wire [19:0] _T_935; // @[Mux.scala 27:72:freechips.rocketchip.system.DefaultRV32Config.fir@199715.4]
  wire [19:0] _T_936; // @[Mux.scala 27:72:freechips.rocketchip.system.DefaultRV32Config.fir@199716.4]
  wire [19:0] ppn; // @[Mux.scala 27:72:freechips.rocketchip.system.DefaultRV32Config.fir@199717.4]
  wire  _T_938; // @[TLB.scala 217:22:freechips.rocketchip.system.DefaultRV32Config.fir@199720.4]
  wire  _T_939; // @[TLB.scala 217:19:freechips.rocketchip.system.DefaultRV32Config.fir@199721.4]
  wire  _T_941; // @[TLB.scala 223:25:freechips.rocketchip.system.DefaultRV32Config.fir@199728.6]
  wire  _T_942; // @[PTW.scala 69:47:freechips.rocketchip.system.DefaultRV32Config.fir@199731.6]
  wire  _T_943; // @[PTW.scala 69:44:freechips.rocketchip.system.DefaultRV32Config.fir@199732.6]
  wire  _T_944; // @[PTW.scala 69:38:freechips.rocketchip.system.DefaultRV32Config.fir@199733.6]
  wire  _T_945; // @[PTW.scala 69:32:freechips.rocketchip.system.DefaultRV32Config.fir@199734.6]
  wire  _T_946; // @[PTW.scala 69:52:freechips.rocketchip.system.DefaultRV32Config.fir@199735.6]
  wire  _T_947; // @[PTW.scala 73:35:freechips.rocketchip.system.DefaultRV32Config.fir@199736.6]
  wire  _T_953; // @[PTW.scala 74:35:freechips.rocketchip.system.DefaultRV32Config.fir@199743.6]
  wire  _T_954; // @[PTW.scala 74:40:freechips.rocketchip.system.DefaultRV32Config.fir@199744.6]
  wire  _T_960; // @[PTW.scala 75:35:freechips.rocketchip.system.DefaultRV32Config.fir@199751.6]
  wire  _T_961; // @[TLB.scala 237:37:freechips.rocketchip.system.DefaultRV32Config.fir@199761.6]
  wire [7:0] _T_970; // @[TLB.scala 123:24:freechips.rocketchip.system.DefaultRV32Config.fir@199774.8]
  wire [34:0] _T_978; // @[TLB.scala 123:24:freechips.rocketchip.system.DefaultRV32Config.fir@199782.8]
  wire  _T_979; // @[TLB.scala 239:40:freechips.rocketchip.system.DefaultRV32Config.fir@199786.8]
  wire  _T_980; // @[TLB.scala 240:82:freechips.rocketchip.system.DefaultRV32Config.fir@199788.10]
  wire  _GEN_66; // @[TLB.scala 240:89:freechips.rocketchip.system.DefaultRV32Config.fir@199789.10]
  wire  _T_996; // @[TLB.scala 240:82:freechips.rocketchip.system.DefaultRV32Config.fir@199810.10]
  wire  _GEN_70; // @[TLB.scala 240:89:freechips.rocketchip.system.DefaultRV32Config.fir@199811.10]
  wire  _T_1012; // @[TLB.scala 240:82:freechips.rocketchip.system.DefaultRV32Config.fir@199832.10]
  wire  _GEN_74; // @[TLB.scala 240:89:freechips.rocketchip.system.DefaultRV32Config.fir@199833.10]
  wire  _T_1028; // @[TLB.scala 240:82:freechips.rocketchip.system.DefaultRV32Config.fir@199854.10]
  wire  _GEN_78; // @[TLB.scala 240:89:freechips.rocketchip.system.DefaultRV32Config.fir@199855.10]
  wire [2:0] _T_1044; // @[TLB.scala 244:22:freechips.rocketchip.system.DefaultRV32Config.fir@199878.10]
  wire  _T_1045; // @[TLB.scala 245:65:freechips.rocketchip.system.DefaultRV32Config.fir@199879.10]
  wire  _T_1046; // @[TLB.scala 246:15:freechips.rocketchip.system.DefaultRV32Config.fir@199881.12]
  wire  _GEN_80; // @[TLB.scala 246:32:freechips.rocketchip.system.DefaultRV32Config.fir@199882.12]
  wire  _GEN_81; // @[TLB.scala 246:32:freechips.rocketchip.system.DefaultRV32Config.fir@199882.12]
  wire  _GEN_82; // @[TLB.scala 246:32:freechips.rocketchip.system.DefaultRV32Config.fir@199882.12]
  wire  _GEN_83; // @[TLB.scala 246:32:freechips.rocketchip.system.DefaultRV32Config.fir@199882.12]
  wire  _GEN_950; // @[TLB.scala 122:16:freechips.rocketchip.system.DefaultRV32Config.fir@199891.12]
  wire  _GEN_84; // @[TLB.scala 122:16:freechips.rocketchip.system.DefaultRV32Config.fir@199891.12]
  wire  _GEN_951; // @[TLB.scala 122:16:freechips.rocketchip.system.DefaultRV32Config.fir@199891.12]
  wire  _GEN_85; // @[TLB.scala 122:16:freechips.rocketchip.system.DefaultRV32Config.fir@199891.12]
  wire  _GEN_952; // @[TLB.scala 122:16:freechips.rocketchip.system.DefaultRV32Config.fir@199891.12]
  wire  _GEN_86; // @[TLB.scala 122:16:freechips.rocketchip.system.DefaultRV32Config.fir@199891.12]
  wire  _GEN_953; // @[TLB.scala 122:16:freechips.rocketchip.system.DefaultRV32Config.fir@199891.12]
  wire  _GEN_87; // @[TLB.scala 122:16:freechips.rocketchip.system.DefaultRV32Config.fir@199891.12]
  wire  _GEN_92; // @[TLB.scala 245:72:freechips.rocketchip.system.DefaultRV32Config.fir@199880.10]
  wire  _GEN_93; // @[TLB.scala 245:72:freechips.rocketchip.system.DefaultRV32Config.fir@199880.10]
  wire  _GEN_94; // @[TLB.scala 245:72:freechips.rocketchip.system.DefaultRV32Config.fir@199880.10]
  wire  _GEN_95; // @[TLB.scala 245:72:freechips.rocketchip.system.DefaultRV32Config.fir@199880.10]
  wire  _T_1063; // @[TLB.scala 245:65:freechips.rocketchip.system.DefaultRV32Config.fir@199909.10]
  wire  _GEN_102; // @[TLB.scala 246:32:freechips.rocketchip.system.DefaultRV32Config.fir@199912.12]
  wire  _GEN_103; // @[TLB.scala 246:32:freechips.rocketchip.system.DefaultRV32Config.fir@199912.12]
  wire  _GEN_104; // @[TLB.scala 246:32:freechips.rocketchip.system.DefaultRV32Config.fir@199912.12]
  wire  _GEN_105; // @[TLB.scala 246:32:freechips.rocketchip.system.DefaultRV32Config.fir@199912.12]
  wire  _GEN_106; // @[TLB.scala 122:16:freechips.rocketchip.system.DefaultRV32Config.fir@199921.12]
  wire  _GEN_107; // @[TLB.scala 122:16:freechips.rocketchip.system.DefaultRV32Config.fir@199921.12]
  wire  _GEN_108; // @[TLB.scala 122:16:freechips.rocketchip.system.DefaultRV32Config.fir@199921.12]
  wire  _GEN_109; // @[TLB.scala 122:16:freechips.rocketchip.system.DefaultRV32Config.fir@199921.12]
  wire  _GEN_114; // @[TLB.scala 245:72:freechips.rocketchip.system.DefaultRV32Config.fir@199910.10]
  wire  _GEN_115; // @[TLB.scala 245:72:freechips.rocketchip.system.DefaultRV32Config.fir@199910.10]
  wire  _GEN_116; // @[TLB.scala 245:72:freechips.rocketchip.system.DefaultRV32Config.fir@199910.10]
  wire  _GEN_117; // @[TLB.scala 245:72:freechips.rocketchip.system.DefaultRV32Config.fir@199910.10]
  wire  _T_1081; // @[TLB.scala 245:65:freechips.rocketchip.system.DefaultRV32Config.fir@199939.10]
  wire  _GEN_124; // @[TLB.scala 246:32:freechips.rocketchip.system.DefaultRV32Config.fir@199942.12]
  wire  _GEN_125; // @[TLB.scala 246:32:freechips.rocketchip.system.DefaultRV32Config.fir@199942.12]
  wire  _GEN_126; // @[TLB.scala 246:32:freechips.rocketchip.system.DefaultRV32Config.fir@199942.12]
  wire  _GEN_127; // @[TLB.scala 246:32:freechips.rocketchip.system.DefaultRV32Config.fir@199942.12]
  wire  _GEN_128; // @[TLB.scala 122:16:freechips.rocketchip.system.DefaultRV32Config.fir@199951.12]
  wire  _GEN_129; // @[TLB.scala 122:16:freechips.rocketchip.system.DefaultRV32Config.fir@199951.12]
  wire  _GEN_130; // @[TLB.scala 122:16:freechips.rocketchip.system.DefaultRV32Config.fir@199951.12]
  wire  _GEN_131; // @[TLB.scala 122:16:freechips.rocketchip.system.DefaultRV32Config.fir@199951.12]
  wire  _GEN_136; // @[TLB.scala 245:72:freechips.rocketchip.system.DefaultRV32Config.fir@199940.10]
  wire  _GEN_137; // @[TLB.scala 245:72:freechips.rocketchip.system.DefaultRV32Config.fir@199940.10]
  wire  _GEN_138; // @[TLB.scala 245:72:freechips.rocketchip.system.DefaultRV32Config.fir@199940.10]
  wire  _GEN_139; // @[TLB.scala 245:72:freechips.rocketchip.system.DefaultRV32Config.fir@199940.10]
  wire  _T_1099; // @[TLB.scala 245:65:freechips.rocketchip.system.DefaultRV32Config.fir@199969.10]
  wire  _GEN_146; // @[TLB.scala 246:32:freechips.rocketchip.system.DefaultRV32Config.fir@199972.12]
  wire  _GEN_147; // @[TLB.scala 246:32:freechips.rocketchip.system.DefaultRV32Config.fir@199972.12]
  wire  _GEN_148; // @[TLB.scala 246:32:freechips.rocketchip.system.DefaultRV32Config.fir@199972.12]
  wire  _GEN_149; // @[TLB.scala 246:32:freechips.rocketchip.system.DefaultRV32Config.fir@199972.12]
  wire  _GEN_150; // @[TLB.scala 122:16:freechips.rocketchip.system.DefaultRV32Config.fir@199981.12]
  wire  _GEN_151; // @[TLB.scala 122:16:freechips.rocketchip.system.DefaultRV32Config.fir@199981.12]
  wire  _GEN_152; // @[TLB.scala 122:16:freechips.rocketchip.system.DefaultRV32Config.fir@199981.12]
  wire  _GEN_153; // @[TLB.scala 122:16:freechips.rocketchip.system.DefaultRV32Config.fir@199981.12]
  wire  _GEN_158; // @[TLB.scala 245:72:freechips.rocketchip.system.DefaultRV32Config.fir@199970.10]
  wire  _GEN_159; // @[TLB.scala 245:72:freechips.rocketchip.system.DefaultRV32Config.fir@199970.10]
  wire  _GEN_160; // @[TLB.scala 245:72:freechips.rocketchip.system.DefaultRV32Config.fir@199970.10]
  wire  _GEN_161; // @[TLB.scala 245:72:freechips.rocketchip.system.DefaultRV32Config.fir@199970.10]
  wire  _T_1117; // @[TLB.scala 245:65:freechips.rocketchip.system.DefaultRV32Config.fir@199999.10]
  wire  _GEN_168; // @[TLB.scala 246:32:freechips.rocketchip.system.DefaultRV32Config.fir@200002.12]
  wire  _GEN_169; // @[TLB.scala 246:32:freechips.rocketchip.system.DefaultRV32Config.fir@200002.12]
  wire  _GEN_170; // @[TLB.scala 246:32:freechips.rocketchip.system.DefaultRV32Config.fir@200002.12]
  wire  _GEN_171; // @[TLB.scala 246:32:freechips.rocketchip.system.DefaultRV32Config.fir@200002.12]
  wire  _GEN_172; // @[TLB.scala 122:16:freechips.rocketchip.system.DefaultRV32Config.fir@200011.12]
  wire  _GEN_173; // @[TLB.scala 122:16:freechips.rocketchip.system.DefaultRV32Config.fir@200011.12]
  wire  _GEN_174; // @[TLB.scala 122:16:freechips.rocketchip.system.DefaultRV32Config.fir@200011.12]
  wire  _GEN_175; // @[TLB.scala 122:16:freechips.rocketchip.system.DefaultRV32Config.fir@200011.12]
  wire  _GEN_180; // @[TLB.scala 245:72:freechips.rocketchip.system.DefaultRV32Config.fir@200000.10]
  wire  _GEN_181; // @[TLB.scala 245:72:freechips.rocketchip.system.DefaultRV32Config.fir@200000.10]
  wire  _GEN_182; // @[TLB.scala 245:72:freechips.rocketchip.system.DefaultRV32Config.fir@200000.10]
  wire  _GEN_183; // @[TLB.scala 245:72:freechips.rocketchip.system.DefaultRV32Config.fir@200000.10]
  wire  _T_1135; // @[TLB.scala 245:65:freechips.rocketchip.system.DefaultRV32Config.fir@200029.10]
  wire  _GEN_190; // @[TLB.scala 246:32:freechips.rocketchip.system.DefaultRV32Config.fir@200032.12]
  wire  _GEN_191; // @[TLB.scala 246:32:freechips.rocketchip.system.DefaultRV32Config.fir@200032.12]
  wire  _GEN_192; // @[TLB.scala 246:32:freechips.rocketchip.system.DefaultRV32Config.fir@200032.12]
  wire  _GEN_193; // @[TLB.scala 246:32:freechips.rocketchip.system.DefaultRV32Config.fir@200032.12]
  wire  _GEN_194; // @[TLB.scala 122:16:freechips.rocketchip.system.DefaultRV32Config.fir@200041.12]
  wire  _GEN_195; // @[TLB.scala 122:16:freechips.rocketchip.system.DefaultRV32Config.fir@200041.12]
  wire  _GEN_196; // @[TLB.scala 122:16:freechips.rocketchip.system.DefaultRV32Config.fir@200041.12]
  wire  _GEN_197; // @[TLB.scala 122:16:freechips.rocketchip.system.DefaultRV32Config.fir@200041.12]
  wire  _GEN_202; // @[TLB.scala 245:72:freechips.rocketchip.system.DefaultRV32Config.fir@200030.10]
  wire  _GEN_203; // @[TLB.scala 245:72:freechips.rocketchip.system.DefaultRV32Config.fir@200030.10]
  wire  _GEN_204; // @[TLB.scala 245:72:freechips.rocketchip.system.DefaultRV32Config.fir@200030.10]
  wire  _GEN_205; // @[TLB.scala 245:72:freechips.rocketchip.system.DefaultRV32Config.fir@200030.10]
  wire  _T_1153; // @[TLB.scala 245:65:freechips.rocketchip.system.DefaultRV32Config.fir@200059.10]
  wire  _GEN_212; // @[TLB.scala 246:32:freechips.rocketchip.system.DefaultRV32Config.fir@200062.12]
  wire  _GEN_213; // @[TLB.scala 246:32:freechips.rocketchip.system.DefaultRV32Config.fir@200062.12]
  wire  _GEN_214; // @[TLB.scala 246:32:freechips.rocketchip.system.DefaultRV32Config.fir@200062.12]
  wire  _GEN_215; // @[TLB.scala 246:32:freechips.rocketchip.system.DefaultRV32Config.fir@200062.12]
  wire  _GEN_216; // @[TLB.scala 122:16:freechips.rocketchip.system.DefaultRV32Config.fir@200071.12]
  wire  _GEN_217; // @[TLB.scala 122:16:freechips.rocketchip.system.DefaultRV32Config.fir@200071.12]
  wire  _GEN_218; // @[TLB.scala 122:16:freechips.rocketchip.system.DefaultRV32Config.fir@200071.12]
  wire  _GEN_219; // @[TLB.scala 122:16:freechips.rocketchip.system.DefaultRV32Config.fir@200071.12]
  wire  _GEN_224; // @[TLB.scala 245:72:freechips.rocketchip.system.DefaultRV32Config.fir@200060.10]
  wire  _GEN_225; // @[TLB.scala 245:72:freechips.rocketchip.system.DefaultRV32Config.fir@200060.10]
  wire  _GEN_226; // @[TLB.scala 245:72:freechips.rocketchip.system.DefaultRV32Config.fir@200060.10]
  wire  _GEN_227; // @[TLB.scala 245:72:freechips.rocketchip.system.DefaultRV32Config.fir@200060.10]
  wire  _T_1171; // @[TLB.scala 245:65:freechips.rocketchip.system.DefaultRV32Config.fir@200089.10]
  wire  _GEN_234; // @[TLB.scala 246:32:freechips.rocketchip.system.DefaultRV32Config.fir@200092.12]
  wire  _GEN_235; // @[TLB.scala 246:32:freechips.rocketchip.system.DefaultRV32Config.fir@200092.12]
  wire  _GEN_236; // @[TLB.scala 246:32:freechips.rocketchip.system.DefaultRV32Config.fir@200092.12]
  wire  _GEN_237; // @[TLB.scala 246:32:freechips.rocketchip.system.DefaultRV32Config.fir@200092.12]
  wire  _GEN_238; // @[TLB.scala 122:16:freechips.rocketchip.system.DefaultRV32Config.fir@200101.12]
  wire  _GEN_239; // @[TLB.scala 122:16:freechips.rocketchip.system.DefaultRV32Config.fir@200101.12]
  wire  _GEN_240; // @[TLB.scala 122:16:freechips.rocketchip.system.DefaultRV32Config.fir@200101.12]
  wire  _GEN_241; // @[TLB.scala 122:16:freechips.rocketchip.system.DefaultRV32Config.fir@200101.12]
  wire  _GEN_246; // @[TLB.scala 245:72:freechips.rocketchip.system.DefaultRV32Config.fir@200090.10]
  wire  _GEN_247; // @[TLB.scala 245:72:freechips.rocketchip.system.DefaultRV32Config.fir@200090.10]
  wire  _GEN_248; // @[TLB.scala 245:72:freechips.rocketchip.system.DefaultRV32Config.fir@200090.10]
  wire  _GEN_249; // @[TLB.scala 245:72:freechips.rocketchip.system.DefaultRV32Config.fir@200090.10]
  wire  _GEN_258; // @[TLB.scala 239:54:freechips.rocketchip.system.DefaultRV32Config.fir@199787.8]
  wire  _GEN_262; // @[TLB.scala 239:54:freechips.rocketchip.system.DefaultRV32Config.fir@199787.8]
  wire  _GEN_266; // @[TLB.scala 239:54:freechips.rocketchip.system.DefaultRV32Config.fir@199787.8]
  wire  _GEN_270; // @[TLB.scala 239:54:freechips.rocketchip.system.DefaultRV32Config.fir@199787.8]
  wire  _GEN_272; // @[TLB.scala 239:54:freechips.rocketchip.system.DefaultRV32Config.fir@199787.8]
  wire  _GEN_273; // @[TLB.scala 239:54:freechips.rocketchip.system.DefaultRV32Config.fir@199787.8]
  wire  _GEN_274; // @[TLB.scala 239:54:freechips.rocketchip.system.DefaultRV32Config.fir@199787.8]
  wire  _GEN_275; // @[TLB.scala 239:54:freechips.rocketchip.system.DefaultRV32Config.fir@199787.8]
  wire  _GEN_282; // @[TLB.scala 239:54:freechips.rocketchip.system.DefaultRV32Config.fir@199787.8]
  wire  _GEN_283; // @[TLB.scala 239:54:freechips.rocketchip.system.DefaultRV32Config.fir@199787.8]
  wire  _GEN_284; // @[TLB.scala 239:54:freechips.rocketchip.system.DefaultRV32Config.fir@199787.8]
  wire  _GEN_285; // @[TLB.scala 239:54:freechips.rocketchip.system.DefaultRV32Config.fir@199787.8]
  wire  _GEN_292; // @[TLB.scala 239:54:freechips.rocketchip.system.DefaultRV32Config.fir@199787.8]
  wire  _GEN_293; // @[TLB.scala 239:54:freechips.rocketchip.system.DefaultRV32Config.fir@199787.8]
  wire  _GEN_294; // @[TLB.scala 239:54:freechips.rocketchip.system.DefaultRV32Config.fir@199787.8]
  wire  _GEN_295; // @[TLB.scala 239:54:freechips.rocketchip.system.DefaultRV32Config.fir@199787.8]
  wire  _GEN_302; // @[TLB.scala 239:54:freechips.rocketchip.system.DefaultRV32Config.fir@199787.8]
  wire  _GEN_303; // @[TLB.scala 239:54:freechips.rocketchip.system.DefaultRV32Config.fir@199787.8]
  wire  _GEN_304; // @[TLB.scala 239:54:freechips.rocketchip.system.DefaultRV32Config.fir@199787.8]
  wire  _GEN_305; // @[TLB.scala 239:54:freechips.rocketchip.system.DefaultRV32Config.fir@199787.8]
  wire  _GEN_312; // @[TLB.scala 239:54:freechips.rocketchip.system.DefaultRV32Config.fir@199787.8]
  wire  _GEN_313; // @[TLB.scala 239:54:freechips.rocketchip.system.DefaultRV32Config.fir@199787.8]
  wire  _GEN_314; // @[TLB.scala 239:54:freechips.rocketchip.system.DefaultRV32Config.fir@199787.8]
  wire  _GEN_315; // @[TLB.scala 239:54:freechips.rocketchip.system.DefaultRV32Config.fir@199787.8]
  wire  _GEN_322; // @[TLB.scala 239:54:freechips.rocketchip.system.DefaultRV32Config.fir@199787.8]
  wire  _GEN_323; // @[TLB.scala 239:54:freechips.rocketchip.system.DefaultRV32Config.fir@199787.8]
  wire  _GEN_324; // @[TLB.scala 239:54:freechips.rocketchip.system.DefaultRV32Config.fir@199787.8]
  wire  _GEN_325; // @[TLB.scala 239:54:freechips.rocketchip.system.DefaultRV32Config.fir@199787.8]
  wire  _GEN_332; // @[TLB.scala 239:54:freechips.rocketchip.system.DefaultRV32Config.fir@199787.8]
  wire  _GEN_333; // @[TLB.scala 239:54:freechips.rocketchip.system.DefaultRV32Config.fir@199787.8]
  wire  _GEN_334; // @[TLB.scala 239:54:freechips.rocketchip.system.DefaultRV32Config.fir@199787.8]
  wire  _GEN_335; // @[TLB.scala 239:54:freechips.rocketchip.system.DefaultRV32Config.fir@199787.8]
  wire  _GEN_342; // @[TLB.scala 239:54:freechips.rocketchip.system.DefaultRV32Config.fir@199787.8]
  wire  _GEN_343; // @[TLB.scala 239:54:freechips.rocketchip.system.DefaultRV32Config.fir@199787.8]
  wire  _GEN_344; // @[TLB.scala 239:54:freechips.rocketchip.system.DefaultRV32Config.fir@199787.8]
  wire  _GEN_345; // @[TLB.scala 239:54:freechips.rocketchip.system.DefaultRV32Config.fir@199787.8]
  wire  _GEN_354; // @[TLB.scala 237:68:freechips.rocketchip.system.DefaultRV32Config.fir@199763.6]
  wire  _GEN_358; // @[TLB.scala 237:68:freechips.rocketchip.system.DefaultRV32Config.fir@199763.6]
  wire  _GEN_362; // @[TLB.scala 237:68:freechips.rocketchip.system.DefaultRV32Config.fir@199763.6]
  wire  _GEN_366; // @[TLB.scala 237:68:freechips.rocketchip.system.DefaultRV32Config.fir@199763.6]
  wire  _GEN_370; // @[TLB.scala 237:68:freechips.rocketchip.system.DefaultRV32Config.fir@199763.6]
  wire  _GEN_372; // @[TLB.scala 237:68:freechips.rocketchip.system.DefaultRV32Config.fir@199763.6]
  wire  _GEN_373; // @[TLB.scala 237:68:freechips.rocketchip.system.DefaultRV32Config.fir@199763.6]
  wire  _GEN_374; // @[TLB.scala 237:68:freechips.rocketchip.system.DefaultRV32Config.fir@199763.6]
  wire  _GEN_375; // @[TLB.scala 237:68:freechips.rocketchip.system.DefaultRV32Config.fir@199763.6]
  wire  _GEN_382; // @[TLB.scala 237:68:freechips.rocketchip.system.DefaultRV32Config.fir@199763.6]
  wire  _GEN_383; // @[TLB.scala 237:68:freechips.rocketchip.system.DefaultRV32Config.fir@199763.6]
  wire  _GEN_384; // @[TLB.scala 237:68:freechips.rocketchip.system.DefaultRV32Config.fir@199763.6]
  wire  _GEN_385; // @[TLB.scala 237:68:freechips.rocketchip.system.DefaultRV32Config.fir@199763.6]
  wire  _GEN_392; // @[TLB.scala 237:68:freechips.rocketchip.system.DefaultRV32Config.fir@199763.6]
  wire  _GEN_393; // @[TLB.scala 237:68:freechips.rocketchip.system.DefaultRV32Config.fir@199763.6]
  wire  _GEN_394; // @[TLB.scala 237:68:freechips.rocketchip.system.DefaultRV32Config.fir@199763.6]
  wire  _GEN_395; // @[TLB.scala 237:68:freechips.rocketchip.system.DefaultRV32Config.fir@199763.6]
  wire  _GEN_402; // @[TLB.scala 237:68:freechips.rocketchip.system.DefaultRV32Config.fir@199763.6]
  wire  _GEN_403; // @[TLB.scala 237:68:freechips.rocketchip.system.DefaultRV32Config.fir@199763.6]
  wire  _GEN_404; // @[TLB.scala 237:68:freechips.rocketchip.system.DefaultRV32Config.fir@199763.6]
  wire  _GEN_405; // @[TLB.scala 237:68:freechips.rocketchip.system.DefaultRV32Config.fir@199763.6]
  wire  _GEN_412; // @[TLB.scala 237:68:freechips.rocketchip.system.DefaultRV32Config.fir@199763.6]
  wire  _GEN_413; // @[TLB.scala 237:68:freechips.rocketchip.system.DefaultRV32Config.fir@199763.6]
  wire  _GEN_414; // @[TLB.scala 237:68:freechips.rocketchip.system.DefaultRV32Config.fir@199763.6]
  wire  _GEN_415; // @[TLB.scala 237:68:freechips.rocketchip.system.DefaultRV32Config.fir@199763.6]
  wire  _GEN_422; // @[TLB.scala 237:68:freechips.rocketchip.system.DefaultRV32Config.fir@199763.6]
  wire  _GEN_423; // @[TLB.scala 237:68:freechips.rocketchip.system.DefaultRV32Config.fir@199763.6]
  wire  _GEN_424; // @[TLB.scala 237:68:freechips.rocketchip.system.DefaultRV32Config.fir@199763.6]
  wire  _GEN_425; // @[TLB.scala 237:68:freechips.rocketchip.system.DefaultRV32Config.fir@199763.6]
  wire  _GEN_432; // @[TLB.scala 237:68:freechips.rocketchip.system.DefaultRV32Config.fir@199763.6]
  wire  _GEN_433; // @[TLB.scala 237:68:freechips.rocketchip.system.DefaultRV32Config.fir@199763.6]
  wire  _GEN_434; // @[TLB.scala 237:68:freechips.rocketchip.system.DefaultRV32Config.fir@199763.6]
  wire  _GEN_435; // @[TLB.scala 237:68:freechips.rocketchip.system.DefaultRV32Config.fir@199763.6]
  wire  _GEN_442; // @[TLB.scala 237:68:freechips.rocketchip.system.DefaultRV32Config.fir@199763.6]
  wire  _GEN_443; // @[TLB.scala 237:68:freechips.rocketchip.system.DefaultRV32Config.fir@199763.6]
  wire  _GEN_444; // @[TLB.scala 237:68:freechips.rocketchip.system.DefaultRV32Config.fir@199763.6]
  wire  _GEN_445; // @[TLB.scala 237:68:freechips.rocketchip.system.DefaultRV32Config.fir@199763.6]
  wire  _GEN_454; // @[TLB.scala 217:42:freechips.rocketchip.system.DefaultRV32Config.fir@199722.4]
  wire  _GEN_458; // @[TLB.scala 217:42:freechips.rocketchip.system.DefaultRV32Config.fir@199722.4]
  wire  _GEN_462; // @[TLB.scala 217:42:freechips.rocketchip.system.DefaultRV32Config.fir@199722.4]
  wire  _GEN_466; // @[TLB.scala 217:42:freechips.rocketchip.system.DefaultRV32Config.fir@199722.4]
  wire  _GEN_470; // @[TLB.scala 217:42:freechips.rocketchip.system.DefaultRV32Config.fir@199722.4]
  wire  _GEN_472; // @[TLB.scala 217:42:freechips.rocketchip.system.DefaultRV32Config.fir@199722.4]
  wire  _GEN_473; // @[TLB.scala 217:42:freechips.rocketchip.system.DefaultRV32Config.fir@199722.4]
  wire  _GEN_474; // @[TLB.scala 217:42:freechips.rocketchip.system.DefaultRV32Config.fir@199722.4]
  wire  _GEN_475; // @[TLB.scala 217:42:freechips.rocketchip.system.DefaultRV32Config.fir@199722.4]
  wire  _GEN_482; // @[TLB.scala 217:42:freechips.rocketchip.system.DefaultRV32Config.fir@199722.4]
  wire  _GEN_483; // @[TLB.scala 217:42:freechips.rocketchip.system.DefaultRV32Config.fir@199722.4]
  wire  _GEN_484; // @[TLB.scala 217:42:freechips.rocketchip.system.DefaultRV32Config.fir@199722.4]
  wire  _GEN_485; // @[TLB.scala 217:42:freechips.rocketchip.system.DefaultRV32Config.fir@199722.4]
  wire  _GEN_492; // @[TLB.scala 217:42:freechips.rocketchip.system.DefaultRV32Config.fir@199722.4]
  wire  _GEN_493; // @[TLB.scala 217:42:freechips.rocketchip.system.DefaultRV32Config.fir@199722.4]
  wire  _GEN_494; // @[TLB.scala 217:42:freechips.rocketchip.system.DefaultRV32Config.fir@199722.4]
  wire  _GEN_495; // @[TLB.scala 217:42:freechips.rocketchip.system.DefaultRV32Config.fir@199722.4]
  wire  _GEN_502; // @[TLB.scala 217:42:freechips.rocketchip.system.DefaultRV32Config.fir@199722.4]
  wire  _GEN_503; // @[TLB.scala 217:42:freechips.rocketchip.system.DefaultRV32Config.fir@199722.4]
  wire  _GEN_504; // @[TLB.scala 217:42:freechips.rocketchip.system.DefaultRV32Config.fir@199722.4]
  wire  _GEN_505; // @[TLB.scala 217:42:freechips.rocketchip.system.DefaultRV32Config.fir@199722.4]
  wire  _GEN_512; // @[TLB.scala 217:42:freechips.rocketchip.system.DefaultRV32Config.fir@199722.4]
  wire  _GEN_513; // @[TLB.scala 217:42:freechips.rocketchip.system.DefaultRV32Config.fir@199722.4]
  wire  _GEN_514; // @[TLB.scala 217:42:freechips.rocketchip.system.DefaultRV32Config.fir@199722.4]
  wire  _GEN_515; // @[TLB.scala 217:42:freechips.rocketchip.system.DefaultRV32Config.fir@199722.4]
  wire  _GEN_522; // @[TLB.scala 217:42:freechips.rocketchip.system.DefaultRV32Config.fir@199722.4]
  wire  _GEN_523; // @[TLB.scala 217:42:freechips.rocketchip.system.DefaultRV32Config.fir@199722.4]
  wire  _GEN_524; // @[TLB.scala 217:42:freechips.rocketchip.system.DefaultRV32Config.fir@199722.4]
  wire  _GEN_525; // @[TLB.scala 217:42:freechips.rocketchip.system.DefaultRV32Config.fir@199722.4]
  wire  _GEN_532; // @[TLB.scala 217:42:freechips.rocketchip.system.DefaultRV32Config.fir@199722.4]
  wire  _GEN_533; // @[TLB.scala 217:42:freechips.rocketchip.system.DefaultRV32Config.fir@199722.4]
  wire  _GEN_534; // @[TLB.scala 217:42:freechips.rocketchip.system.DefaultRV32Config.fir@199722.4]
  wire  _GEN_535; // @[TLB.scala 217:42:freechips.rocketchip.system.DefaultRV32Config.fir@199722.4]
  wire  _GEN_542; // @[TLB.scala 217:42:freechips.rocketchip.system.DefaultRV32Config.fir@199722.4]
  wire  _GEN_543; // @[TLB.scala 217:42:freechips.rocketchip.system.DefaultRV32Config.fir@199722.4]
  wire  _GEN_544; // @[TLB.scala 217:42:freechips.rocketchip.system.DefaultRV32Config.fir@199722.4]
  wire  _GEN_545; // @[TLB.scala 217:42:freechips.rocketchip.system.DefaultRV32Config.fir@199722.4]
  wire [5:0] _T_1659; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@201191.4]
  wire [13:0] ptw_ae_array; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@201199.4]
  wire [5:0] _T_1673; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@201206.4]
  wire [12:0] _T_1680; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@201213.4]
  wire [12:0] _T_1694; // @[TLB.scala 256:98:freechips.rocketchip.system.DefaultRV32Config.fir@201227.4]
  wire [12:0] priv_x_ok; // @[TLB.scala 257:22:freechips.rocketchip.system.DefaultRV32Config.fir@201255.4]
  wire [5:0] _T_1737; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@201272.4]
  wire [12:0] _T_1744; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@201279.4]
  wire [12:0] _T_1773; // @[TLB.scala 260:39:freechips.rocketchip.system.DefaultRV32Config.fir@201310.4]
  wire [13:0] x_array; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@201311.4]
  wire [13:0] _T_1788; // @[TLB.scala 261:89:freechips.rocketchip.system.DefaultRV32Config.fir@201326.4]
  wire [1:0] _T_1805; // @[Bitwise.scala 72:12:freechips.rocketchip.system.DefaultRV32Config.fir@201345.4]
  wire [5:0] _T_1810; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@201350.4]
  wire [13:0] _T_1817; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@201357.4]
  wire [13:0] px_array; // @[TLB.scala 263:87:freechips.rocketchip.system.DefaultRV32Config.fir@201359.4]
  wire [1:0] _T_1833; // @[Bitwise.scala 72:12:freechips.rocketchip.system.DefaultRV32Config.fir@201375.4]
  wire [5:0] _T_1838; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@201380.4]
  wire [13:0] c_array; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@201387.4]
  wire [13:0] _T_2003; // @[TLB.scala 313:33:freechips.rocketchip.system.DefaultRV32Config.fir@201570.4]
  wire [13:0] pf_inst_array; // @[TLB.scala 313:23:freechips.rocketchip.system.DefaultRV32Config.fir@201571.4]
  wire  tlb_hit; // @[TLB.scala 315:27:freechips.rocketchip.system.DefaultRV32Config.fir@201572.4]
  wire  _T_2006; // @[TLB.scala 316:43:freechips.rocketchip.system.DefaultRV32Config.fir@201575.4]
  wire  tlb_miss; // @[TLB.scala 316:40:freechips.rocketchip.system.DefaultRV32Config.fir@201576.4]
  reg [6:0] _T_2007; // @[Replacement.scala 158:30:freechips.rocketchip.system.DefaultRV32Config.fir@201577.4]
  reg [2:0] _T_2008; // @[Replacement.scala 158:30:freechips.rocketchip.system.DefaultRV32Config.fir@201578.4]
  wire  _T_2009; // @[TLB.scala 320:22:freechips.rocketchip.system.DefaultRV32Config.fir@201579.4]
  wire  _T_2010; // @[package.scala 64:59:freechips.rocketchip.system.DefaultRV32Config.fir@201581.6]
  wire  _T_2011; // @[package.scala 64:59:freechips.rocketchip.system.DefaultRV32Config.fir@201582.6]
  wire  _T_2012; // @[package.scala 64:59:freechips.rocketchip.system.DefaultRV32Config.fir@201583.6]
  wire  _T_2013; // @[package.scala 64:59:freechips.rocketchip.system.DefaultRV32Config.fir@201584.6]
  wire  _T_2014; // @[package.scala 64:59:freechips.rocketchip.system.DefaultRV32Config.fir@201585.6]
  wire  _T_2015; // @[package.scala 64:59:freechips.rocketchip.system.DefaultRV32Config.fir@201586.6]
  wire  _T_2016; // @[package.scala 64:59:freechips.rocketchip.system.DefaultRV32Config.fir@201587.6]
  wire [7:0] _T_2023; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@201595.8]
  wire  _T_2026; // @[OneHot.scala 32:14:freechips.rocketchip.system.DefaultRV32Config.fir@201598.8]
  wire [3:0] _T_2027; // @[OneHot.scala 32:28:freechips.rocketchip.system.DefaultRV32Config.fir@201599.8]
  wire  _T_2030; // @[OneHot.scala 32:14:freechips.rocketchip.system.DefaultRV32Config.fir@201602.8]
  wire [1:0] _T_2031; // @[OneHot.scala 32:28:freechips.rocketchip.system.DefaultRV32Config.fir@201603.8]
  wire [2:0] _T_2034; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@201606.8]
  wire  _T_2037; // @[Replacement.scala 186:33:freechips.rocketchip.system.DefaultRV32Config.fir@201609.8]
  wire  _T_2042; // @[Replacement.scala 186:33:freechips.rocketchip.system.DefaultRV32Config.fir@201614.8]
  wire  _T_2047; // @[Replacement.scala 208:7:freechips.rocketchip.system.DefaultRV32Config.fir@201619.8]
  wire  _T_2048; // @[Replacement.scala 193:16:freechips.rocketchip.system.DefaultRV32Config.fir@201620.8]
  wire  _T_2052; // @[Replacement.scala 196:16:freechips.rocketchip.system.DefaultRV32Config.fir@201624.8]
  wire [2:0] _T_2054; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@201626.8]
  wire [2:0] _T_2055; // @[Replacement.scala 193:16:freechips.rocketchip.system.DefaultRV32Config.fir@201627.8]
  wire  _T_2064; // @[Replacement.scala 193:16:freechips.rocketchip.system.DefaultRV32Config.fir@201636.8]
  wire  _T_2068; // @[Replacement.scala 196:16:freechips.rocketchip.system.DefaultRV32Config.fir@201640.8]
  wire [2:0] _T_2070; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@201642.8]
  wire [2:0] _T_2071; // @[Replacement.scala 196:16:freechips.rocketchip.system.DefaultRV32Config.fir@201643.8]
  wire [6:0] _T_2073; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@201645.8]
  wire  _T_2074; // @[package.scala 64:59:freechips.rocketchip.system.DefaultRV32Config.fir@201648.6]
  wire  _T_2075; // @[package.scala 64:59:freechips.rocketchip.system.DefaultRV32Config.fir@201649.6]
  wire  _T_2076; // @[package.scala 64:59:freechips.rocketchip.system.DefaultRV32Config.fir@201650.6]
  wire [3:0] _T_2079; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@201654.8]
  wire  _T_2082; // @[OneHot.scala 32:14:freechips.rocketchip.system.DefaultRV32Config.fir@201657.8]
  wire [1:0] _T_2083; // @[OneHot.scala 32:28:freechips.rocketchip.system.DefaultRV32Config.fir@201658.8]
  wire [1:0] _T_2085; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@201660.8]
  wire  _T_2088; // @[Replacement.scala 186:33:freechips.rocketchip.system.DefaultRV32Config.fir@201663.8]
  wire  _T_2093; // @[Replacement.scala 208:7:freechips.rocketchip.system.DefaultRV32Config.fir@201668.8]
  wire  _T_2094; // @[Replacement.scala 193:16:freechips.rocketchip.system.DefaultRV32Config.fir@201669.8]
  wire  _T_2098; // @[Replacement.scala 196:16:freechips.rocketchip.system.DefaultRV32Config.fir@201673.8]
  wire [2:0] _T_2100; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@201675.8]
  wire  _T_2110; // @[Misc.scala 182:16:freechips.rocketchip.system.DefaultRV32Config.fir@201688.4]
  wire  _T_2112; // @[Misc.scala 182:61:freechips.rocketchip.system.DefaultRV32Config.fir@201690.4]
  wire  _T_2114; // @[Misc.scala 182:16:freechips.rocketchip.system.DefaultRV32Config.fir@201692.4]
  wire  _T_2116; // @[Misc.scala 182:61:freechips.rocketchip.system.DefaultRV32Config.fir@201694.4]
  wire  _T_2117; // @[Misc.scala 182:49:freechips.rocketchip.system.DefaultRV32Config.fir@201695.4]
  wire  _T_2126; // @[Misc.scala 182:16:freechips.rocketchip.system.DefaultRV32Config.fir@201704.4]
  wire  _T_2128; // @[Misc.scala 182:61:freechips.rocketchip.system.DefaultRV32Config.fir@201706.4]
  wire  _T_2130; // @[Misc.scala 182:16:freechips.rocketchip.system.DefaultRV32Config.fir@201708.4]
  wire  _T_2132; // @[Misc.scala 182:61:freechips.rocketchip.system.DefaultRV32Config.fir@201710.4]
  wire  _T_2133; // @[Misc.scala 182:49:freechips.rocketchip.system.DefaultRV32Config.fir@201711.4]
  wire  _T_2134; // @[Misc.scala 182:16:freechips.rocketchip.system.DefaultRV32Config.fir@201712.4]
  wire  _T_2135; // @[Misc.scala 182:37:freechips.rocketchip.system.DefaultRV32Config.fir@201713.4]
  wire  _T_2136; // @[Misc.scala 182:61:freechips.rocketchip.system.DefaultRV32Config.fir@201714.4]
  wire  _T_2137; // @[Misc.scala 182:49:freechips.rocketchip.system.DefaultRV32Config.fir@201715.4]
  wire  _T_2147; // @[Misc.scala 182:16:freechips.rocketchip.system.DefaultRV32Config.fir@201725.4]
  wire  _T_2149; // @[Misc.scala 182:61:freechips.rocketchip.system.DefaultRV32Config.fir@201727.4]
  wire  _T_2151; // @[Misc.scala 182:16:freechips.rocketchip.system.DefaultRV32Config.fir@201729.4]
  wire  _T_2153; // @[Misc.scala 182:61:freechips.rocketchip.system.DefaultRV32Config.fir@201731.4]
  wire  _T_2154; // @[Misc.scala 182:49:freechips.rocketchip.system.DefaultRV32Config.fir@201732.4]
  wire  _T_2161; // @[Misc.scala 182:16:freechips.rocketchip.system.DefaultRV32Config.fir@201739.4]
  wire  _T_2163; // @[Misc.scala 182:61:freechips.rocketchip.system.DefaultRV32Config.fir@201741.4]
  wire  _T_2170; // @[Misc.scala 182:16:freechips.rocketchip.system.DefaultRV32Config.fir@201748.4]
  wire  _T_2172; // @[Misc.scala 182:61:freechips.rocketchip.system.DefaultRV32Config.fir@201750.4]
  wire  _T_2174; // @[Misc.scala 182:16:freechips.rocketchip.system.DefaultRV32Config.fir@201752.4]
  wire  _T_2175; // @[Misc.scala 182:37:freechips.rocketchip.system.DefaultRV32Config.fir@201753.4]
  wire  _T_2176; // @[Misc.scala 182:61:freechips.rocketchip.system.DefaultRV32Config.fir@201754.4]
  wire  _T_2177; // @[Misc.scala 182:49:freechips.rocketchip.system.DefaultRV32Config.fir@201755.4]
  wire  _T_2178; // @[Misc.scala 182:16:freechips.rocketchip.system.DefaultRV32Config.fir@201756.4]
  wire  _T_2179; // @[Misc.scala 182:37:freechips.rocketchip.system.DefaultRV32Config.fir@201757.4]
  wire  _T_2180; // @[Misc.scala 182:61:freechips.rocketchip.system.DefaultRV32Config.fir@201758.4]
  wire  _T_2181; // @[Misc.scala 182:49:freechips.rocketchip.system.DefaultRV32Config.fir@201759.4]
  wire  _T_2183; // @[Misc.scala 182:37:freechips.rocketchip.system.DefaultRV32Config.fir@201761.4]
  wire  _T_2184; // @[Misc.scala 182:61:freechips.rocketchip.system.DefaultRV32Config.fir@201762.4]
  wire  multipleHits; // @[Misc.scala 182:49:freechips.rocketchip.system.DefaultRV32Config.fir@201763.4]
  wire [13:0] _T_2194; // @[TLB.scala 335:47:freechips.rocketchip.system.DefaultRV32Config.fir@201776.4]
  wire [13:0] _T_2201; // @[TLB.scala 338:23:freechips.rocketchip.system.DefaultRV32Config.fir@201786.4]
  wire [13:0] _T_2202; // @[TLB.scala 338:33:freechips.rocketchip.system.DefaultRV32Config.fir@201787.4]
  wire [13:0] _T_2208; // @[TLB.scala 342:33:freechips.rocketchip.system.DefaultRV32Config.fir@201797.4]
  wire  _T_2215; // @[TLB.scala 345:29:freechips.rocketchip.system.DefaultRV32Config.fir@201807.4]
  wire  _T_2221; // @[Decoupled.scala 40:37:freechips.rocketchip.system.DefaultRV32Config.fir@201818.4]
  wire  _T_2222; // @[TLB.scala 354:25:freechips.rocketchip.system.DefaultRV32Config.fir@201819.4]
  wire  _T_2228; // @[Replacement.scala 240:16:freechips.rocketchip.system.DefaultRV32Config.fir@201828.6]
  wire [1:0] _T_2229; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@201829.6]
  wire [3:0] _T_2232; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@201832.6]
  wire  _T_2233; // @[TLB.scala 402:16:freechips.rocketchip.system.DefaultRV32Config.fir@201833.6]
  wire [3:0] _T_2234; // @[TLB.scala 402:43:freechips.rocketchip.system.DefaultRV32Config.fir@201834.6]
  wire  _T_2251; // @[Replacement.scala 240:16:freechips.rocketchip.system.DefaultRV32Config.fir@201852.6]
  wire [1:0] _T_2252; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@201853.6]
  wire  _T_2258; // @[Replacement.scala 240:16:freechips.rocketchip.system.DefaultRV32Config.fir@201859.6]
  wire [1:0] _T_2259; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@201860.6]
  wire [1:0] _T_2260; // @[Replacement.scala 240:16:freechips.rocketchip.system.DefaultRV32Config.fir@201861.6]
  wire [2:0] _T_2261; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@201862.6]
  wire [7:0] _T_2292; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@201893.6]
  wire  _T_2293; // @[TLB.scala 402:16:freechips.rocketchip.system.DefaultRV32Config.fir@201894.6]
  wire [7:0] _T_2294; // @[TLB.scala 402:43:freechips.rocketchip.system.DefaultRV32Config.fir@201895.6]
  wire  _T_2338; // @[TLB.scala 368:17:freechips.rocketchip.system.DefaultRV32Config.fir@201954.4]
  wire  _T_2339; // @[TLB.scala 368:28:freechips.rocketchip.system.DefaultRV32Config.fir@201955.4]
  wire  _T_2340; // @[TLB.scala 376:14:freechips.rocketchip.system.DefaultRV32Config.fir@201963.6]
  wire  _T_2342; // @[TLB.scala 376:72:freechips.rocketchip.system.DefaultRV32Config.fir@201965.6]
  wire  _T_2343; // @[TLB.scala 376:34:freechips.rocketchip.system.DefaultRV32Config.fir@201966.6]
  wire  _T_2345; // @[TLB.scala 376:13:freechips.rocketchip.system.DefaultRV32Config.fir@201968.6]
  wire  _T_2346; // @[TLB.scala 376:13:freechips.rocketchip.system.DefaultRV32Config.fir@201969.6]
  wire  _T_2353; // @[TLB.scala 135:61:freechips.rocketchip.system.DefaultRV32Config.fir@201984.8]
  wire  _T_2498; // @[TLB.scala 143:13:freechips.rocketchip.system.DefaultRV32Config.fir@202298.10]
  wire  _GEN_648; // @[TLB.scala 143:19:freechips.rocketchip.system.DefaultRV32Config.fir@202299.10]
  wire  _T_2499; // @[TLB.scala 143:13:freechips.rocketchip.system.DefaultRV32Config.fir@202302.10]
  wire  _GEN_649; // @[TLB.scala 143:19:freechips.rocketchip.system.DefaultRV32Config.fir@202303.10]
  wire  _T_2500; // @[TLB.scala 143:13:freechips.rocketchip.system.DefaultRV32Config.fir@202306.10]
  wire  _GEN_650; // @[TLB.scala 143:19:freechips.rocketchip.system.DefaultRV32Config.fir@202307.10]
  wire  _T_2501; // @[TLB.scala 143:13:freechips.rocketchip.system.DefaultRV32Config.fir@202310.10]
  wire  _GEN_651; // @[TLB.scala 143:19:freechips.rocketchip.system.DefaultRV32Config.fir@202311.10]
  wire  _GEN_652; // @[TLB.scala 379:40:freechips.rocketchip.system.DefaultRV32Config.fir@202149.8]
  wire  _GEN_653; // @[TLB.scala 379:40:freechips.rocketchip.system.DefaultRV32Config.fir@202149.8]
  wire  _GEN_654; // @[TLB.scala 379:40:freechips.rocketchip.system.DefaultRV32Config.fir@202149.8]
  wire  _GEN_655; // @[TLB.scala 379:40:freechips.rocketchip.system.DefaultRV32Config.fir@202149.8]
  wire  _T_2508; // @[TLB.scala 135:61:freechips.rocketchip.system.DefaultRV32Config.fir@202331.8]
  wire  _T_2653; // @[TLB.scala 143:13:freechips.rocketchip.system.DefaultRV32Config.fir@202645.10]
  wire  _GEN_676; // @[TLB.scala 143:19:freechips.rocketchip.system.DefaultRV32Config.fir@202646.10]
  wire  _T_2654; // @[TLB.scala 143:13:freechips.rocketchip.system.DefaultRV32Config.fir@202649.10]
  wire  _GEN_677; // @[TLB.scala 143:19:freechips.rocketchip.system.DefaultRV32Config.fir@202650.10]
  wire  _T_2655; // @[TLB.scala 143:13:freechips.rocketchip.system.DefaultRV32Config.fir@202653.10]
  wire  _GEN_678; // @[TLB.scala 143:19:freechips.rocketchip.system.DefaultRV32Config.fir@202654.10]
  wire  _T_2656; // @[TLB.scala 143:13:freechips.rocketchip.system.DefaultRV32Config.fir@202657.10]
  wire  _GEN_679; // @[TLB.scala 143:19:freechips.rocketchip.system.DefaultRV32Config.fir@202658.10]
  wire  _GEN_680; // @[TLB.scala 379:40:freechips.rocketchip.system.DefaultRV32Config.fir@202496.8]
  wire  _GEN_681; // @[TLB.scala 379:40:freechips.rocketchip.system.DefaultRV32Config.fir@202496.8]
  wire  _GEN_682; // @[TLB.scala 379:40:freechips.rocketchip.system.DefaultRV32Config.fir@202496.8]
  wire  _GEN_683; // @[TLB.scala 379:40:freechips.rocketchip.system.DefaultRV32Config.fir@202496.8]
  wire  _T_2663; // @[TLB.scala 135:61:freechips.rocketchip.system.DefaultRV32Config.fir@202678.8]
  wire  _T_2808; // @[TLB.scala 143:13:freechips.rocketchip.system.DefaultRV32Config.fir@202992.10]
  wire  _GEN_704; // @[TLB.scala 143:19:freechips.rocketchip.system.DefaultRV32Config.fir@202993.10]
  wire  _T_2809; // @[TLB.scala 143:13:freechips.rocketchip.system.DefaultRV32Config.fir@202996.10]
  wire  _GEN_705; // @[TLB.scala 143:19:freechips.rocketchip.system.DefaultRV32Config.fir@202997.10]
  wire  _T_2810; // @[TLB.scala 143:13:freechips.rocketchip.system.DefaultRV32Config.fir@203000.10]
  wire  _GEN_706; // @[TLB.scala 143:19:freechips.rocketchip.system.DefaultRV32Config.fir@203001.10]
  wire  _T_2811; // @[TLB.scala 143:13:freechips.rocketchip.system.DefaultRV32Config.fir@203004.10]
  wire  _GEN_707; // @[TLB.scala 143:19:freechips.rocketchip.system.DefaultRV32Config.fir@203005.10]
  wire  _GEN_708; // @[TLB.scala 379:40:freechips.rocketchip.system.DefaultRV32Config.fir@202843.8]
  wire  _GEN_709; // @[TLB.scala 379:40:freechips.rocketchip.system.DefaultRV32Config.fir@202843.8]
  wire  _GEN_710; // @[TLB.scala 379:40:freechips.rocketchip.system.DefaultRV32Config.fir@202843.8]
  wire  _GEN_711; // @[TLB.scala 379:40:freechips.rocketchip.system.DefaultRV32Config.fir@202843.8]
  wire  _T_2818; // @[TLB.scala 135:61:freechips.rocketchip.system.DefaultRV32Config.fir@203025.8]
  wire  _T_2963; // @[TLB.scala 143:13:freechips.rocketchip.system.DefaultRV32Config.fir@203339.10]
  wire  _GEN_732; // @[TLB.scala 143:19:freechips.rocketchip.system.DefaultRV32Config.fir@203340.10]
  wire  _T_2964; // @[TLB.scala 143:13:freechips.rocketchip.system.DefaultRV32Config.fir@203343.10]
  wire  _GEN_733; // @[TLB.scala 143:19:freechips.rocketchip.system.DefaultRV32Config.fir@203344.10]
  wire  _T_2965; // @[TLB.scala 143:13:freechips.rocketchip.system.DefaultRV32Config.fir@203347.10]
  wire  _GEN_734; // @[TLB.scala 143:19:freechips.rocketchip.system.DefaultRV32Config.fir@203348.10]
  wire  _T_2966; // @[TLB.scala 143:13:freechips.rocketchip.system.DefaultRV32Config.fir@203351.10]
  wire  _GEN_735; // @[TLB.scala 143:19:freechips.rocketchip.system.DefaultRV32Config.fir@203352.10]
  wire  _GEN_736; // @[TLB.scala 379:40:freechips.rocketchip.system.DefaultRV32Config.fir@203190.8]
  wire  _GEN_737; // @[TLB.scala 379:40:freechips.rocketchip.system.DefaultRV32Config.fir@203190.8]
  wire  _GEN_738; // @[TLB.scala 379:40:freechips.rocketchip.system.DefaultRV32Config.fir@203190.8]
  wire  _GEN_739; // @[TLB.scala 379:40:freechips.rocketchip.system.DefaultRV32Config.fir@203190.8]
  wire  _T_2973; // @[TLB.scala 135:61:freechips.rocketchip.system.DefaultRV32Config.fir@203372.8]
  wire  _T_3118; // @[TLB.scala 143:13:freechips.rocketchip.system.DefaultRV32Config.fir@203686.10]
  wire  _GEN_760; // @[TLB.scala 143:19:freechips.rocketchip.system.DefaultRV32Config.fir@203687.10]
  wire  _T_3119; // @[TLB.scala 143:13:freechips.rocketchip.system.DefaultRV32Config.fir@203690.10]
  wire  _GEN_761; // @[TLB.scala 143:19:freechips.rocketchip.system.DefaultRV32Config.fir@203691.10]
  wire  _T_3120; // @[TLB.scala 143:13:freechips.rocketchip.system.DefaultRV32Config.fir@203694.10]
  wire  _GEN_762; // @[TLB.scala 143:19:freechips.rocketchip.system.DefaultRV32Config.fir@203695.10]
  wire  _T_3121; // @[TLB.scala 143:13:freechips.rocketchip.system.DefaultRV32Config.fir@203698.10]
  wire  _GEN_763; // @[TLB.scala 143:19:freechips.rocketchip.system.DefaultRV32Config.fir@203699.10]
  wire  _GEN_764; // @[TLB.scala 379:40:freechips.rocketchip.system.DefaultRV32Config.fir@203537.8]
  wire  _GEN_765; // @[TLB.scala 379:40:freechips.rocketchip.system.DefaultRV32Config.fir@203537.8]
  wire  _GEN_766; // @[TLB.scala 379:40:freechips.rocketchip.system.DefaultRV32Config.fir@203537.8]
  wire  _GEN_767; // @[TLB.scala 379:40:freechips.rocketchip.system.DefaultRV32Config.fir@203537.8]
  wire  _T_3128; // @[TLB.scala 135:61:freechips.rocketchip.system.DefaultRV32Config.fir@203719.8]
  wire  _T_3273; // @[TLB.scala 143:13:freechips.rocketchip.system.DefaultRV32Config.fir@204033.10]
  wire  _GEN_788; // @[TLB.scala 143:19:freechips.rocketchip.system.DefaultRV32Config.fir@204034.10]
  wire  _T_3274; // @[TLB.scala 143:13:freechips.rocketchip.system.DefaultRV32Config.fir@204037.10]
  wire  _GEN_789; // @[TLB.scala 143:19:freechips.rocketchip.system.DefaultRV32Config.fir@204038.10]
  wire  _T_3275; // @[TLB.scala 143:13:freechips.rocketchip.system.DefaultRV32Config.fir@204041.10]
  wire  _GEN_790; // @[TLB.scala 143:19:freechips.rocketchip.system.DefaultRV32Config.fir@204042.10]
  wire  _T_3276; // @[TLB.scala 143:13:freechips.rocketchip.system.DefaultRV32Config.fir@204045.10]
  wire  _GEN_791; // @[TLB.scala 143:19:freechips.rocketchip.system.DefaultRV32Config.fir@204046.10]
  wire  _GEN_792; // @[TLB.scala 379:40:freechips.rocketchip.system.DefaultRV32Config.fir@203884.8]
  wire  _GEN_793; // @[TLB.scala 379:40:freechips.rocketchip.system.DefaultRV32Config.fir@203884.8]
  wire  _GEN_794; // @[TLB.scala 379:40:freechips.rocketchip.system.DefaultRV32Config.fir@203884.8]
  wire  _GEN_795; // @[TLB.scala 379:40:freechips.rocketchip.system.DefaultRV32Config.fir@203884.8]
  wire  _T_3283; // @[TLB.scala 135:61:freechips.rocketchip.system.DefaultRV32Config.fir@204066.8]
  wire  _T_3428; // @[TLB.scala 143:13:freechips.rocketchip.system.DefaultRV32Config.fir@204380.10]
  wire  _GEN_816; // @[TLB.scala 143:19:freechips.rocketchip.system.DefaultRV32Config.fir@204381.10]
  wire  _T_3429; // @[TLB.scala 143:13:freechips.rocketchip.system.DefaultRV32Config.fir@204384.10]
  wire  _GEN_817; // @[TLB.scala 143:19:freechips.rocketchip.system.DefaultRV32Config.fir@204385.10]
  wire  _T_3430; // @[TLB.scala 143:13:freechips.rocketchip.system.DefaultRV32Config.fir@204388.10]
  wire  _GEN_818; // @[TLB.scala 143:19:freechips.rocketchip.system.DefaultRV32Config.fir@204389.10]
  wire  _T_3431; // @[TLB.scala 143:13:freechips.rocketchip.system.DefaultRV32Config.fir@204392.10]
  wire  _GEN_819; // @[TLB.scala 143:19:freechips.rocketchip.system.DefaultRV32Config.fir@204393.10]
  wire  _GEN_820; // @[TLB.scala 379:40:freechips.rocketchip.system.DefaultRV32Config.fir@204231.8]
  wire  _GEN_821; // @[TLB.scala 379:40:freechips.rocketchip.system.DefaultRV32Config.fir@204231.8]
  wire  _GEN_822; // @[TLB.scala 379:40:freechips.rocketchip.system.DefaultRV32Config.fir@204231.8]
  wire  _GEN_823; // @[TLB.scala 379:40:freechips.rocketchip.system.DefaultRV32Config.fir@204231.8]
  wire  _T_3438; // @[TLB.scala 135:61:freechips.rocketchip.system.DefaultRV32Config.fir@204413.8]
  wire  _T_3583; // @[TLB.scala 143:13:freechips.rocketchip.system.DefaultRV32Config.fir@204727.10]
  wire  _GEN_844; // @[TLB.scala 143:19:freechips.rocketchip.system.DefaultRV32Config.fir@204728.10]
  wire  _T_3584; // @[TLB.scala 143:13:freechips.rocketchip.system.DefaultRV32Config.fir@204731.10]
  wire  _GEN_845; // @[TLB.scala 143:19:freechips.rocketchip.system.DefaultRV32Config.fir@204732.10]
  wire  _T_3585; // @[TLB.scala 143:13:freechips.rocketchip.system.DefaultRV32Config.fir@204735.10]
  wire  _GEN_846; // @[TLB.scala 143:19:freechips.rocketchip.system.DefaultRV32Config.fir@204736.10]
  wire  _T_3586; // @[TLB.scala 143:13:freechips.rocketchip.system.DefaultRV32Config.fir@204739.10]
  wire  _GEN_847; // @[TLB.scala 143:19:freechips.rocketchip.system.DefaultRV32Config.fir@204740.10]
  wire  _GEN_848; // @[TLB.scala 379:40:freechips.rocketchip.system.DefaultRV32Config.fir@204578.8]
  wire  _GEN_849; // @[TLB.scala 379:40:freechips.rocketchip.system.DefaultRV32Config.fir@204578.8]
  wire  _GEN_850; // @[TLB.scala 379:40:freechips.rocketchip.system.DefaultRV32Config.fir@204578.8]
  wire  _GEN_851; // @[TLB.scala 379:40:freechips.rocketchip.system.DefaultRV32Config.fir@204578.8]
  wire  _T_3619; // @[TLB.scala 143:13:freechips.rocketchip.system.DefaultRV32Config.fir@204808.10]
  wire  _GEN_857; // @[TLB.scala 143:19:freechips.rocketchip.system.DefaultRV32Config.fir@204809.10]
  wire  _GEN_858; // @[TLB.scala 379:40:freechips.rocketchip.system.DefaultRV32Config.fir@204770.8]
  wire  _T_3652; // @[TLB.scala 143:13:freechips.rocketchip.system.DefaultRV32Config.fir@204874.10]
  wire  _GEN_861; // @[TLB.scala 143:19:freechips.rocketchip.system.DefaultRV32Config.fir@204875.10]
  wire  _GEN_862; // @[TLB.scala 379:40:freechips.rocketchip.system.DefaultRV32Config.fir@204836.8]
  wire  _T_3685; // @[TLB.scala 143:13:freechips.rocketchip.system.DefaultRV32Config.fir@204940.10]
  wire  _GEN_865; // @[TLB.scala 143:19:freechips.rocketchip.system.DefaultRV32Config.fir@204941.10]
  wire  _GEN_866; // @[TLB.scala 379:40:freechips.rocketchip.system.DefaultRV32Config.fir@204902.8]
  wire  _T_3718; // @[TLB.scala 143:13:freechips.rocketchip.system.DefaultRV32Config.fir@205006.10]
  wire  _GEN_869; // @[TLB.scala 143:19:freechips.rocketchip.system.DefaultRV32Config.fir@205007.10]
  wire  _GEN_870; // @[TLB.scala 379:40:freechips.rocketchip.system.DefaultRV32Config.fir@204968.8]
  wire  _T_3751; // @[TLB.scala 143:13:freechips.rocketchip.system.DefaultRV32Config.fir@205072.10]
  wire  _GEN_873; // @[TLB.scala 143:19:freechips.rocketchip.system.DefaultRV32Config.fir@205073.10]
  wire  _GEN_874; // @[TLB.scala 379:40:freechips.rocketchip.system.DefaultRV32Config.fir@205034.8]
  wire  _T_3753; // @[TLB.scala 383:24:freechips.rocketchip.system.DefaultRV32Config.fir@205082.4]
  OptimizationBarrier OptimizationBarrier ( // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@198417.4]
    .io_x_ppn(OptimizationBarrier_io_x_ppn),
    .io_x_u(OptimizationBarrier_io_x_u),
    .io_x_ae(OptimizationBarrier_io_x_ae),
    .io_x_sw(OptimizationBarrier_io_x_sw),
    .io_x_sx(OptimizationBarrier_io_x_sx),
    .io_x_sr(OptimizationBarrier_io_x_sr),
    .io_x_pw(OptimizationBarrier_io_x_pw),
    .io_x_px(OptimizationBarrier_io_x_px),
    .io_x_pr(OptimizationBarrier_io_x_pr),
    .io_x_ppp(OptimizationBarrier_io_x_ppp),
    .io_x_pal(OptimizationBarrier_io_x_pal),
    .io_x_paa(OptimizationBarrier_io_x_paa),
    .io_x_eff(OptimizationBarrier_io_x_eff),
    .io_x_c(OptimizationBarrier_io_x_c),
    .io_y_ppn(OptimizationBarrier_io_y_ppn),
    .io_y_u(OptimizationBarrier_io_y_u),
    .io_y_ae(OptimizationBarrier_io_y_ae),
    .io_y_sw(OptimizationBarrier_io_y_sw),
    .io_y_sx(OptimizationBarrier_io_y_sx),
    .io_y_sr(OptimizationBarrier_io_y_sr),
    .io_y_pw(OptimizationBarrier_io_y_pw),
    .io_y_px(OptimizationBarrier_io_y_px),
    .io_y_pr(OptimizationBarrier_io_y_pr),
    .io_y_ppp(OptimizationBarrier_io_y_ppp),
    .io_y_pal(OptimizationBarrier_io_y_pal),
    .io_y_paa(OptimizationBarrier_io_y_paa),
    .io_y_eff(OptimizationBarrier_io_y_eff),
    .io_y_c(OptimizationBarrier_io_y_c)
  );
  PMPChecker pmp ( // @[TLB.scala 190:19:freechips.rocketchip.system.DefaultRV32Config.fir@198438.4]
    .io_prv(pmp_io_prv),
    .io_pmp_0_cfg_l(pmp_io_pmp_0_cfg_l),
    .io_pmp_0_cfg_a(pmp_io_pmp_0_cfg_a),
    .io_pmp_0_cfg_x(pmp_io_pmp_0_cfg_x),
    .io_pmp_0_cfg_w(pmp_io_pmp_0_cfg_w),
    .io_pmp_0_cfg_r(pmp_io_pmp_0_cfg_r),
    .io_pmp_0_addr(pmp_io_pmp_0_addr),
    .io_pmp_0_mask(pmp_io_pmp_0_mask),
    .io_pmp_1_cfg_l(pmp_io_pmp_1_cfg_l),
    .io_pmp_1_cfg_a(pmp_io_pmp_1_cfg_a),
    .io_pmp_1_cfg_x(pmp_io_pmp_1_cfg_x),
    .io_pmp_1_cfg_w(pmp_io_pmp_1_cfg_w),
    .io_pmp_1_cfg_r(pmp_io_pmp_1_cfg_r),
    .io_pmp_1_addr(pmp_io_pmp_1_addr),
    .io_pmp_1_mask(pmp_io_pmp_1_mask),
    .io_pmp_2_cfg_l(pmp_io_pmp_2_cfg_l),
    .io_pmp_2_cfg_a(pmp_io_pmp_2_cfg_a),
    .io_pmp_2_cfg_x(pmp_io_pmp_2_cfg_x),
    .io_pmp_2_cfg_w(pmp_io_pmp_2_cfg_w),
    .io_pmp_2_cfg_r(pmp_io_pmp_2_cfg_r),
    .io_pmp_2_addr(pmp_io_pmp_2_addr),
    .io_pmp_2_mask(pmp_io_pmp_2_mask),
    .io_pmp_3_cfg_l(pmp_io_pmp_3_cfg_l),
    .io_pmp_3_cfg_a(pmp_io_pmp_3_cfg_a),
    .io_pmp_3_cfg_x(pmp_io_pmp_3_cfg_x),
    .io_pmp_3_cfg_w(pmp_io_pmp_3_cfg_w),
    .io_pmp_3_cfg_r(pmp_io_pmp_3_cfg_r),
    .io_pmp_3_addr(pmp_io_pmp_3_addr),
    .io_pmp_3_mask(pmp_io_pmp_3_mask),
    .io_pmp_4_cfg_l(pmp_io_pmp_4_cfg_l),
    .io_pmp_4_cfg_a(pmp_io_pmp_4_cfg_a),
    .io_pmp_4_cfg_x(pmp_io_pmp_4_cfg_x),
    .io_pmp_4_cfg_w(pmp_io_pmp_4_cfg_w),
    .io_pmp_4_cfg_r(pmp_io_pmp_4_cfg_r),
    .io_pmp_4_addr(pmp_io_pmp_4_addr),
    .io_pmp_4_mask(pmp_io_pmp_4_mask),
    .io_pmp_5_cfg_l(pmp_io_pmp_5_cfg_l),
    .io_pmp_5_cfg_a(pmp_io_pmp_5_cfg_a),
    .io_pmp_5_cfg_x(pmp_io_pmp_5_cfg_x),
    .io_pmp_5_cfg_w(pmp_io_pmp_5_cfg_w),
    .io_pmp_5_cfg_r(pmp_io_pmp_5_cfg_r),
    .io_pmp_5_addr(pmp_io_pmp_5_addr),
    .io_pmp_5_mask(pmp_io_pmp_5_mask),
    .io_pmp_6_cfg_l(pmp_io_pmp_6_cfg_l),
    .io_pmp_6_cfg_a(pmp_io_pmp_6_cfg_a),
    .io_pmp_6_cfg_x(pmp_io_pmp_6_cfg_x),
    .io_pmp_6_cfg_w(pmp_io_pmp_6_cfg_w),
    .io_pmp_6_cfg_r(pmp_io_pmp_6_cfg_r),
    .io_pmp_6_addr(pmp_io_pmp_6_addr),
    .io_pmp_6_mask(pmp_io_pmp_6_mask),
    .io_pmp_7_cfg_l(pmp_io_pmp_7_cfg_l),
    .io_pmp_7_cfg_a(pmp_io_pmp_7_cfg_a),
    .io_pmp_7_cfg_x(pmp_io_pmp_7_cfg_x),
    .io_pmp_7_cfg_w(pmp_io_pmp_7_cfg_w),
    .io_pmp_7_cfg_r(pmp_io_pmp_7_cfg_r),
    .io_pmp_7_addr(pmp_io_pmp_7_addr),
    .io_pmp_7_mask(pmp_io_pmp_7_mask),
    .io_addr(pmp_io_addr),
    .io_r(pmp_io_r),
    .io_w(pmp_io_w),
    .io_x(pmp_io_x)
  );
  OptimizationBarrier OptimizationBarrier_1 ( // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@199139.4]
    .io_x_ppn(OptimizationBarrier_1_io_x_ppn),
    .io_x_u(OptimizationBarrier_1_io_x_u),
    .io_x_ae(OptimizationBarrier_1_io_x_ae),
    .io_x_sw(OptimizationBarrier_1_io_x_sw),
    .io_x_sx(OptimizationBarrier_1_io_x_sx),
    .io_x_sr(OptimizationBarrier_1_io_x_sr),
    .io_x_pw(OptimizationBarrier_1_io_x_pw),
    .io_x_px(OptimizationBarrier_1_io_x_px),
    .io_x_pr(OptimizationBarrier_1_io_x_pr),
    .io_x_ppp(OptimizationBarrier_1_io_x_ppp),
    .io_x_pal(OptimizationBarrier_1_io_x_pal),
    .io_x_paa(OptimizationBarrier_1_io_x_paa),
    .io_x_eff(OptimizationBarrier_1_io_x_eff),
    .io_x_c(OptimizationBarrier_1_io_x_c),
    .io_y_ppn(OptimizationBarrier_1_io_y_ppn),
    .io_y_u(OptimizationBarrier_1_io_y_u),
    .io_y_ae(OptimizationBarrier_1_io_y_ae),
    .io_y_sw(OptimizationBarrier_1_io_y_sw),
    .io_y_sx(OptimizationBarrier_1_io_y_sx),
    .io_y_sr(OptimizationBarrier_1_io_y_sr),
    .io_y_pw(OptimizationBarrier_1_io_y_pw),
    .io_y_px(OptimizationBarrier_1_io_y_px),
    .io_y_pr(OptimizationBarrier_1_io_y_pr),
    .io_y_ppp(OptimizationBarrier_1_io_y_ppp),
    .io_y_pal(OptimizationBarrier_1_io_y_pal),
    .io_y_paa(OptimizationBarrier_1_io_y_paa),
    .io_y_eff(OptimizationBarrier_1_io_y_eff),
    .io_y_c(OptimizationBarrier_1_io_y_c)
  );
  OptimizationBarrier OptimizationBarrier_2 ( // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@199182.4]
    .io_x_ppn(OptimizationBarrier_2_io_x_ppn),
    .io_x_u(OptimizationBarrier_2_io_x_u),
    .io_x_ae(OptimizationBarrier_2_io_x_ae),
    .io_x_sw(OptimizationBarrier_2_io_x_sw),
    .io_x_sx(OptimizationBarrier_2_io_x_sx),
    .io_x_sr(OptimizationBarrier_2_io_x_sr),
    .io_x_pw(OptimizationBarrier_2_io_x_pw),
    .io_x_px(OptimizationBarrier_2_io_x_px),
    .io_x_pr(OptimizationBarrier_2_io_x_pr),
    .io_x_ppp(OptimizationBarrier_2_io_x_ppp),
    .io_x_pal(OptimizationBarrier_2_io_x_pal),
    .io_x_paa(OptimizationBarrier_2_io_x_paa),
    .io_x_eff(OptimizationBarrier_2_io_x_eff),
    .io_x_c(OptimizationBarrier_2_io_x_c),
    .io_y_ppn(OptimizationBarrier_2_io_y_ppn),
    .io_y_u(OptimizationBarrier_2_io_y_u),
    .io_y_ae(OptimizationBarrier_2_io_y_ae),
    .io_y_sw(OptimizationBarrier_2_io_y_sw),
    .io_y_sx(OptimizationBarrier_2_io_y_sx),
    .io_y_sr(OptimizationBarrier_2_io_y_sr),
    .io_y_pw(OptimizationBarrier_2_io_y_pw),
    .io_y_px(OptimizationBarrier_2_io_y_px),
    .io_y_pr(OptimizationBarrier_2_io_y_pr),
    .io_y_ppp(OptimizationBarrier_2_io_y_ppp),
    .io_y_pal(OptimizationBarrier_2_io_y_pal),
    .io_y_paa(OptimizationBarrier_2_io_y_paa),
    .io_y_eff(OptimizationBarrier_2_io_y_eff),
    .io_y_c(OptimizationBarrier_2_io_y_c)
  );
  OptimizationBarrier OptimizationBarrier_3 ( // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@199225.4]
    .io_x_ppn(OptimizationBarrier_3_io_x_ppn),
    .io_x_u(OptimizationBarrier_3_io_x_u),
    .io_x_ae(OptimizationBarrier_3_io_x_ae),
    .io_x_sw(OptimizationBarrier_3_io_x_sw),
    .io_x_sx(OptimizationBarrier_3_io_x_sx),
    .io_x_sr(OptimizationBarrier_3_io_x_sr),
    .io_x_pw(OptimizationBarrier_3_io_x_pw),
    .io_x_px(OptimizationBarrier_3_io_x_px),
    .io_x_pr(OptimizationBarrier_3_io_x_pr),
    .io_x_ppp(OptimizationBarrier_3_io_x_ppp),
    .io_x_pal(OptimizationBarrier_3_io_x_pal),
    .io_x_paa(OptimizationBarrier_3_io_x_paa),
    .io_x_eff(OptimizationBarrier_3_io_x_eff),
    .io_x_c(OptimizationBarrier_3_io_x_c),
    .io_y_ppn(OptimizationBarrier_3_io_y_ppn),
    .io_y_u(OptimizationBarrier_3_io_y_u),
    .io_y_ae(OptimizationBarrier_3_io_y_ae),
    .io_y_sw(OptimizationBarrier_3_io_y_sw),
    .io_y_sx(OptimizationBarrier_3_io_y_sx),
    .io_y_sr(OptimizationBarrier_3_io_y_sr),
    .io_y_pw(OptimizationBarrier_3_io_y_pw),
    .io_y_px(OptimizationBarrier_3_io_y_px),
    .io_y_pr(OptimizationBarrier_3_io_y_pr),
    .io_y_ppp(OptimizationBarrier_3_io_y_ppp),
    .io_y_pal(OptimizationBarrier_3_io_y_pal),
    .io_y_paa(OptimizationBarrier_3_io_y_paa),
    .io_y_eff(OptimizationBarrier_3_io_y_eff),
    .io_y_c(OptimizationBarrier_3_io_y_c)
  );
  OptimizationBarrier OptimizationBarrier_4 ( // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@199268.4]
    .io_x_ppn(OptimizationBarrier_4_io_x_ppn),
    .io_x_u(OptimizationBarrier_4_io_x_u),
    .io_x_ae(OptimizationBarrier_4_io_x_ae),
    .io_x_sw(OptimizationBarrier_4_io_x_sw),
    .io_x_sx(OptimizationBarrier_4_io_x_sx),
    .io_x_sr(OptimizationBarrier_4_io_x_sr),
    .io_x_pw(OptimizationBarrier_4_io_x_pw),
    .io_x_px(OptimizationBarrier_4_io_x_px),
    .io_x_pr(OptimizationBarrier_4_io_x_pr),
    .io_x_ppp(OptimizationBarrier_4_io_x_ppp),
    .io_x_pal(OptimizationBarrier_4_io_x_pal),
    .io_x_paa(OptimizationBarrier_4_io_x_paa),
    .io_x_eff(OptimizationBarrier_4_io_x_eff),
    .io_x_c(OptimizationBarrier_4_io_x_c),
    .io_y_ppn(OptimizationBarrier_4_io_y_ppn),
    .io_y_u(OptimizationBarrier_4_io_y_u),
    .io_y_ae(OptimizationBarrier_4_io_y_ae),
    .io_y_sw(OptimizationBarrier_4_io_y_sw),
    .io_y_sx(OptimizationBarrier_4_io_y_sx),
    .io_y_sr(OptimizationBarrier_4_io_y_sr),
    .io_y_pw(OptimizationBarrier_4_io_y_pw),
    .io_y_px(OptimizationBarrier_4_io_y_px),
    .io_y_pr(OptimizationBarrier_4_io_y_pr),
    .io_y_ppp(OptimizationBarrier_4_io_y_ppp),
    .io_y_pal(OptimizationBarrier_4_io_y_pal),
    .io_y_paa(OptimizationBarrier_4_io_y_paa),
    .io_y_eff(OptimizationBarrier_4_io_y_eff),
    .io_y_c(OptimizationBarrier_4_io_y_c)
  );
  OptimizationBarrier OptimizationBarrier_5 ( // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@199311.4]
    .io_x_ppn(OptimizationBarrier_5_io_x_ppn),
    .io_x_u(OptimizationBarrier_5_io_x_u),
    .io_x_ae(OptimizationBarrier_5_io_x_ae),
    .io_x_sw(OptimizationBarrier_5_io_x_sw),
    .io_x_sx(OptimizationBarrier_5_io_x_sx),
    .io_x_sr(OptimizationBarrier_5_io_x_sr),
    .io_x_pw(OptimizationBarrier_5_io_x_pw),
    .io_x_px(OptimizationBarrier_5_io_x_px),
    .io_x_pr(OptimizationBarrier_5_io_x_pr),
    .io_x_ppp(OptimizationBarrier_5_io_x_ppp),
    .io_x_pal(OptimizationBarrier_5_io_x_pal),
    .io_x_paa(OptimizationBarrier_5_io_x_paa),
    .io_x_eff(OptimizationBarrier_5_io_x_eff),
    .io_x_c(OptimizationBarrier_5_io_x_c),
    .io_y_ppn(OptimizationBarrier_5_io_y_ppn),
    .io_y_u(OptimizationBarrier_5_io_y_u),
    .io_y_ae(OptimizationBarrier_5_io_y_ae),
    .io_y_sw(OptimizationBarrier_5_io_y_sw),
    .io_y_sx(OptimizationBarrier_5_io_y_sx),
    .io_y_sr(OptimizationBarrier_5_io_y_sr),
    .io_y_pw(OptimizationBarrier_5_io_y_pw),
    .io_y_px(OptimizationBarrier_5_io_y_px),
    .io_y_pr(OptimizationBarrier_5_io_y_pr),
    .io_y_ppp(OptimizationBarrier_5_io_y_ppp),
    .io_y_pal(OptimizationBarrier_5_io_y_pal),
    .io_y_paa(OptimizationBarrier_5_io_y_paa),
    .io_y_eff(OptimizationBarrier_5_io_y_eff),
    .io_y_c(OptimizationBarrier_5_io_y_c)
  );
  OptimizationBarrier OptimizationBarrier_6 ( // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@199354.4]
    .io_x_ppn(OptimizationBarrier_6_io_x_ppn),
    .io_x_u(OptimizationBarrier_6_io_x_u),
    .io_x_ae(OptimizationBarrier_6_io_x_ae),
    .io_x_sw(OptimizationBarrier_6_io_x_sw),
    .io_x_sx(OptimizationBarrier_6_io_x_sx),
    .io_x_sr(OptimizationBarrier_6_io_x_sr),
    .io_x_pw(OptimizationBarrier_6_io_x_pw),
    .io_x_px(OptimizationBarrier_6_io_x_px),
    .io_x_pr(OptimizationBarrier_6_io_x_pr),
    .io_x_ppp(OptimizationBarrier_6_io_x_ppp),
    .io_x_pal(OptimizationBarrier_6_io_x_pal),
    .io_x_paa(OptimizationBarrier_6_io_x_paa),
    .io_x_eff(OptimizationBarrier_6_io_x_eff),
    .io_x_c(OptimizationBarrier_6_io_x_c),
    .io_y_ppn(OptimizationBarrier_6_io_y_ppn),
    .io_y_u(OptimizationBarrier_6_io_y_u),
    .io_y_ae(OptimizationBarrier_6_io_y_ae),
    .io_y_sw(OptimizationBarrier_6_io_y_sw),
    .io_y_sx(OptimizationBarrier_6_io_y_sx),
    .io_y_sr(OptimizationBarrier_6_io_y_sr),
    .io_y_pw(OptimizationBarrier_6_io_y_pw),
    .io_y_px(OptimizationBarrier_6_io_y_px),
    .io_y_pr(OptimizationBarrier_6_io_y_pr),
    .io_y_ppp(OptimizationBarrier_6_io_y_ppp),
    .io_y_pal(OptimizationBarrier_6_io_y_pal),
    .io_y_paa(OptimizationBarrier_6_io_y_paa),
    .io_y_eff(OptimizationBarrier_6_io_y_eff),
    .io_y_c(OptimizationBarrier_6_io_y_c)
  );
  OptimizationBarrier OptimizationBarrier_7 ( // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@199397.4]
    .io_x_ppn(OptimizationBarrier_7_io_x_ppn),
    .io_x_u(OptimizationBarrier_7_io_x_u),
    .io_x_ae(OptimizationBarrier_7_io_x_ae),
    .io_x_sw(OptimizationBarrier_7_io_x_sw),
    .io_x_sx(OptimizationBarrier_7_io_x_sx),
    .io_x_sr(OptimizationBarrier_7_io_x_sr),
    .io_x_pw(OptimizationBarrier_7_io_x_pw),
    .io_x_px(OptimizationBarrier_7_io_x_px),
    .io_x_pr(OptimizationBarrier_7_io_x_pr),
    .io_x_ppp(OptimizationBarrier_7_io_x_ppp),
    .io_x_pal(OptimizationBarrier_7_io_x_pal),
    .io_x_paa(OptimizationBarrier_7_io_x_paa),
    .io_x_eff(OptimizationBarrier_7_io_x_eff),
    .io_x_c(OptimizationBarrier_7_io_x_c),
    .io_y_ppn(OptimizationBarrier_7_io_y_ppn),
    .io_y_u(OptimizationBarrier_7_io_y_u),
    .io_y_ae(OptimizationBarrier_7_io_y_ae),
    .io_y_sw(OptimizationBarrier_7_io_y_sw),
    .io_y_sx(OptimizationBarrier_7_io_y_sx),
    .io_y_sr(OptimizationBarrier_7_io_y_sr),
    .io_y_pw(OptimizationBarrier_7_io_y_pw),
    .io_y_px(OptimizationBarrier_7_io_y_px),
    .io_y_pr(OptimizationBarrier_7_io_y_pr),
    .io_y_ppp(OptimizationBarrier_7_io_y_ppp),
    .io_y_pal(OptimizationBarrier_7_io_y_pal),
    .io_y_paa(OptimizationBarrier_7_io_y_paa),
    .io_y_eff(OptimizationBarrier_7_io_y_eff),
    .io_y_c(OptimizationBarrier_7_io_y_c)
  );
  OptimizationBarrier OptimizationBarrier_8 ( // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@199440.4]
    .io_x_ppn(OptimizationBarrier_8_io_x_ppn),
    .io_x_u(OptimizationBarrier_8_io_x_u),
    .io_x_ae(OptimizationBarrier_8_io_x_ae),
    .io_x_sw(OptimizationBarrier_8_io_x_sw),
    .io_x_sx(OptimizationBarrier_8_io_x_sx),
    .io_x_sr(OptimizationBarrier_8_io_x_sr),
    .io_x_pw(OptimizationBarrier_8_io_x_pw),
    .io_x_px(OptimizationBarrier_8_io_x_px),
    .io_x_pr(OptimizationBarrier_8_io_x_pr),
    .io_x_ppp(OptimizationBarrier_8_io_x_ppp),
    .io_x_pal(OptimizationBarrier_8_io_x_pal),
    .io_x_paa(OptimizationBarrier_8_io_x_paa),
    .io_x_eff(OptimizationBarrier_8_io_x_eff),
    .io_x_c(OptimizationBarrier_8_io_x_c),
    .io_y_ppn(OptimizationBarrier_8_io_y_ppn),
    .io_y_u(OptimizationBarrier_8_io_y_u),
    .io_y_ae(OptimizationBarrier_8_io_y_ae),
    .io_y_sw(OptimizationBarrier_8_io_y_sw),
    .io_y_sx(OptimizationBarrier_8_io_y_sx),
    .io_y_sr(OptimizationBarrier_8_io_y_sr),
    .io_y_pw(OptimizationBarrier_8_io_y_pw),
    .io_y_px(OptimizationBarrier_8_io_y_px),
    .io_y_pr(OptimizationBarrier_8_io_y_pr),
    .io_y_ppp(OptimizationBarrier_8_io_y_ppp),
    .io_y_pal(OptimizationBarrier_8_io_y_pal),
    .io_y_paa(OptimizationBarrier_8_io_y_paa),
    .io_y_eff(OptimizationBarrier_8_io_y_eff),
    .io_y_c(OptimizationBarrier_8_io_y_c)
  );
  OptimizationBarrier OptimizationBarrier_9 ( // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@199482.4]
    .io_x_ppn(OptimizationBarrier_9_io_x_ppn),
    .io_x_u(OptimizationBarrier_9_io_x_u),
    .io_x_ae(OptimizationBarrier_9_io_x_ae),
    .io_x_sw(OptimizationBarrier_9_io_x_sw),
    .io_x_sx(OptimizationBarrier_9_io_x_sx),
    .io_x_sr(OptimizationBarrier_9_io_x_sr),
    .io_x_pw(OptimizationBarrier_9_io_x_pw),
    .io_x_px(OptimizationBarrier_9_io_x_px),
    .io_x_pr(OptimizationBarrier_9_io_x_pr),
    .io_x_ppp(OptimizationBarrier_9_io_x_ppp),
    .io_x_pal(OptimizationBarrier_9_io_x_pal),
    .io_x_paa(OptimizationBarrier_9_io_x_paa),
    .io_x_eff(OptimizationBarrier_9_io_x_eff),
    .io_x_c(OptimizationBarrier_9_io_x_c),
    .io_y_ppn(OptimizationBarrier_9_io_y_ppn),
    .io_y_u(OptimizationBarrier_9_io_y_u),
    .io_y_ae(OptimizationBarrier_9_io_y_ae),
    .io_y_sw(OptimizationBarrier_9_io_y_sw),
    .io_y_sx(OptimizationBarrier_9_io_y_sx),
    .io_y_sr(OptimizationBarrier_9_io_y_sr),
    .io_y_pw(OptimizationBarrier_9_io_y_pw),
    .io_y_px(OptimizationBarrier_9_io_y_px),
    .io_y_pr(OptimizationBarrier_9_io_y_pr),
    .io_y_ppp(OptimizationBarrier_9_io_y_ppp),
    .io_y_pal(OptimizationBarrier_9_io_y_pal),
    .io_y_paa(OptimizationBarrier_9_io_y_paa),
    .io_y_eff(OptimizationBarrier_9_io_y_eff),
    .io_y_c(OptimizationBarrier_9_io_y_c)
  );
  OptimizationBarrier OptimizationBarrier_10 ( // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@199531.4]
    .io_x_ppn(OptimizationBarrier_10_io_x_ppn),
    .io_x_u(OptimizationBarrier_10_io_x_u),
    .io_x_ae(OptimizationBarrier_10_io_x_ae),
    .io_x_sw(OptimizationBarrier_10_io_x_sw),
    .io_x_sx(OptimizationBarrier_10_io_x_sx),
    .io_x_sr(OptimizationBarrier_10_io_x_sr),
    .io_x_pw(OptimizationBarrier_10_io_x_pw),
    .io_x_px(OptimizationBarrier_10_io_x_px),
    .io_x_pr(OptimizationBarrier_10_io_x_pr),
    .io_x_ppp(OptimizationBarrier_10_io_x_ppp),
    .io_x_pal(OptimizationBarrier_10_io_x_pal),
    .io_x_paa(OptimizationBarrier_10_io_x_paa),
    .io_x_eff(OptimizationBarrier_10_io_x_eff),
    .io_x_c(OptimizationBarrier_10_io_x_c),
    .io_y_ppn(OptimizationBarrier_10_io_y_ppn),
    .io_y_u(OptimizationBarrier_10_io_y_u),
    .io_y_ae(OptimizationBarrier_10_io_y_ae),
    .io_y_sw(OptimizationBarrier_10_io_y_sw),
    .io_y_sx(OptimizationBarrier_10_io_y_sx),
    .io_y_sr(OptimizationBarrier_10_io_y_sr),
    .io_y_pw(OptimizationBarrier_10_io_y_pw),
    .io_y_px(OptimizationBarrier_10_io_y_px),
    .io_y_pr(OptimizationBarrier_10_io_y_pr),
    .io_y_ppp(OptimizationBarrier_10_io_y_ppp),
    .io_y_pal(OptimizationBarrier_10_io_y_pal),
    .io_y_paa(OptimizationBarrier_10_io_y_paa),
    .io_y_eff(OptimizationBarrier_10_io_y_eff),
    .io_y_c(OptimizationBarrier_10_io_y_c)
  );
  OptimizationBarrier OptimizationBarrier_11 ( // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@199580.4]
    .io_x_ppn(OptimizationBarrier_11_io_x_ppn),
    .io_x_u(OptimizationBarrier_11_io_x_u),
    .io_x_ae(OptimizationBarrier_11_io_x_ae),
    .io_x_sw(OptimizationBarrier_11_io_x_sw),
    .io_x_sx(OptimizationBarrier_11_io_x_sx),
    .io_x_sr(OptimizationBarrier_11_io_x_sr),
    .io_x_pw(OptimizationBarrier_11_io_x_pw),
    .io_x_px(OptimizationBarrier_11_io_x_px),
    .io_x_pr(OptimizationBarrier_11_io_x_pr),
    .io_x_ppp(OptimizationBarrier_11_io_x_ppp),
    .io_x_pal(OptimizationBarrier_11_io_x_pal),
    .io_x_paa(OptimizationBarrier_11_io_x_paa),
    .io_x_eff(OptimizationBarrier_11_io_x_eff),
    .io_x_c(OptimizationBarrier_11_io_x_c),
    .io_y_ppn(OptimizationBarrier_11_io_y_ppn),
    .io_y_u(OptimizationBarrier_11_io_y_u),
    .io_y_ae(OptimizationBarrier_11_io_y_ae),
    .io_y_sw(OptimizationBarrier_11_io_y_sw),
    .io_y_sx(OptimizationBarrier_11_io_y_sx),
    .io_y_sr(OptimizationBarrier_11_io_y_sr),
    .io_y_pw(OptimizationBarrier_11_io_y_pw),
    .io_y_px(OptimizationBarrier_11_io_y_px),
    .io_y_pr(OptimizationBarrier_11_io_y_pr),
    .io_y_ppp(OptimizationBarrier_11_io_y_ppp),
    .io_y_pal(OptimizationBarrier_11_io_y_pal),
    .io_y_paa(OptimizationBarrier_11_io_y_paa),
    .io_y_eff(OptimizationBarrier_11_io_y_eff),
    .io_y_c(OptimizationBarrier_11_io_y_c)
  );
  OptimizationBarrier OptimizationBarrier_12 ( // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@199629.4]
    .io_x_ppn(OptimizationBarrier_12_io_x_ppn),
    .io_x_u(OptimizationBarrier_12_io_x_u),
    .io_x_ae(OptimizationBarrier_12_io_x_ae),
    .io_x_sw(OptimizationBarrier_12_io_x_sw),
    .io_x_sx(OptimizationBarrier_12_io_x_sx),
    .io_x_sr(OptimizationBarrier_12_io_x_sr),
    .io_x_pw(OptimizationBarrier_12_io_x_pw),
    .io_x_px(OptimizationBarrier_12_io_x_px),
    .io_x_pr(OptimizationBarrier_12_io_x_pr),
    .io_x_ppp(OptimizationBarrier_12_io_x_ppp),
    .io_x_pal(OptimizationBarrier_12_io_x_pal),
    .io_x_paa(OptimizationBarrier_12_io_x_paa),
    .io_x_eff(OptimizationBarrier_12_io_x_eff),
    .io_x_c(OptimizationBarrier_12_io_x_c),
    .io_y_ppn(OptimizationBarrier_12_io_y_ppn),
    .io_y_u(OptimizationBarrier_12_io_y_u),
    .io_y_ae(OptimizationBarrier_12_io_y_ae),
    .io_y_sw(OptimizationBarrier_12_io_y_sw),
    .io_y_sx(OptimizationBarrier_12_io_y_sx),
    .io_y_sr(OptimizationBarrier_12_io_y_sr),
    .io_y_pw(OptimizationBarrier_12_io_y_pw),
    .io_y_px(OptimizationBarrier_12_io_y_px),
    .io_y_pr(OptimizationBarrier_12_io_y_pr),
    .io_y_ppp(OptimizationBarrier_12_io_y_ppp),
    .io_y_pal(OptimizationBarrier_12_io_y_pal),
    .io_y_paa(OptimizationBarrier_12_io_y_paa),
    .io_y_eff(OptimizationBarrier_12_io_y_eff),
    .io_y_c(OptimizationBarrier_12_io_y_c)
  );
  OptimizationBarrier OptimizationBarrier_13 ( // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@199678.4]
    .io_x_ppn(OptimizationBarrier_13_io_x_ppn),
    .io_x_u(OptimizationBarrier_13_io_x_u),
    .io_x_ae(OptimizationBarrier_13_io_x_ae),
    .io_x_sw(OptimizationBarrier_13_io_x_sw),
    .io_x_sx(OptimizationBarrier_13_io_x_sx),
    .io_x_sr(OptimizationBarrier_13_io_x_sr),
    .io_x_pw(OptimizationBarrier_13_io_x_pw),
    .io_x_px(OptimizationBarrier_13_io_x_px),
    .io_x_pr(OptimizationBarrier_13_io_x_pr),
    .io_x_ppp(OptimizationBarrier_13_io_x_ppp),
    .io_x_pal(OptimizationBarrier_13_io_x_pal),
    .io_x_paa(OptimizationBarrier_13_io_x_paa),
    .io_x_eff(OptimizationBarrier_13_io_x_eff),
    .io_x_c(OptimizationBarrier_13_io_x_c),
    .io_y_ppn(OptimizationBarrier_13_io_y_ppn),
    .io_y_u(OptimizationBarrier_13_io_y_u),
    .io_y_ae(OptimizationBarrier_13_io_y_ae),
    .io_y_sw(OptimizationBarrier_13_io_y_sw),
    .io_y_sx(OptimizationBarrier_13_io_y_sx),
    .io_y_sr(OptimizationBarrier_13_io_y_sr),
    .io_y_pw(OptimizationBarrier_13_io_y_pw),
    .io_y_px(OptimizationBarrier_13_io_y_px),
    .io_y_pr(OptimizationBarrier_13_io_y_pr),
    .io_y_ppp(OptimizationBarrier_13_io_y_ppp),
    .io_y_pal(OptimizationBarrier_13_io_y_pal),
    .io_y_paa(OptimizationBarrier_13_io_y_paa),
    .io_y_eff(OptimizationBarrier_13_io_y_eff),
    .io_y_c(OptimizationBarrier_13_io_y_c)
  );
  OptimizationBarrier OptimizationBarrier_14 ( // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@200159.4]
    .io_x_ppn(OptimizationBarrier_14_io_x_ppn),
    .io_x_u(OptimizationBarrier_14_io_x_u),
    .io_x_ae(OptimizationBarrier_14_io_x_ae),
    .io_x_sw(OptimizationBarrier_14_io_x_sw),
    .io_x_sx(OptimizationBarrier_14_io_x_sx),
    .io_x_sr(OptimizationBarrier_14_io_x_sr),
    .io_x_pw(OptimizationBarrier_14_io_x_pw),
    .io_x_px(OptimizationBarrier_14_io_x_px),
    .io_x_pr(OptimizationBarrier_14_io_x_pr),
    .io_x_ppp(OptimizationBarrier_14_io_x_ppp),
    .io_x_pal(OptimizationBarrier_14_io_x_pal),
    .io_x_paa(OptimizationBarrier_14_io_x_paa),
    .io_x_eff(OptimizationBarrier_14_io_x_eff),
    .io_x_c(OptimizationBarrier_14_io_x_c),
    .io_y_ppn(OptimizationBarrier_14_io_y_ppn),
    .io_y_u(OptimizationBarrier_14_io_y_u),
    .io_y_ae(OptimizationBarrier_14_io_y_ae),
    .io_y_sw(OptimizationBarrier_14_io_y_sw),
    .io_y_sx(OptimizationBarrier_14_io_y_sx),
    .io_y_sr(OptimizationBarrier_14_io_y_sr),
    .io_y_pw(OptimizationBarrier_14_io_y_pw),
    .io_y_px(OptimizationBarrier_14_io_y_px),
    .io_y_pr(OptimizationBarrier_14_io_y_pr),
    .io_y_ppp(OptimizationBarrier_14_io_y_ppp),
    .io_y_pal(OptimizationBarrier_14_io_y_pal),
    .io_y_paa(OptimizationBarrier_14_io_y_paa),
    .io_y_eff(OptimizationBarrier_14_io_y_eff),
    .io_y_c(OptimizationBarrier_14_io_y_c)
  );
  OptimizationBarrier OptimizationBarrier_15 ( // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@200202.4]
    .io_x_ppn(OptimizationBarrier_15_io_x_ppn),
    .io_x_u(OptimizationBarrier_15_io_x_u),
    .io_x_ae(OptimizationBarrier_15_io_x_ae),
    .io_x_sw(OptimizationBarrier_15_io_x_sw),
    .io_x_sx(OptimizationBarrier_15_io_x_sx),
    .io_x_sr(OptimizationBarrier_15_io_x_sr),
    .io_x_pw(OptimizationBarrier_15_io_x_pw),
    .io_x_px(OptimizationBarrier_15_io_x_px),
    .io_x_pr(OptimizationBarrier_15_io_x_pr),
    .io_x_ppp(OptimizationBarrier_15_io_x_ppp),
    .io_x_pal(OptimizationBarrier_15_io_x_pal),
    .io_x_paa(OptimizationBarrier_15_io_x_paa),
    .io_x_eff(OptimizationBarrier_15_io_x_eff),
    .io_x_c(OptimizationBarrier_15_io_x_c),
    .io_y_ppn(OptimizationBarrier_15_io_y_ppn),
    .io_y_u(OptimizationBarrier_15_io_y_u),
    .io_y_ae(OptimizationBarrier_15_io_y_ae),
    .io_y_sw(OptimizationBarrier_15_io_y_sw),
    .io_y_sx(OptimizationBarrier_15_io_y_sx),
    .io_y_sr(OptimizationBarrier_15_io_y_sr),
    .io_y_pw(OptimizationBarrier_15_io_y_pw),
    .io_y_px(OptimizationBarrier_15_io_y_px),
    .io_y_pr(OptimizationBarrier_15_io_y_pr),
    .io_y_ppp(OptimizationBarrier_15_io_y_ppp),
    .io_y_pal(OptimizationBarrier_15_io_y_pal),
    .io_y_paa(OptimizationBarrier_15_io_y_paa),
    .io_y_eff(OptimizationBarrier_15_io_y_eff),
    .io_y_c(OptimizationBarrier_15_io_y_c)
  );
  OptimizationBarrier OptimizationBarrier_16 ( // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@200245.4]
    .io_x_ppn(OptimizationBarrier_16_io_x_ppn),
    .io_x_u(OptimizationBarrier_16_io_x_u),
    .io_x_ae(OptimizationBarrier_16_io_x_ae),
    .io_x_sw(OptimizationBarrier_16_io_x_sw),
    .io_x_sx(OptimizationBarrier_16_io_x_sx),
    .io_x_sr(OptimizationBarrier_16_io_x_sr),
    .io_x_pw(OptimizationBarrier_16_io_x_pw),
    .io_x_px(OptimizationBarrier_16_io_x_px),
    .io_x_pr(OptimizationBarrier_16_io_x_pr),
    .io_x_ppp(OptimizationBarrier_16_io_x_ppp),
    .io_x_pal(OptimizationBarrier_16_io_x_pal),
    .io_x_paa(OptimizationBarrier_16_io_x_paa),
    .io_x_eff(OptimizationBarrier_16_io_x_eff),
    .io_x_c(OptimizationBarrier_16_io_x_c),
    .io_y_ppn(OptimizationBarrier_16_io_y_ppn),
    .io_y_u(OptimizationBarrier_16_io_y_u),
    .io_y_ae(OptimizationBarrier_16_io_y_ae),
    .io_y_sw(OptimizationBarrier_16_io_y_sw),
    .io_y_sx(OptimizationBarrier_16_io_y_sx),
    .io_y_sr(OptimizationBarrier_16_io_y_sr),
    .io_y_pw(OptimizationBarrier_16_io_y_pw),
    .io_y_px(OptimizationBarrier_16_io_y_px),
    .io_y_pr(OptimizationBarrier_16_io_y_pr),
    .io_y_ppp(OptimizationBarrier_16_io_y_ppp),
    .io_y_pal(OptimizationBarrier_16_io_y_pal),
    .io_y_paa(OptimizationBarrier_16_io_y_paa),
    .io_y_eff(OptimizationBarrier_16_io_y_eff),
    .io_y_c(OptimizationBarrier_16_io_y_c)
  );
  OptimizationBarrier OptimizationBarrier_17 ( // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@200288.4]
    .io_x_ppn(OptimizationBarrier_17_io_x_ppn),
    .io_x_u(OptimizationBarrier_17_io_x_u),
    .io_x_ae(OptimizationBarrier_17_io_x_ae),
    .io_x_sw(OptimizationBarrier_17_io_x_sw),
    .io_x_sx(OptimizationBarrier_17_io_x_sx),
    .io_x_sr(OptimizationBarrier_17_io_x_sr),
    .io_x_pw(OptimizationBarrier_17_io_x_pw),
    .io_x_px(OptimizationBarrier_17_io_x_px),
    .io_x_pr(OptimizationBarrier_17_io_x_pr),
    .io_x_ppp(OptimizationBarrier_17_io_x_ppp),
    .io_x_pal(OptimizationBarrier_17_io_x_pal),
    .io_x_paa(OptimizationBarrier_17_io_x_paa),
    .io_x_eff(OptimizationBarrier_17_io_x_eff),
    .io_x_c(OptimizationBarrier_17_io_x_c),
    .io_y_ppn(OptimizationBarrier_17_io_y_ppn),
    .io_y_u(OptimizationBarrier_17_io_y_u),
    .io_y_ae(OptimizationBarrier_17_io_y_ae),
    .io_y_sw(OptimizationBarrier_17_io_y_sw),
    .io_y_sx(OptimizationBarrier_17_io_y_sx),
    .io_y_sr(OptimizationBarrier_17_io_y_sr),
    .io_y_pw(OptimizationBarrier_17_io_y_pw),
    .io_y_px(OptimizationBarrier_17_io_y_px),
    .io_y_pr(OptimizationBarrier_17_io_y_pr),
    .io_y_ppp(OptimizationBarrier_17_io_y_ppp),
    .io_y_pal(OptimizationBarrier_17_io_y_pal),
    .io_y_paa(OptimizationBarrier_17_io_y_paa),
    .io_y_eff(OptimizationBarrier_17_io_y_eff),
    .io_y_c(OptimizationBarrier_17_io_y_c)
  );
  OptimizationBarrier OptimizationBarrier_18 ( // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@200331.4]
    .io_x_ppn(OptimizationBarrier_18_io_x_ppn),
    .io_x_u(OptimizationBarrier_18_io_x_u),
    .io_x_ae(OptimizationBarrier_18_io_x_ae),
    .io_x_sw(OptimizationBarrier_18_io_x_sw),
    .io_x_sx(OptimizationBarrier_18_io_x_sx),
    .io_x_sr(OptimizationBarrier_18_io_x_sr),
    .io_x_pw(OptimizationBarrier_18_io_x_pw),
    .io_x_px(OptimizationBarrier_18_io_x_px),
    .io_x_pr(OptimizationBarrier_18_io_x_pr),
    .io_x_ppp(OptimizationBarrier_18_io_x_ppp),
    .io_x_pal(OptimizationBarrier_18_io_x_pal),
    .io_x_paa(OptimizationBarrier_18_io_x_paa),
    .io_x_eff(OptimizationBarrier_18_io_x_eff),
    .io_x_c(OptimizationBarrier_18_io_x_c),
    .io_y_ppn(OptimizationBarrier_18_io_y_ppn),
    .io_y_u(OptimizationBarrier_18_io_y_u),
    .io_y_ae(OptimizationBarrier_18_io_y_ae),
    .io_y_sw(OptimizationBarrier_18_io_y_sw),
    .io_y_sx(OptimizationBarrier_18_io_y_sx),
    .io_y_sr(OptimizationBarrier_18_io_y_sr),
    .io_y_pw(OptimizationBarrier_18_io_y_pw),
    .io_y_px(OptimizationBarrier_18_io_y_px),
    .io_y_pr(OptimizationBarrier_18_io_y_pr),
    .io_y_ppp(OptimizationBarrier_18_io_y_ppp),
    .io_y_pal(OptimizationBarrier_18_io_y_pal),
    .io_y_paa(OptimizationBarrier_18_io_y_paa),
    .io_y_eff(OptimizationBarrier_18_io_y_eff),
    .io_y_c(OptimizationBarrier_18_io_y_c)
  );
  OptimizationBarrier OptimizationBarrier_19 ( // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@200374.4]
    .io_x_ppn(OptimizationBarrier_19_io_x_ppn),
    .io_x_u(OptimizationBarrier_19_io_x_u),
    .io_x_ae(OptimizationBarrier_19_io_x_ae),
    .io_x_sw(OptimizationBarrier_19_io_x_sw),
    .io_x_sx(OptimizationBarrier_19_io_x_sx),
    .io_x_sr(OptimizationBarrier_19_io_x_sr),
    .io_x_pw(OptimizationBarrier_19_io_x_pw),
    .io_x_px(OptimizationBarrier_19_io_x_px),
    .io_x_pr(OptimizationBarrier_19_io_x_pr),
    .io_x_ppp(OptimizationBarrier_19_io_x_ppp),
    .io_x_pal(OptimizationBarrier_19_io_x_pal),
    .io_x_paa(OptimizationBarrier_19_io_x_paa),
    .io_x_eff(OptimizationBarrier_19_io_x_eff),
    .io_x_c(OptimizationBarrier_19_io_x_c),
    .io_y_ppn(OptimizationBarrier_19_io_y_ppn),
    .io_y_u(OptimizationBarrier_19_io_y_u),
    .io_y_ae(OptimizationBarrier_19_io_y_ae),
    .io_y_sw(OptimizationBarrier_19_io_y_sw),
    .io_y_sx(OptimizationBarrier_19_io_y_sx),
    .io_y_sr(OptimizationBarrier_19_io_y_sr),
    .io_y_pw(OptimizationBarrier_19_io_y_pw),
    .io_y_px(OptimizationBarrier_19_io_y_px),
    .io_y_pr(OptimizationBarrier_19_io_y_pr),
    .io_y_ppp(OptimizationBarrier_19_io_y_ppp),
    .io_y_pal(OptimizationBarrier_19_io_y_pal),
    .io_y_paa(OptimizationBarrier_19_io_y_paa),
    .io_y_eff(OptimizationBarrier_19_io_y_eff),
    .io_y_c(OptimizationBarrier_19_io_y_c)
  );
  OptimizationBarrier OptimizationBarrier_20 ( // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@200417.4]
    .io_x_ppn(OptimizationBarrier_20_io_x_ppn),
    .io_x_u(OptimizationBarrier_20_io_x_u),
    .io_x_ae(OptimizationBarrier_20_io_x_ae),
    .io_x_sw(OptimizationBarrier_20_io_x_sw),
    .io_x_sx(OptimizationBarrier_20_io_x_sx),
    .io_x_sr(OptimizationBarrier_20_io_x_sr),
    .io_x_pw(OptimizationBarrier_20_io_x_pw),
    .io_x_px(OptimizationBarrier_20_io_x_px),
    .io_x_pr(OptimizationBarrier_20_io_x_pr),
    .io_x_ppp(OptimizationBarrier_20_io_x_ppp),
    .io_x_pal(OptimizationBarrier_20_io_x_pal),
    .io_x_paa(OptimizationBarrier_20_io_x_paa),
    .io_x_eff(OptimizationBarrier_20_io_x_eff),
    .io_x_c(OptimizationBarrier_20_io_x_c),
    .io_y_ppn(OptimizationBarrier_20_io_y_ppn),
    .io_y_u(OptimizationBarrier_20_io_y_u),
    .io_y_ae(OptimizationBarrier_20_io_y_ae),
    .io_y_sw(OptimizationBarrier_20_io_y_sw),
    .io_y_sx(OptimizationBarrier_20_io_y_sx),
    .io_y_sr(OptimizationBarrier_20_io_y_sr),
    .io_y_pw(OptimizationBarrier_20_io_y_pw),
    .io_y_px(OptimizationBarrier_20_io_y_px),
    .io_y_pr(OptimizationBarrier_20_io_y_pr),
    .io_y_ppp(OptimizationBarrier_20_io_y_ppp),
    .io_y_pal(OptimizationBarrier_20_io_y_pal),
    .io_y_paa(OptimizationBarrier_20_io_y_paa),
    .io_y_eff(OptimizationBarrier_20_io_y_eff),
    .io_y_c(OptimizationBarrier_20_io_y_c)
  );
  OptimizationBarrier OptimizationBarrier_21 ( // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@200460.4]
    .io_x_ppn(OptimizationBarrier_21_io_x_ppn),
    .io_x_u(OptimizationBarrier_21_io_x_u),
    .io_x_ae(OptimizationBarrier_21_io_x_ae),
    .io_x_sw(OptimizationBarrier_21_io_x_sw),
    .io_x_sx(OptimizationBarrier_21_io_x_sx),
    .io_x_sr(OptimizationBarrier_21_io_x_sr),
    .io_x_pw(OptimizationBarrier_21_io_x_pw),
    .io_x_px(OptimizationBarrier_21_io_x_px),
    .io_x_pr(OptimizationBarrier_21_io_x_pr),
    .io_x_ppp(OptimizationBarrier_21_io_x_ppp),
    .io_x_pal(OptimizationBarrier_21_io_x_pal),
    .io_x_paa(OptimizationBarrier_21_io_x_paa),
    .io_x_eff(OptimizationBarrier_21_io_x_eff),
    .io_x_c(OptimizationBarrier_21_io_x_c),
    .io_y_ppn(OptimizationBarrier_21_io_y_ppn),
    .io_y_u(OptimizationBarrier_21_io_y_u),
    .io_y_ae(OptimizationBarrier_21_io_y_ae),
    .io_y_sw(OptimizationBarrier_21_io_y_sw),
    .io_y_sx(OptimizationBarrier_21_io_y_sx),
    .io_y_sr(OptimizationBarrier_21_io_y_sr),
    .io_y_pw(OptimizationBarrier_21_io_y_pw),
    .io_y_px(OptimizationBarrier_21_io_y_px),
    .io_y_pr(OptimizationBarrier_21_io_y_pr),
    .io_y_ppp(OptimizationBarrier_21_io_y_ppp),
    .io_y_pal(OptimizationBarrier_21_io_y_pal),
    .io_y_paa(OptimizationBarrier_21_io_y_paa),
    .io_y_eff(OptimizationBarrier_21_io_y_eff),
    .io_y_c(OptimizationBarrier_21_io_y_c)
  );
  OptimizationBarrier OptimizationBarrier_22 ( // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@200502.4]
    .io_x_ppn(OptimizationBarrier_22_io_x_ppn),
    .io_x_u(OptimizationBarrier_22_io_x_u),
    .io_x_ae(OptimizationBarrier_22_io_x_ae),
    .io_x_sw(OptimizationBarrier_22_io_x_sw),
    .io_x_sx(OptimizationBarrier_22_io_x_sx),
    .io_x_sr(OptimizationBarrier_22_io_x_sr),
    .io_x_pw(OptimizationBarrier_22_io_x_pw),
    .io_x_px(OptimizationBarrier_22_io_x_px),
    .io_x_pr(OptimizationBarrier_22_io_x_pr),
    .io_x_ppp(OptimizationBarrier_22_io_x_ppp),
    .io_x_pal(OptimizationBarrier_22_io_x_pal),
    .io_x_paa(OptimizationBarrier_22_io_x_paa),
    .io_x_eff(OptimizationBarrier_22_io_x_eff),
    .io_x_c(OptimizationBarrier_22_io_x_c),
    .io_y_ppn(OptimizationBarrier_22_io_y_ppn),
    .io_y_u(OptimizationBarrier_22_io_y_u),
    .io_y_ae(OptimizationBarrier_22_io_y_ae),
    .io_y_sw(OptimizationBarrier_22_io_y_sw),
    .io_y_sx(OptimizationBarrier_22_io_y_sx),
    .io_y_sr(OptimizationBarrier_22_io_y_sr),
    .io_y_pw(OptimizationBarrier_22_io_y_pw),
    .io_y_px(OptimizationBarrier_22_io_y_px),
    .io_y_pr(OptimizationBarrier_22_io_y_pr),
    .io_y_ppp(OptimizationBarrier_22_io_y_ppp),
    .io_y_pal(OptimizationBarrier_22_io_y_pal),
    .io_y_paa(OptimizationBarrier_22_io_y_paa),
    .io_y_eff(OptimizationBarrier_22_io_y_eff),
    .io_y_c(OptimizationBarrier_22_io_y_c)
  );
  OptimizationBarrier OptimizationBarrier_23 ( // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@200544.4]
    .io_x_ppn(OptimizationBarrier_23_io_x_ppn),
    .io_x_u(OptimizationBarrier_23_io_x_u),
    .io_x_ae(OptimizationBarrier_23_io_x_ae),
    .io_x_sw(OptimizationBarrier_23_io_x_sw),
    .io_x_sx(OptimizationBarrier_23_io_x_sx),
    .io_x_sr(OptimizationBarrier_23_io_x_sr),
    .io_x_pw(OptimizationBarrier_23_io_x_pw),
    .io_x_px(OptimizationBarrier_23_io_x_px),
    .io_x_pr(OptimizationBarrier_23_io_x_pr),
    .io_x_ppp(OptimizationBarrier_23_io_x_ppp),
    .io_x_pal(OptimizationBarrier_23_io_x_pal),
    .io_x_paa(OptimizationBarrier_23_io_x_paa),
    .io_x_eff(OptimizationBarrier_23_io_x_eff),
    .io_x_c(OptimizationBarrier_23_io_x_c),
    .io_y_ppn(OptimizationBarrier_23_io_y_ppn),
    .io_y_u(OptimizationBarrier_23_io_y_u),
    .io_y_ae(OptimizationBarrier_23_io_y_ae),
    .io_y_sw(OptimizationBarrier_23_io_y_sw),
    .io_y_sx(OptimizationBarrier_23_io_y_sx),
    .io_y_sr(OptimizationBarrier_23_io_y_sr),
    .io_y_pw(OptimizationBarrier_23_io_y_pw),
    .io_y_px(OptimizationBarrier_23_io_y_px),
    .io_y_pr(OptimizationBarrier_23_io_y_pr),
    .io_y_ppp(OptimizationBarrier_23_io_y_ppp),
    .io_y_pal(OptimizationBarrier_23_io_y_pal),
    .io_y_paa(OptimizationBarrier_23_io_y_paa),
    .io_y_eff(OptimizationBarrier_23_io_y_eff),
    .io_y_c(OptimizationBarrier_23_io_y_c)
  );
  OptimizationBarrier OptimizationBarrier_24 ( // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@200586.4]
    .io_x_ppn(OptimizationBarrier_24_io_x_ppn),
    .io_x_u(OptimizationBarrier_24_io_x_u),
    .io_x_ae(OptimizationBarrier_24_io_x_ae),
    .io_x_sw(OptimizationBarrier_24_io_x_sw),
    .io_x_sx(OptimizationBarrier_24_io_x_sx),
    .io_x_sr(OptimizationBarrier_24_io_x_sr),
    .io_x_pw(OptimizationBarrier_24_io_x_pw),
    .io_x_px(OptimizationBarrier_24_io_x_px),
    .io_x_pr(OptimizationBarrier_24_io_x_pr),
    .io_x_ppp(OptimizationBarrier_24_io_x_ppp),
    .io_x_pal(OptimizationBarrier_24_io_x_pal),
    .io_x_paa(OptimizationBarrier_24_io_x_paa),
    .io_x_eff(OptimizationBarrier_24_io_x_eff),
    .io_x_c(OptimizationBarrier_24_io_x_c),
    .io_y_ppn(OptimizationBarrier_24_io_y_ppn),
    .io_y_u(OptimizationBarrier_24_io_y_u),
    .io_y_ae(OptimizationBarrier_24_io_y_ae),
    .io_y_sw(OptimizationBarrier_24_io_y_sw),
    .io_y_sx(OptimizationBarrier_24_io_y_sx),
    .io_y_sr(OptimizationBarrier_24_io_y_sr),
    .io_y_pw(OptimizationBarrier_24_io_y_pw),
    .io_y_px(OptimizationBarrier_24_io_y_px),
    .io_y_pr(OptimizationBarrier_24_io_y_pr),
    .io_y_ppp(OptimizationBarrier_24_io_y_ppp),
    .io_y_pal(OptimizationBarrier_24_io_y_pal),
    .io_y_paa(OptimizationBarrier_24_io_y_paa),
    .io_y_eff(OptimizationBarrier_24_io_y_eff),
    .io_y_c(OptimizationBarrier_24_io_y_c)
  );
  OptimizationBarrier OptimizationBarrier_25 ( // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@200628.4]
    .io_x_ppn(OptimizationBarrier_25_io_x_ppn),
    .io_x_u(OptimizationBarrier_25_io_x_u),
    .io_x_ae(OptimizationBarrier_25_io_x_ae),
    .io_x_sw(OptimizationBarrier_25_io_x_sw),
    .io_x_sx(OptimizationBarrier_25_io_x_sx),
    .io_x_sr(OptimizationBarrier_25_io_x_sr),
    .io_x_pw(OptimizationBarrier_25_io_x_pw),
    .io_x_px(OptimizationBarrier_25_io_x_px),
    .io_x_pr(OptimizationBarrier_25_io_x_pr),
    .io_x_ppp(OptimizationBarrier_25_io_x_ppp),
    .io_x_pal(OptimizationBarrier_25_io_x_pal),
    .io_x_paa(OptimizationBarrier_25_io_x_paa),
    .io_x_eff(OptimizationBarrier_25_io_x_eff),
    .io_x_c(OptimizationBarrier_25_io_x_c),
    .io_y_ppn(OptimizationBarrier_25_io_y_ppn),
    .io_y_u(OptimizationBarrier_25_io_y_u),
    .io_y_ae(OptimizationBarrier_25_io_y_ae),
    .io_y_sw(OptimizationBarrier_25_io_y_sw),
    .io_y_sx(OptimizationBarrier_25_io_y_sx),
    .io_y_sr(OptimizationBarrier_25_io_y_sr),
    .io_y_pw(OptimizationBarrier_25_io_y_pw),
    .io_y_px(OptimizationBarrier_25_io_y_px),
    .io_y_pr(OptimizationBarrier_25_io_y_pr),
    .io_y_ppp(OptimizationBarrier_25_io_y_ppp),
    .io_y_pal(OptimizationBarrier_25_io_y_pal),
    .io_y_paa(OptimizationBarrier_25_io_y_paa),
    .io_y_eff(OptimizationBarrier_25_io_y_eff),
    .io_y_c(OptimizationBarrier_25_io_y_c)
  );
  OptimizationBarrier OptimizationBarrier_26 ( // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@200670.4]
    .io_x_ppn(OptimizationBarrier_26_io_x_ppn),
    .io_x_u(OptimizationBarrier_26_io_x_u),
    .io_x_ae(OptimizationBarrier_26_io_x_ae),
    .io_x_sw(OptimizationBarrier_26_io_x_sw),
    .io_x_sx(OptimizationBarrier_26_io_x_sx),
    .io_x_sr(OptimizationBarrier_26_io_x_sr),
    .io_x_pw(OptimizationBarrier_26_io_x_pw),
    .io_x_px(OptimizationBarrier_26_io_x_px),
    .io_x_pr(OptimizationBarrier_26_io_x_pr),
    .io_x_ppp(OptimizationBarrier_26_io_x_ppp),
    .io_x_pal(OptimizationBarrier_26_io_x_pal),
    .io_x_paa(OptimizationBarrier_26_io_x_paa),
    .io_x_eff(OptimizationBarrier_26_io_x_eff),
    .io_x_c(OptimizationBarrier_26_io_x_c),
    .io_y_ppn(OptimizationBarrier_26_io_y_ppn),
    .io_y_u(OptimizationBarrier_26_io_y_u),
    .io_y_ae(OptimizationBarrier_26_io_y_ae),
    .io_y_sw(OptimizationBarrier_26_io_y_sw),
    .io_y_sx(OptimizationBarrier_26_io_y_sx),
    .io_y_sr(OptimizationBarrier_26_io_y_sr),
    .io_y_pw(OptimizationBarrier_26_io_y_pw),
    .io_y_px(OptimizationBarrier_26_io_y_px),
    .io_y_pr(OptimizationBarrier_26_io_y_pr),
    .io_y_ppp(OptimizationBarrier_26_io_y_ppp),
    .io_y_pal(OptimizationBarrier_26_io_y_pal),
    .io_y_paa(OptimizationBarrier_26_io_y_paa),
    .io_y_eff(OptimizationBarrier_26_io_y_eff),
    .io_y_c(OptimizationBarrier_26_io_y_c)
  );
  OptimizationBarrier OptimizationBarrier_27 ( // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@200713.4]
    .io_x_ppn(OptimizationBarrier_27_io_x_ppn),
    .io_x_u(OptimizationBarrier_27_io_x_u),
    .io_x_ae(OptimizationBarrier_27_io_x_ae),
    .io_x_sw(OptimizationBarrier_27_io_x_sw),
    .io_x_sx(OptimizationBarrier_27_io_x_sx),
    .io_x_sr(OptimizationBarrier_27_io_x_sr),
    .io_x_pw(OptimizationBarrier_27_io_x_pw),
    .io_x_px(OptimizationBarrier_27_io_x_px),
    .io_x_pr(OptimizationBarrier_27_io_x_pr),
    .io_x_ppp(OptimizationBarrier_27_io_x_ppp),
    .io_x_pal(OptimizationBarrier_27_io_x_pal),
    .io_x_paa(OptimizationBarrier_27_io_x_paa),
    .io_x_eff(OptimizationBarrier_27_io_x_eff),
    .io_x_c(OptimizationBarrier_27_io_x_c),
    .io_y_ppn(OptimizationBarrier_27_io_y_ppn),
    .io_y_u(OptimizationBarrier_27_io_y_u),
    .io_y_ae(OptimizationBarrier_27_io_y_ae),
    .io_y_sw(OptimizationBarrier_27_io_y_sw),
    .io_y_sx(OptimizationBarrier_27_io_y_sx),
    .io_y_sr(OptimizationBarrier_27_io_y_sr),
    .io_y_pw(OptimizationBarrier_27_io_y_pw),
    .io_y_px(OptimizationBarrier_27_io_y_px),
    .io_y_pr(OptimizationBarrier_27_io_y_pr),
    .io_y_ppp(OptimizationBarrier_27_io_y_ppp),
    .io_y_pal(OptimizationBarrier_27_io_y_pal),
    .io_y_paa(OptimizationBarrier_27_io_y_paa),
    .io_y_eff(OptimizationBarrier_27_io_y_eff),
    .io_y_c(OptimizationBarrier_27_io_y_c)
  );
  OptimizationBarrier OptimizationBarrier_28 ( // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@200756.4]
    .io_x_ppn(OptimizationBarrier_28_io_x_ppn),
    .io_x_u(OptimizationBarrier_28_io_x_u),
    .io_x_ae(OptimizationBarrier_28_io_x_ae),
    .io_x_sw(OptimizationBarrier_28_io_x_sw),
    .io_x_sx(OptimizationBarrier_28_io_x_sx),
    .io_x_sr(OptimizationBarrier_28_io_x_sr),
    .io_x_pw(OptimizationBarrier_28_io_x_pw),
    .io_x_px(OptimizationBarrier_28_io_x_px),
    .io_x_pr(OptimizationBarrier_28_io_x_pr),
    .io_x_ppp(OptimizationBarrier_28_io_x_ppp),
    .io_x_pal(OptimizationBarrier_28_io_x_pal),
    .io_x_paa(OptimizationBarrier_28_io_x_paa),
    .io_x_eff(OptimizationBarrier_28_io_x_eff),
    .io_x_c(OptimizationBarrier_28_io_x_c),
    .io_y_ppn(OptimizationBarrier_28_io_y_ppn),
    .io_y_u(OptimizationBarrier_28_io_y_u),
    .io_y_ae(OptimizationBarrier_28_io_y_ae),
    .io_y_sw(OptimizationBarrier_28_io_y_sw),
    .io_y_sx(OptimizationBarrier_28_io_y_sx),
    .io_y_sr(OptimizationBarrier_28_io_y_sr),
    .io_y_pw(OptimizationBarrier_28_io_y_pw),
    .io_y_px(OptimizationBarrier_28_io_y_px),
    .io_y_pr(OptimizationBarrier_28_io_y_pr),
    .io_y_ppp(OptimizationBarrier_28_io_y_ppp),
    .io_y_pal(OptimizationBarrier_28_io_y_pal),
    .io_y_paa(OptimizationBarrier_28_io_y_paa),
    .io_y_eff(OptimizationBarrier_28_io_y_eff),
    .io_y_c(OptimizationBarrier_28_io_y_c)
  );
  OptimizationBarrier OptimizationBarrier_29 ( // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@200799.4]
    .io_x_ppn(OptimizationBarrier_29_io_x_ppn),
    .io_x_u(OptimizationBarrier_29_io_x_u),
    .io_x_ae(OptimizationBarrier_29_io_x_ae),
    .io_x_sw(OptimizationBarrier_29_io_x_sw),
    .io_x_sx(OptimizationBarrier_29_io_x_sx),
    .io_x_sr(OptimizationBarrier_29_io_x_sr),
    .io_x_pw(OptimizationBarrier_29_io_x_pw),
    .io_x_px(OptimizationBarrier_29_io_x_px),
    .io_x_pr(OptimizationBarrier_29_io_x_pr),
    .io_x_ppp(OptimizationBarrier_29_io_x_ppp),
    .io_x_pal(OptimizationBarrier_29_io_x_pal),
    .io_x_paa(OptimizationBarrier_29_io_x_paa),
    .io_x_eff(OptimizationBarrier_29_io_x_eff),
    .io_x_c(OptimizationBarrier_29_io_x_c),
    .io_y_ppn(OptimizationBarrier_29_io_y_ppn),
    .io_y_u(OptimizationBarrier_29_io_y_u),
    .io_y_ae(OptimizationBarrier_29_io_y_ae),
    .io_y_sw(OptimizationBarrier_29_io_y_sw),
    .io_y_sx(OptimizationBarrier_29_io_y_sx),
    .io_y_sr(OptimizationBarrier_29_io_y_sr),
    .io_y_pw(OptimizationBarrier_29_io_y_pw),
    .io_y_px(OptimizationBarrier_29_io_y_px),
    .io_y_pr(OptimizationBarrier_29_io_y_pr),
    .io_y_ppp(OptimizationBarrier_29_io_y_ppp),
    .io_y_pal(OptimizationBarrier_29_io_y_pal),
    .io_y_paa(OptimizationBarrier_29_io_y_paa),
    .io_y_eff(OptimizationBarrier_29_io_y_eff),
    .io_y_c(OptimizationBarrier_29_io_y_c)
  );
  OptimizationBarrier OptimizationBarrier_30 ( // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@200842.4]
    .io_x_ppn(OptimizationBarrier_30_io_x_ppn),
    .io_x_u(OptimizationBarrier_30_io_x_u),
    .io_x_ae(OptimizationBarrier_30_io_x_ae),
    .io_x_sw(OptimizationBarrier_30_io_x_sw),
    .io_x_sx(OptimizationBarrier_30_io_x_sx),
    .io_x_sr(OptimizationBarrier_30_io_x_sr),
    .io_x_pw(OptimizationBarrier_30_io_x_pw),
    .io_x_px(OptimizationBarrier_30_io_x_px),
    .io_x_pr(OptimizationBarrier_30_io_x_pr),
    .io_x_ppp(OptimizationBarrier_30_io_x_ppp),
    .io_x_pal(OptimizationBarrier_30_io_x_pal),
    .io_x_paa(OptimizationBarrier_30_io_x_paa),
    .io_x_eff(OptimizationBarrier_30_io_x_eff),
    .io_x_c(OptimizationBarrier_30_io_x_c),
    .io_y_ppn(OptimizationBarrier_30_io_y_ppn),
    .io_y_u(OptimizationBarrier_30_io_y_u),
    .io_y_ae(OptimizationBarrier_30_io_y_ae),
    .io_y_sw(OptimizationBarrier_30_io_y_sw),
    .io_y_sx(OptimizationBarrier_30_io_y_sx),
    .io_y_sr(OptimizationBarrier_30_io_y_sr),
    .io_y_pw(OptimizationBarrier_30_io_y_pw),
    .io_y_px(OptimizationBarrier_30_io_y_px),
    .io_y_pr(OptimizationBarrier_30_io_y_pr),
    .io_y_ppp(OptimizationBarrier_30_io_y_ppp),
    .io_y_pal(OptimizationBarrier_30_io_y_pal),
    .io_y_paa(OptimizationBarrier_30_io_y_paa),
    .io_y_eff(OptimizationBarrier_30_io_y_eff),
    .io_y_c(OptimizationBarrier_30_io_y_c)
  );
  OptimizationBarrier OptimizationBarrier_31 ( // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@200885.4]
    .io_x_ppn(OptimizationBarrier_31_io_x_ppn),
    .io_x_u(OptimizationBarrier_31_io_x_u),
    .io_x_ae(OptimizationBarrier_31_io_x_ae),
    .io_x_sw(OptimizationBarrier_31_io_x_sw),
    .io_x_sx(OptimizationBarrier_31_io_x_sx),
    .io_x_sr(OptimizationBarrier_31_io_x_sr),
    .io_x_pw(OptimizationBarrier_31_io_x_pw),
    .io_x_px(OptimizationBarrier_31_io_x_px),
    .io_x_pr(OptimizationBarrier_31_io_x_pr),
    .io_x_ppp(OptimizationBarrier_31_io_x_ppp),
    .io_x_pal(OptimizationBarrier_31_io_x_pal),
    .io_x_paa(OptimizationBarrier_31_io_x_paa),
    .io_x_eff(OptimizationBarrier_31_io_x_eff),
    .io_x_c(OptimizationBarrier_31_io_x_c),
    .io_y_ppn(OptimizationBarrier_31_io_y_ppn),
    .io_y_u(OptimizationBarrier_31_io_y_u),
    .io_y_ae(OptimizationBarrier_31_io_y_ae),
    .io_y_sw(OptimizationBarrier_31_io_y_sw),
    .io_y_sx(OptimizationBarrier_31_io_y_sx),
    .io_y_sr(OptimizationBarrier_31_io_y_sr),
    .io_y_pw(OptimizationBarrier_31_io_y_pw),
    .io_y_px(OptimizationBarrier_31_io_y_px),
    .io_y_pr(OptimizationBarrier_31_io_y_pr),
    .io_y_ppp(OptimizationBarrier_31_io_y_ppp),
    .io_y_pal(OptimizationBarrier_31_io_y_pal),
    .io_y_paa(OptimizationBarrier_31_io_y_paa),
    .io_y_eff(OptimizationBarrier_31_io_y_eff),
    .io_y_c(OptimizationBarrier_31_io_y_c)
  );
  OptimizationBarrier OptimizationBarrier_32 ( // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@200928.4]
    .io_x_ppn(OptimizationBarrier_32_io_x_ppn),
    .io_x_u(OptimizationBarrier_32_io_x_u),
    .io_x_ae(OptimizationBarrier_32_io_x_ae),
    .io_x_sw(OptimizationBarrier_32_io_x_sw),
    .io_x_sx(OptimizationBarrier_32_io_x_sx),
    .io_x_sr(OptimizationBarrier_32_io_x_sr),
    .io_x_pw(OptimizationBarrier_32_io_x_pw),
    .io_x_px(OptimizationBarrier_32_io_x_px),
    .io_x_pr(OptimizationBarrier_32_io_x_pr),
    .io_x_ppp(OptimizationBarrier_32_io_x_ppp),
    .io_x_pal(OptimizationBarrier_32_io_x_pal),
    .io_x_paa(OptimizationBarrier_32_io_x_paa),
    .io_x_eff(OptimizationBarrier_32_io_x_eff),
    .io_x_c(OptimizationBarrier_32_io_x_c),
    .io_y_ppn(OptimizationBarrier_32_io_y_ppn),
    .io_y_u(OptimizationBarrier_32_io_y_u),
    .io_y_ae(OptimizationBarrier_32_io_y_ae),
    .io_y_sw(OptimizationBarrier_32_io_y_sw),
    .io_y_sx(OptimizationBarrier_32_io_y_sx),
    .io_y_sr(OptimizationBarrier_32_io_y_sr),
    .io_y_pw(OptimizationBarrier_32_io_y_pw),
    .io_y_px(OptimizationBarrier_32_io_y_px),
    .io_y_pr(OptimizationBarrier_32_io_y_pr),
    .io_y_ppp(OptimizationBarrier_32_io_y_ppp),
    .io_y_pal(OptimizationBarrier_32_io_y_pal),
    .io_y_paa(OptimizationBarrier_32_io_y_paa),
    .io_y_eff(OptimizationBarrier_32_io_y_eff),
    .io_y_c(OptimizationBarrier_32_io_y_c)
  );
  OptimizationBarrier OptimizationBarrier_33 ( // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@200971.4]
    .io_x_ppn(OptimizationBarrier_33_io_x_ppn),
    .io_x_u(OptimizationBarrier_33_io_x_u),
    .io_x_ae(OptimizationBarrier_33_io_x_ae),
    .io_x_sw(OptimizationBarrier_33_io_x_sw),
    .io_x_sx(OptimizationBarrier_33_io_x_sx),
    .io_x_sr(OptimizationBarrier_33_io_x_sr),
    .io_x_pw(OptimizationBarrier_33_io_x_pw),
    .io_x_px(OptimizationBarrier_33_io_x_px),
    .io_x_pr(OptimizationBarrier_33_io_x_pr),
    .io_x_ppp(OptimizationBarrier_33_io_x_ppp),
    .io_x_pal(OptimizationBarrier_33_io_x_pal),
    .io_x_paa(OptimizationBarrier_33_io_x_paa),
    .io_x_eff(OptimizationBarrier_33_io_x_eff),
    .io_x_c(OptimizationBarrier_33_io_x_c),
    .io_y_ppn(OptimizationBarrier_33_io_y_ppn),
    .io_y_u(OptimizationBarrier_33_io_y_u),
    .io_y_ae(OptimizationBarrier_33_io_y_ae),
    .io_y_sw(OptimizationBarrier_33_io_y_sw),
    .io_y_sx(OptimizationBarrier_33_io_y_sx),
    .io_y_sr(OptimizationBarrier_33_io_y_sr),
    .io_y_pw(OptimizationBarrier_33_io_y_pw),
    .io_y_px(OptimizationBarrier_33_io_y_px),
    .io_y_pr(OptimizationBarrier_33_io_y_pr),
    .io_y_ppp(OptimizationBarrier_33_io_y_ppp),
    .io_y_pal(OptimizationBarrier_33_io_y_pal),
    .io_y_paa(OptimizationBarrier_33_io_y_paa),
    .io_y_eff(OptimizationBarrier_33_io_y_eff),
    .io_y_c(OptimizationBarrier_33_io_y_c)
  );
  OptimizationBarrier OptimizationBarrier_34 ( // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@201014.4]
    .io_x_ppn(OptimizationBarrier_34_io_x_ppn),
    .io_x_u(OptimizationBarrier_34_io_x_u),
    .io_x_ae(OptimizationBarrier_34_io_x_ae),
    .io_x_sw(OptimizationBarrier_34_io_x_sw),
    .io_x_sx(OptimizationBarrier_34_io_x_sx),
    .io_x_sr(OptimizationBarrier_34_io_x_sr),
    .io_x_pw(OptimizationBarrier_34_io_x_pw),
    .io_x_px(OptimizationBarrier_34_io_x_px),
    .io_x_pr(OptimizationBarrier_34_io_x_pr),
    .io_x_ppp(OptimizationBarrier_34_io_x_ppp),
    .io_x_pal(OptimizationBarrier_34_io_x_pal),
    .io_x_paa(OptimizationBarrier_34_io_x_paa),
    .io_x_eff(OptimizationBarrier_34_io_x_eff),
    .io_x_c(OptimizationBarrier_34_io_x_c),
    .io_y_ppn(OptimizationBarrier_34_io_y_ppn),
    .io_y_u(OptimizationBarrier_34_io_y_u),
    .io_y_ae(OptimizationBarrier_34_io_y_ae),
    .io_y_sw(OptimizationBarrier_34_io_y_sw),
    .io_y_sx(OptimizationBarrier_34_io_y_sx),
    .io_y_sr(OptimizationBarrier_34_io_y_sr),
    .io_y_pw(OptimizationBarrier_34_io_y_pw),
    .io_y_px(OptimizationBarrier_34_io_y_px),
    .io_y_pr(OptimizationBarrier_34_io_y_pr),
    .io_y_ppp(OptimizationBarrier_34_io_y_ppp),
    .io_y_pal(OptimizationBarrier_34_io_y_pal),
    .io_y_paa(OptimizationBarrier_34_io_y_paa),
    .io_y_eff(OptimizationBarrier_34_io_y_eff),
    .io_y_c(OptimizationBarrier_34_io_y_c)
  );
  OptimizationBarrier OptimizationBarrier_35 ( // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@201056.4]
    .io_x_ppn(OptimizationBarrier_35_io_x_ppn),
    .io_x_u(OptimizationBarrier_35_io_x_u),
    .io_x_ae(OptimizationBarrier_35_io_x_ae),
    .io_x_sw(OptimizationBarrier_35_io_x_sw),
    .io_x_sx(OptimizationBarrier_35_io_x_sx),
    .io_x_sr(OptimizationBarrier_35_io_x_sr),
    .io_x_pw(OptimizationBarrier_35_io_x_pw),
    .io_x_px(OptimizationBarrier_35_io_x_px),
    .io_x_pr(OptimizationBarrier_35_io_x_pr),
    .io_x_ppp(OptimizationBarrier_35_io_x_ppp),
    .io_x_pal(OptimizationBarrier_35_io_x_pal),
    .io_x_paa(OptimizationBarrier_35_io_x_paa),
    .io_x_eff(OptimizationBarrier_35_io_x_eff),
    .io_x_c(OptimizationBarrier_35_io_x_c),
    .io_y_ppn(OptimizationBarrier_35_io_y_ppn),
    .io_y_u(OptimizationBarrier_35_io_y_u),
    .io_y_ae(OptimizationBarrier_35_io_y_ae),
    .io_y_sw(OptimizationBarrier_35_io_y_sw),
    .io_y_sx(OptimizationBarrier_35_io_y_sx),
    .io_y_sr(OptimizationBarrier_35_io_y_sr),
    .io_y_pw(OptimizationBarrier_35_io_y_pw),
    .io_y_px(OptimizationBarrier_35_io_y_px),
    .io_y_pr(OptimizationBarrier_35_io_y_pr),
    .io_y_ppp(OptimizationBarrier_35_io_y_ppp),
    .io_y_pal(OptimizationBarrier_35_io_y_pal),
    .io_y_paa(OptimizationBarrier_35_io_y_paa),
    .io_y_eff(OptimizationBarrier_35_io_y_eff),
    .io_y_c(OptimizationBarrier_35_io_y_c)
  );
  OptimizationBarrier OptimizationBarrier_36 ( // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@201098.4]
    .io_x_ppn(OptimizationBarrier_36_io_x_ppn),
    .io_x_u(OptimizationBarrier_36_io_x_u),
    .io_x_ae(OptimizationBarrier_36_io_x_ae),
    .io_x_sw(OptimizationBarrier_36_io_x_sw),
    .io_x_sx(OptimizationBarrier_36_io_x_sx),
    .io_x_sr(OptimizationBarrier_36_io_x_sr),
    .io_x_pw(OptimizationBarrier_36_io_x_pw),
    .io_x_px(OptimizationBarrier_36_io_x_px),
    .io_x_pr(OptimizationBarrier_36_io_x_pr),
    .io_x_ppp(OptimizationBarrier_36_io_x_ppp),
    .io_x_pal(OptimizationBarrier_36_io_x_pal),
    .io_x_paa(OptimizationBarrier_36_io_x_paa),
    .io_x_eff(OptimizationBarrier_36_io_x_eff),
    .io_x_c(OptimizationBarrier_36_io_x_c),
    .io_y_ppn(OptimizationBarrier_36_io_y_ppn),
    .io_y_u(OptimizationBarrier_36_io_y_u),
    .io_y_ae(OptimizationBarrier_36_io_y_ae),
    .io_y_sw(OptimizationBarrier_36_io_y_sw),
    .io_y_sx(OptimizationBarrier_36_io_y_sx),
    .io_y_sr(OptimizationBarrier_36_io_y_sr),
    .io_y_pw(OptimizationBarrier_36_io_y_pw),
    .io_y_px(OptimizationBarrier_36_io_y_px),
    .io_y_pr(OptimizationBarrier_36_io_y_pr),
    .io_y_ppp(OptimizationBarrier_36_io_y_ppp),
    .io_y_pal(OptimizationBarrier_36_io_y_pal),
    .io_y_paa(OptimizationBarrier_36_io_y_paa),
    .io_y_eff(OptimizationBarrier_36_io_y_eff),
    .io_y_c(OptimizationBarrier_36_io_y_c)
  );
  OptimizationBarrier OptimizationBarrier_37 ( // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@201140.4]
    .io_x_ppn(OptimizationBarrier_37_io_x_ppn),
    .io_x_u(OptimizationBarrier_37_io_x_u),
    .io_x_ae(OptimizationBarrier_37_io_x_ae),
    .io_x_sw(OptimizationBarrier_37_io_x_sw),
    .io_x_sx(OptimizationBarrier_37_io_x_sx),
    .io_x_sr(OptimizationBarrier_37_io_x_sr),
    .io_x_pw(OptimizationBarrier_37_io_x_pw),
    .io_x_px(OptimizationBarrier_37_io_x_px),
    .io_x_pr(OptimizationBarrier_37_io_x_pr),
    .io_x_ppp(OptimizationBarrier_37_io_x_ppp),
    .io_x_pal(OptimizationBarrier_37_io_x_pal),
    .io_x_paa(OptimizationBarrier_37_io_x_paa),
    .io_x_eff(OptimizationBarrier_37_io_x_eff),
    .io_x_c(OptimizationBarrier_37_io_x_c),
    .io_y_ppn(OptimizationBarrier_37_io_y_ppn),
    .io_y_u(OptimizationBarrier_37_io_y_u),
    .io_y_ae(OptimizationBarrier_37_io_y_ae),
    .io_y_sw(OptimizationBarrier_37_io_y_sw),
    .io_y_sx(OptimizationBarrier_37_io_y_sx),
    .io_y_sr(OptimizationBarrier_37_io_y_sr),
    .io_y_pw(OptimizationBarrier_37_io_y_pw),
    .io_y_px(OptimizationBarrier_37_io_y_px),
    .io_y_pr(OptimizationBarrier_37_io_y_pr),
    .io_y_ppp(OptimizationBarrier_37_io_y_ppp),
    .io_y_pal(OptimizationBarrier_37_io_y_pal),
    .io_y_paa(OptimizationBarrier_37_io_y_paa),
    .io_y_eff(OptimizationBarrier_37_io_y_eff),
    .io_y_c(OptimizationBarrier_37_io_y_c)
  );
  OptimizationBarrier OptimizationBarrier_38 ( // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@201182.4]
    .io_x_ppn(OptimizationBarrier_38_io_x_ppn),
    .io_x_u(OptimizationBarrier_38_io_x_u),
    .io_x_ae(OptimizationBarrier_38_io_x_ae),
    .io_x_sw(OptimizationBarrier_38_io_x_sw),
    .io_x_sx(OptimizationBarrier_38_io_x_sx),
    .io_x_sr(OptimizationBarrier_38_io_x_sr),
    .io_x_pw(OptimizationBarrier_38_io_x_pw),
    .io_x_px(OptimizationBarrier_38_io_x_px),
    .io_x_pr(OptimizationBarrier_38_io_x_pr),
    .io_x_ppp(OptimizationBarrier_38_io_x_ppp),
    .io_x_pal(OptimizationBarrier_38_io_x_pal),
    .io_x_paa(OptimizationBarrier_38_io_x_paa),
    .io_x_eff(OptimizationBarrier_38_io_x_eff),
    .io_x_c(OptimizationBarrier_38_io_x_c),
    .io_y_ppn(OptimizationBarrier_38_io_y_ppn),
    .io_y_u(OptimizationBarrier_38_io_y_u),
    .io_y_ae(OptimizationBarrier_38_io_y_ae),
    .io_y_sw(OptimizationBarrier_38_io_y_sw),
    .io_y_sx(OptimizationBarrier_38_io_y_sx),
    .io_y_sr(OptimizationBarrier_38_io_y_sr),
    .io_y_pw(OptimizationBarrier_38_io_y_pw),
    .io_y_px(OptimizationBarrier_38_io_y_px),
    .io_y_pr(OptimizationBarrier_38_io_y_pr),
    .io_y_ppp(OptimizationBarrier_38_io_y_ppp),
    .io_y_pal(OptimizationBarrier_38_io_y_pal),
    .io_y_paa(OptimizationBarrier_38_io_y_paa),
    .io_y_eff(OptimizationBarrier_38_io_y_eff),
    .io_y_c(OptimizationBarrier_38_io_y_c)
  );
  assign priv_s = io_ptw_status_prv[0]; // @[TLB.scala 177:20:freechips.rocketchip.system.DefaultRV32Config.fir@198366.4]
  assign priv_uses_vm = io_ptw_status_prv <= 2'h1; // @[TLB.scala 178:27:freechips.rocketchip.system.DefaultRV32Config.fir@198367.4]
  assign vm_enabled = io_ptw_ptbr_mode & priv_uses_vm; // @[TLB.scala 179:83:freechips.rocketchip.system.DefaultRV32Config.fir@198370.4]
  assign vpn = io_req_bits_vaddr[31:12]; // @[TLB.scala 182:30:freechips.rocketchip.system.DefaultRV32Config.fir@198373.4]
  assign refill_ppn = io_ptw_resp_bits_pte_ppn[19:0]; // @[TLB.scala 183:44:freechips.rocketchip.system.DefaultRV32Config.fir@198374.4]
  assign _T_4 = state == 2'h1; // @[package.scala 15:47:freechips.rocketchip.system.DefaultRV32Config.fir@198376.4]
  assign _T_5 = state == 2'h3; // @[package.scala 15:47:freechips.rocketchip.system.DefaultRV32Config.fir@198377.4]
  assign invalidate_refill = _T_4 | _T_5; // @[package.scala 64:59:freechips.rocketchip.system.DefaultRV32Config.fir@198378.4]
  assign _T_26 = special_entry_level < 1'h1; // @[TLB.scala 108:28:freechips.rocketchip.system.DefaultRV32Config.fir@198423.4]
  assign _T_28 = _T_26 ? vpn : 20'h0; // @[TLB.scala 109:28:freechips.rocketchip.system.DefaultRV32Config.fir@198425.4]
  assign _T_29 = _T_28 | OptimizationBarrier_io_y_ppn; // @[TLB.scala 109:47:freechips.rocketchip.system.DefaultRV32Config.fir@198426.4]
  assign _T_31 = {OptimizationBarrier_io_y_ppn[19:10],_T_29[9:0]}; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@198428.4]
  assign _T_33 = vm_enabled ? _T_31 : io_req_bits_vaddr[31:12]; // @[TLB.scala 187:20:freechips.rocketchip.system.DefaultRV32Config.fir@198430.4]
  assign mpu_ppn = io_ptw_resp_valid ? refill_ppn : _T_33; // @[TLB.scala 186:20:freechips.rocketchip.system.DefaultRV32Config.fir@198431.4]
  assign mpu_physaddr = {mpu_ppn,io_req_bits_vaddr[11:0]}; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@198433.4]
  assign _T_37 = {io_ptw_status_debug,io_ptw_status_prv}; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@198436.4]
  assign mpu_priv = io_ptw_resp_valid ? 3'h1 : _T_37; // @[TLB.scala 189:27:freechips.rocketchip.system.DefaultRV32Config.fir@198437.4]
  assign _T_38 = mpu_physaddr ^ 32'h3000; // @[Parameters.scala 137:31:freechips.rocketchip.system.DefaultRV32Config.fir@198453.4]
  assign _T_39 = {1'b0,$signed(_T_38)}; // @[Parameters.scala 137:49:freechips.rocketchip.system.DefaultRV32Config.fir@198454.4]
  assign _T_41 = $signed(_T_39) & -33'sh1000; // @[Parameters.scala 137:52:freechips.rocketchip.system.DefaultRV32Config.fir@198456.4]
  assign _T_42 = $signed(_T_41) == 33'sh0; // @[Parameters.scala 137:67:freechips.rocketchip.system.DefaultRV32Config.fir@198457.4]
  assign _T_43 = mpu_physaddr ^ 32'hc000000; // @[Parameters.scala 137:31:freechips.rocketchip.system.DefaultRV32Config.fir@198458.4]
  assign _T_44 = {1'b0,$signed(_T_43)}; // @[Parameters.scala 137:49:freechips.rocketchip.system.DefaultRV32Config.fir@198459.4]
  assign _T_46 = $signed(_T_44) & -33'sh4000000; // @[Parameters.scala 137:52:freechips.rocketchip.system.DefaultRV32Config.fir@198461.4]
  assign _T_47 = $signed(_T_46) == 33'sh0; // @[Parameters.scala 137:67:freechips.rocketchip.system.DefaultRV32Config.fir@198462.4]
  assign _T_48 = mpu_physaddr ^ 32'h2000000; // @[Parameters.scala 137:31:freechips.rocketchip.system.DefaultRV32Config.fir@198463.4]
  assign _T_49 = {1'b0,$signed(_T_48)}; // @[Parameters.scala 137:49:freechips.rocketchip.system.DefaultRV32Config.fir@198464.4]
  assign _T_51 = $signed(_T_49) & -33'sh10000; // @[Parameters.scala 137:52:freechips.rocketchip.system.DefaultRV32Config.fir@198466.4]
  assign _T_52 = $signed(_T_51) == 33'sh0; // @[Parameters.scala 137:67:freechips.rocketchip.system.DefaultRV32Config.fir@198467.4]
  assign _T_54 = {1'b0,$signed(mpu_physaddr)}; // @[Parameters.scala 137:49:freechips.rocketchip.system.DefaultRV32Config.fir@198469.4]
  assign _T_56 = $signed(_T_54) & -33'sh1000; // @[Parameters.scala 137:52:freechips.rocketchip.system.DefaultRV32Config.fir@198471.4]
  assign _T_57 = $signed(_T_56) == 33'sh0; // @[Parameters.scala 137:67:freechips.rocketchip.system.DefaultRV32Config.fir@198472.4]
  assign _T_58 = mpu_physaddr ^ 32'h10000; // @[Parameters.scala 137:31:freechips.rocketchip.system.DefaultRV32Config.fir@198473.4]
  assign _T_59 = {1'b0,$signed(_T_58)}; // @[Parameters.scala 137:49:freechips.rocketchip.system.DefaultRV32Config.fir@198474.4]
  assign _T_61 = $signed(_T_59) & -33'sh10000; // @[Parameters.scala 137:52:freechips.rocketchip.system.DefaultRV32Config.fir@198476.4]
  assign _T_62 = $signed(_T_61) == 33'sh0; // @[Parameters.scala 137:67:freechips.rocketchip.system.DefaultRV32Config.fir@198477.4]
  assign _T_63 = mpu_physaddr ^ 32'h80000000; // @[Parameters.scala 137:31:freechips.rocketchip.system.DefaultRV32Config.fir@198478.4]
  assign _T_64 = {1'b0,$signed(_T_63)}; // @[Parameters.scala 137:49:freechips.rocketchip.system.DefaultRV32Config.fir@198479.4]
  assign _T_66 = $signed(_T_64) & -33'sh10000000; // @[Parameters.scala 137:52:freechips.rocketchip.system.DefaultRV32Config.fir@198481.4]
  assign _T_67 = $signed(_T_66) == 33'sh0; // @[Parameters.scala 137:67:freechips.rocketchip.system.DefaultRV32Config.fir@198482.4]
  assign _T_68 = mpu_physaddr ^ 32'h60000000; // @[Parameters.scala 137:31:freechips.rocketchip.system.DefaultRV32Config.fir@198483.4]
  assign _T_69 = {1'b0,$signed(_T_68)}; // @[Parameters.scala 137:49:freechips.rocketchip.system.DefaultRV32Config.fir@198484.4]
  assign _T_71 = $signed(_T_69) & -33'sh20000000; // @[Parameters.scala 137:52:freechips.rocketchip.system.DefaultRV32Config.fir@198486.4]
  assign _T_72 = $signed(_T_71) == 33'sh0; // @[Parameters.scala 137:67:freechips.rocketchip.system.DefaultRV32Config.fir@198487.4]
  assign _T_74 = _T_42 | _T_47; // @[TLB.scala 195:67:freechips.rocketchip.system.DefaultRV32Config.fir@198497.4]
  assign _T_75 = _T_74 | _T_52; // @[TLB.scala 195:67:freechips.rocketchip.system.DefaultRV32Config.fir@198498.4]
  assign _T_76 = _T_75 | _T_57; // @[TLB.scala 195:67:freechips.rocketchip.system.DefaultRV32Config.fir@198499.4]
  assign _T_77 = _T_76 | _T_62; // @[TLB.scala 195:67:freechips.rocketchip.system.DefaultRV32Config.fir@198500.4]
  assign _T_78 = _T_77 | _T_67; // @[TLB.scala 195:67:freechips.rocketchip.system.DefaultRV32Config.fir@198501.4]
  assign legal_address = _T_78 | _T_72; // @[TLB.scala 195:67:freechips.rocketchip.system.DefaultRV32Config.fir@198502.4]
  assign _T_87 = $signed(_T_64) & 33'sh80000000; // @[Parameters.scala 137:52:freechips.rocketchip.system.DefaultRV32Config.fir@198511.4]
  assign _T_88 = $signed(_T_87) == 33'sh0; // @[Parameters.scala 137:67:freechips.rocketchip.system.DefaultRV32Config.fir@198512.4]
  assign cacheable = legal_address & _T_88; // @[TLB.scala 197:19:freechips.rocketchip.system.DefaultRV32Config.fir@198518.4]
  assign _T_148 = mpu_physaddr ^ 32'h8000000; // @[Parameters.scala 137:31:freechips.rocketchip.system.DefaultRV32Config.fir@198575.4]
  assign _T_149 = {1'b0,$signed(_T_148)}; // @[Parameters.scala 137:49:freechips.rocketchip.system.DefaultRV32Config.fir@198576.4]
  assign _T_151 = $signed(_T_149) & 33'shc8000000; // @[Parameters.scala 137:52:freechips.rocketchip.system.DefaultRV32Config.fir@198578.4]
  assign _T_152 = $signed(_T_151) == 33'sh0; // @[Parameters.scala 137:67:freechips.rocketchip.system.DefaultRV32Config.fir@198579.4]
  assign _T_165 = $signed(_T_54) & 33'shc8010000; // @[Parameters.scala 137:52:freechips.rocketchip.system.DefaultRV32Config.fir@198592.4]
  assign _T_166 = $signed(_T_165) == 33'sh0; // @[Parameters.scala 137:67:freechips.rocketchip.system.DefaultRV32Config.fir@198593.4]
  assign _T_173 = _T_166 | _T_152; // @[TLBPermissions.scala 82:66:freechips.rocketchip.system.DefaultRV32Config.fir@198600.4]
  assign _T_186 = mpu_priv <= 3'h3; // @[TLB.scala 200:39:freechips.rocketchip.system.DefaultRV32Config.fir@198613.4]
  assign deny_access_to_debug = _T_186 & _T_57; // @[TLB.scala 200:48:freechips.rocketchip.system.DefaultRV32Config.fir@198619.4]
  assign _T_198 = ~deny_access_to_debug; // @[TLB.scala 201:44:freechips.rocketchip.system.DefaultRV32Config.fir@198626.4]
  assign _T_199 = legal_address & _T_198; // @[TLB.scala 201:41:freechips.rocketchip.system.DefaultRV32Config.fir@198627.4]
  assign prot_r = _T_199 & pmp_io_r; // @[TLB.scala 201:66:freechips.rocketchip.system.DefaultRV32Config.fir@198628.4]
  assign _T_210 = mpu_physaddr ^ 32'h40000000; // @[Parameters.scala 137:31:freechips.rocketchip.system.DefaultRV32Config.fir@198639.4]
  assign _T_211 = {1'b0,$signed(_T_210)}; // @[Parameters.scala 137:49:freechips.rocketchip.system.DefaultRV32Config.fir@198640.4]
  assign _T_213 = $signed(_T_211) & 33'shc0000000; // @[Parameters.scala 137:52:freechips.rocketchip.system.DefaultRV32Config.fir@198642.4]
  assign _T_214 = $signed(_T_213) == 33'sh0; // @[Parameters.scala 137:67:freechips.rocketchip.system.DefaultRV32Config.fir@198643.4]
  assign _T_218 = $signed(_T_64) & 33'shc0000000; // @[Parameters.scala 137:52:freechips.rocketchip.system.DefaultRV32Config.fir@198647.4]
  assign _T_219 = $signed(_T_218) == 33'sh0; // @[Parameters.scala 137:67:freechips.rocketchip.system.DefaultRV32Config.fir@198648.4]
  assign _T_221 = _T_173 | _T_214; // @[Parameters.scala 528:89:freechips.rocketchip.system.DefaultRV32Config.fir@198650.4]
  assign _T_222 = _T_221 | _T_219; // @[Parameters.scala 528:89:freechips.rocketchip.system.DefaultRV32Config.fir@198651.4]
  assign _T_232 = legal_address & _T_222; // @[TLB.scala 197:19:freechips.rocketchip.system.DefaultRV32Config.fir@198662.4]
  assign _T_234 = _T_232 & _T_198; // @[TLB.scala 202:45:freechips.rocketchip.system.DefaultRV32Config.fir@198664.4]
  assign prot_w = _T_234 & pmp_io_w; // @[TLB.scala 202:70:freechips.rocketchip.system.DefaultRV32Config.fir@198665.4]
  assign prot_al = legal_address & _T_173; // @[TLB.scala 197:19:freechips.rocketchip.system.DefaultRV32Config.fir@198733.4]
  assign _T_334 = $signed(_T_54) & 33'shca000000; // @[Parameters.scala 137:52:freechips.rocketchip.system.DefaultRV32Config.fir@198771.4]
  assign _T_335 = $signed(_T_334) == 33'sh0; // @[Parameters.scala 137:67:freechips.rocketchip.system.DefaultRV32Config.fir@198772.4]
  assign _T_346 = _T_335 | _T_214; // @[Parameters.scala 528:89:freechips.rocketchip.system.DefaultRV32Config.fir@198783.4]
  assign _T_347 = _T_346 | _T_219; // @[Parameters.scala 528:89:freechips.rocketchip.system.DefaultRV32Config.fir@198784.4]
  assign _T_363 = legal_address & _T_347; // @[TLB.scala 197:19:freechips.rocketchip.system.DefaultRV32Config.fir@198801.4]
  assign _T_365 = _T_363 & _T_198; // @[TLB.scala 206:40:freechips.rocketchip.system.DefaultRV32Config.fir@198803.4]
  assign prot_x = _T_365 & pmp_io_x; // @[TLB.scala 206:65:freechips.rocketchip.system.DefaultRV32Config.fir@198804.4]
  assign _T_386 = $signed(_T_54) & 33'shca012000; // @[Parameters.scala 137:52:freechips.rocketchip.system.DefaultRV32Config.fir@198825.4]
  assign _T_387 = $signed(_T_386) == 33'sh0; // @[Parameters.scala 137:67:freechips.rocketchip.system.DefaultRV32Config.fir@198826.4]
  assign _T_391 = $signed(_T_49) & 33'shca010000; // @[Parameters.scala 137:52:freechips.rocketchip.system.DefaultRV32Config.fir@198830.4]
  assign _T_392 = $signed(_T_391) == 33'sh0; // @[Parameters.scala 137:67:freechips.rocketchip.system.DefaultRV32Config.fir@198831.4]
  assign _T_403 = _T_387 | _T_392; // @[Parameters.scala 528:89:freechips.rocketchip.system.DefaultRV32Config.fir@198842.4]
  assign _T_404 = _T_403 | _T_152; // @[Parameters.scala 528:89:freechips.rocketchip.system.DefaultRV32Config.fir@198843.4]
  assign _T_405 = _T_404 | _T_214; // @[Parameters.scala 528:89:freechips.rocketchip.system.DefaultRV32Config.fir@198844.4]
  assign prot_eff = legal_address & _T_405; // @[TLB.scala 197:19:freechips.rocketchip.system.DefaultRV32Config.fir@198850.4]
  assign _T_410 = sectored_entries_0_valid_0 | sectored_entries_0_valid_1; // @[package.scala 64:59:freechips.rocketchip.system.DefaultRV32Config.fir@198851.4]
  assign _T_411 = _T_410 | sectored_entries_0_valid_2; // @[package.scala 64:59:freechips.rocketchip.system.DefaultRV32Config.fir@198852.4]
  assign _T_412 = _T_411 | sectored_entries_0_valid_3; // @[package.scala 64:59:freechips.rocketchip.system.DefaultRV32Config.fir@198853.4]
  assign _T_413 = sectored_entries_0_tag ^ vpn; // @[TLB.scala 88:41:freechips.rocketchip.system.DefaultRV32Config.fir@198854.4]
  assign _T_415 = _T_413[19:2] == 18'h0; // @[TLB.scala 88:66:freechips.rocketchip.system.DefaultRV32Config.fir@198856.4]
  assign sector_hits_0 = _T_412 & _T_415; // @[TLB.scala 87:40:freechips.rocketchip.system.DefaultRV32Config.fir@198857.4]
  assign _T_416 = sectored_entries_1_valid_0 | sectored_entries_1_valid_1; // @[package.scala 64:59:freechips.rocketchip.system.DefaultRV32Config.fir@198858.4]
  assign _T_417 = _T_416 | sectored_entries_1_valid_2; // @[package.scala 64:59:freechips.rocketchip.system.DefaultRV32Config.fir@198859.4]
  assign _T_418 = _T_417 | sectored_entries_1_valid_3; // @[package.scala 64:59:freechips.rocketchip.system.DefaultRV32Config.fir@198860.4]
  assign _T_419 = sectored_entries_1_tag ^ vpn; // @[TLB.scala 88:41:freechips.rocketchip.system.DefaultRV32Config.fir@198861.4]
  assign _T_421 = _T_419[19:2] == 18'h0; // @[TLB.scala 88:66:freechips.rocketchip.system.DefaultRV32Config.fir@198863.4]
  assign sector_hits_1 = _T_418 & _T_421; // @[TLB.scala 87:40:freechips.rocketchip.system.DefaultRV32Config.fir@198864.4]
  assign _T_422 = sectored_entries_2_valid_0 | sectored_entries_2_valid_1; // @[package.scala 64:59:freechips.rocketchip.system.DefaultRV32Config.fir@198865.4]
  assign _T_423 = _T_422 | sectored_entries_2_valid_2; // @[package.scala 64:59:freechips.rocketchip.system.DefaultRV32Config.fir@198866.4]
  assign _T_424 = _T_423 | sectored_entries_2_valid_3; // @[package.scala 64:59:freechips.rocketchip.system.DefaultRV32Config.fir@198867.4]
  assign _T_425 = sectored_entries_2_tag ^ vpn; // @[TLB.scala 88:41:freechips.rocketchip.system.DefaultRV32Config.fir@198868.4]
  assign _T_427 = _T_425[19:2] == 18'h0; // @[TLB.scala 88:66:freechips.rocketchip.system.DefaultRV32Config.fir@198870.4]
  assign sector_hits_2 = _T_424 & _T_427; // @[TLB.scala 87:40:freechips.rocketchip.system.DefaultRV32Config.fir@198871.4]
  assign _T_428 = sectored_entries_3_valid_0 | sectored_entries_3_valid_1; // @[package.scala 64:59:freechips.rocketchip.system.DefaultRV32Config.fir@198872.4]
  assign _T_429 = _T_428 | sectored_entries_3_valid_2; // @[package.scala 64:59:freechips.rocketchip.system.DefaultRV32Config.fir@198873.4]
  assign _T_430 = _T_429 | sectored_entries_3_valid_3; // @[package.scala 64:59:freechips.rocketchip.system.DefaultRV32Config.fir@198874.4]
  assign _T_431 = sectored_entries_3_tag ^ vpn; // @[TLB.scala 88:41:freechips.rocketchip.system.DefaultRV32Config.fir@198875.4]
  assign _T_433 = _T_431[19:2] == 18'h0; // @[TLB.scala 88:66:freechips.rocketchip.system.DefaultRV32Config.fir@198877.4]
  assign sector_hits_3 = _T_430 & _T_433; // @[TLB.scala 87:40:freechips.rocketchip.system.DefaultRV32Config.fir@198878.4]
  assign _T_434 = sectored_entries_4_valid_0 | sectored_entries_4_valid_1; // @[package.scala 64:59:freechips.rocketchip.system.DefaultRV32Config.fir@198879.4]
  assign _T_435 = _T_434 | sectored_entries_4_valid_2; // @[package.scala 64:59:freechips.rocketchip.system.DefaultRV32Config.fir@198880.4]
  assign _T_436 = _T_435 | sectored_entries_4_valid_3; // @[package.scala 64:59:freechips.rocketchip.system.DefaultRV32Config.fir@198881.4]
  assign _T_437 = sectored_entries_4_tag ^ vpn; // @[TLB.scala 88:41:freechips.rocketchip.system.DefaultRV32Config.fir@198882.4]
  assign _T_439 = _T_437[19:2] == 18'h0; // @[TLB.scala 88:66:freechips.rocketchip.system.DefaultRV32Config.fir@198884.4]
  assign sector_hits_4 = _T_436 & _T_439; // @[TLB.scala 87:40:freechips.rocketchip.system.DefaultRV32Config.fir@198885.4]
  assign _T_440 = sectored_entries_5_valid_0 | sectored_entries_5_valid_1; // @[package.scala 64:59:freechips.rocketchip.system.DefaultRV32Config.fir@198886.4]
  assign _T_441 = _T_440 | sectored_entries_5_valid_2; // @[package.scala 64:59:freechips.rocketchip.system.DefaultRV32Config.fir@198887.4]
  assign _T_442 = _T_441 | sectored_entries_5_valid_3; // @[package.scala 64:59:freechips.rocketchip.system.DefaultRV32Config.fir@198888.4]
  assign _T_443 = sectored_entries_5_tag ^ vpn; // @[TLB.scala 88:41:freechips.rocketchip.system.DefaultRV32Config.fir@198889.4]
  assign _T_445 = _T_443[19:2] == 18'h0; // @[TLB.scala 88:66:freechips.rocketchip.system.DefaultRV32Config.fir@198891.4]
  assign sector_hits_5 = _T_442 & _T_445; // @[TLB.scala 87:40:freechips.rocketchip.system.DefaultRV32Config.fir@198892.4]
  assign _T_446 = sectored_entries_6_valid_0 | sectored_entries_6_valid_1; // @[package.scala 64:59:freechips.rocketchip.system.DefaultRV32Config.fir@198893.4]
  assign _T_447 = _T_446 | sectored_entries_6_valid_2; // @[package.scala 64:59:freechips.rocketchip.system.DefaultRV32Config.fir@198894.4]
  assign _T_448 = _T_447 | sectored_entries_6_valid_3; // @[package.scala 64:59:freechips.rocketchip.system.DefaultRV32Config.fir@198895.4]
  assign _T_449 = sectored_entries_6_tag ^ vpn; // @[TLB.scala 88:41:freechips.rocketchip.system.DefaultRV32Config.fir@198896.4]
  assign _T_451 = _T_449[19:2] == 18'h0; // @[TLB.scala 88:66:freechips.rocketchip.system.DefaultRV32Config.fir@198898.4]
  assign sector_hits_6 = _T_448 & _T_451; // @[TLB.scala 87:40:freechips.rocketchip.system.DefaultRV32Config.fir@198899.4]
  assign _T_452 = sectored_entries_7_valid_0 | sectored_entries_7_valid_1; // @[package.scala 64:59:freechips.rocketchip.system.DefaultRV32Config.fir@198900.4]
  assign _T_453 = _T_452 | sectored_entries_7_valid_2; // @[package.scala 64:59:freechips.rocketchip.system.DefaultRV32Config.fir@198901.4]
  assign _T_454 = _T_453 | sectored_entries_7_valid_3; // @[package.scala 64:59:freechips.rocketchip.system.DefaultRV32Config.fir@198902.4]
  assign _T_455 = sectored_entries_7_tag ^ vpn; // @[TLB.scala 88:41:freechips.rocketchip.system.DefaultRV32Config.fir@198903.4]
  assign _T_457 = _T_455[19:2] == 18'h0; // @[TLB.scala 88:66:freechips.rocketchip.system.DefaultRV32Config.fir@198905.4]
  assign sector_hits_7 = _T_454 & _T_457; // @[TLB.scala 87:40:freechips.rocketchip.system.DefaultRV32Config.fir@198906.4]
  assign _T_462 = superpage_entries_0_tag[19:10] == vpn[19:10]; // @[TLB.scala 95:77:freechips.rocketchip.system.DefaultRV32Config.fir@198911.4]
  assign superpage_hits_0 = superpage_entries_0_valid_0 & _T_462; // @[TLB.scala 95:29:freechips.rocketchip.system.DefaultRV32Config.fir@198913.4]
  assign _T_475 = superpage_entries_1_tag[19:10] == vpn[19:10]; // @[TLB.scala 95:77:freechips.rocketchip.system.DefaultRV32Config.fir@198925.4]
  assign superpage_hits_1 = superpage_entries_1_valid_0 & _T_475; // @[TLB.scala 95:29:freechips.rocketchip.system.DefaultRV32Config.fir@198927.4]
  assign _T_488 = superpage_entries_2_tag[19:10] == vpn[19:10]; // @[TLB.scala 95:77:freechips.rocketchip.system.DefaultRV32Config.fir@198939.4]
  assign superpage_hits_2 = superpage_entries_2_valid_0 & _T_488; // @[TLB.scala 95:29:freechips.rocketchip.system.DefaultRV32Config.fir@198941.4]
  assign _T_501 = superpage_entries_3_tag[19:10] == vpn[19:10]; // @[TLB.scala 95:77:freechips.rocketchip.system.DefaultRV32Config.fir@198953.4]
  assign superpage_hits_3 = superpage_entries_3_valid_0 & _T_501; // @[TLB.scala 95:29:freechips.rocketchip.system.DefaultRV32Config.fir@198955.4]
  assign _GEN_1 = 2'h1 == vpn[1:0] ? sectored_entries_0_valid_1 : sectored_entries_0_valid_0; // @[TLB.scala 100:18:freechips.rocketchip.system.DefaultRV32Config.fir@198967.4]
  assign _GEN_2 = 2'h2 == vpn[1:0] ? sectored_entries_0_valid_2 : _GEN_1; // @[TLB.scala 100:18:freechips.rocketchip.system.DefaultRV32Config.fir@198967.4]
  assign _GEN_3 = 2'h3 == vpn[1:0] ? sectored_entries_0_valid_3 : _GEN_2; // @[TLB.scala 100:18:freechips.rocketchip.system.DefaultRV32Config.fir@198967.4]
  assign _T_514 = _GEN_3 & _T_415; // @[TLB.scala 100:18:freechips.rocketchip.system.DefaultRV32Config.fir@198967.4]
  assign hitsVec_0 = vm_enabled & _T_514; // @[TLB.scala 211:44:freechips.rocketchip.system.DefaultRV32Config.fir@198968.4]
  assign _GEN_5 = 2'h1 == vpn[1:0] ? sectored_entries_1_valid_1 : sectored_entries_1_valid_0; // @[TLB.scala 100:18:freechips.rocketchip.system.DefaultRV32Config.fir@198973.4]
  assign _GEN_6 = 2'h2 == vpn[1:0] ? sectored_entries_1_valid_2 : _GEN_5; // @[TLB.scala 100:18:freechips.rocketchip.system.DefaultRV32Config.fir@198973.4]
  assign _GEN_7 = 2'h3 == vpn[1:0] ? sectored_entries_1_valid_3 : _GEN_6; // @[TLB.scala 100:18:freechips.rocketchip.system.DefaultRV32Config.fir@198973.4]
  assign _T_519 = _GEN_7 & _T_421; // @[TLB.scala 100:18:freechips.rocketchip.system.DefaultRV32Config.fir@198973.4]
  assign hitsVec_1 = vm_enabled & _T_519; // @[TLB.scala 211:44:freechips.rocketchip.system.DefaultRV32Config.fir@198974.4]
  assign _GEN_9 = 2'h1 == vpn[1:0] ? sectored_entries_2_valid_1 : sectored_entries_2_valid_0; // @[TLB.scala 100:18:freechips.rocketchip.system.DefaultRV32Config.fir@198979.4]
  assign _GEN_10 = 2'h2 == vpn[1:0] ? sectored_entries_2_valid_2 : _GEN_9; // @[TLB.scala 100:18:freechips.rocketchip.system.DefaultRV32Config.fir@198979.4]
  assign _GEN_11 = 2'h3 == vpn[1:0] ? sectored_entries_2_valid_3 : _GEN_10; // @[TLB.scala 100:18:freechips.rocketchip.system.DefaultRV32Config.fir@198979.4]
  assign _T_524 = _GEN_11 & _T_427; // @[TLB.scala 100:18:freechips.rocketchip.system.DefaultRV32Config.fir@198979.4]
  assign hitsVec_2 = vm_enabled & _T_524; // @[TLB.scala 211:44:freechips.rocketchip.system.DefaultRV32Config.fir@198980.4]
  assign _GEN_13 = 2'h1 == vpn[1:0] ? sectored_entries_3_valid_1 : sectored_entries_3_valid_0; // @[TLB.scala 100:18:freechips.rocketchip.system.DefaultRV32Config.fir@198985.4]
  assign _GEN_14 = 2'h2 == vpn[1:0] ? sectored_entries_3_valid_2 : _GEN_13; // @[TLB.scala 100:18:freechips.rocketchip.system.DefaultRV32Config.fir@198985.4]
  assign _GEN_15 = 2'h3 == vpn[1:0] ? sectored_entries_3_valid_3 : _GEN_14; // @[TLB.scala 100:18:freechips.rocketchip.system.DefaultRV32Config.fir@198985.4]
  assign _T_529 = _GEN_15 & _T_433; // @[TLB.scala 100:18:freechips.rocketchip.system.DefaultRV32Config.fir@198985.4]
  assign hitsVec_3 = vm_enabled & _T_529; // @[TLB.scala 211:44:freechips.rocketchip.system.DefaultRV32Config.fir@198986.4]
  assign _GEN_17 = 2'h1 == vpn[1:0] ? sectored_entries_4_valid_1 : sectored_entries_4_valid_0; // @[TLB.scala 100:18:freechips.rocketchip.system.DefaultRV32Config.fir@198991.4]
  assign _GEN_18 = 2'h2 == vpn[1:0] ? sectored_entries_4_valid_2 : _GEN_17; // @[TLB.scala 100:18:freechips.rocketchip.system.DefaultRV32Config.fir@198991.4]
  assign _GEN_19 = 2'h3 == vpn[1:0] ? sectored_entries_4_valid_3 : _GEN_18; // @[TLB.scala 100:18:freechips.rocketchip.system.DefaultRV32Config.fir@198991.4]
  assign _T_534 = _GEN_19 & _T_439; // @[TLB.scala 100:18:freechips.rocketchip.system.DefaultRV32Config.fir@198991.4]
  assign hitsVec_4 = vm_enabled & _T_534; // @[TLB.scala 211:44:freechips.rocketchip.system.DefaultRV32Config.fir@198992.4]
  assign _GEN_21 = 2'h1 == vpn[1:0] ? sectored_entries_5_valid_1 : sectored_entries_5_valid_0; // @[TLB.scala 100:18:freechips.rocketchip.system.DefaultRV32Config.fir@198997.4]
  assign _GEN_22 = 2'h2 == vpn[1:0] ? sectored_entries_5_valid_2 : _GEN_21; // @[TLB.scala 100:18:freechips.rocketchip.system.DefaultRV32Config.fir@198997.4]
  assign _GEN_23 = 2'h3 == vpn[1:0] ? sectored_entries_5_valid_3 : _GEN_22; // @[TLB.scala 100:18:freechips.rocketchip.system.DefaultRV32Config.fir@198997.4]
  assign _T_539 = _GEN_23 & _T_445; // @[TLB.scala 100:18:freechips.rocketchip.system.DefaultRV32Config.fir@198997.4]
  assign hitsVec_5 = vm_enabled & _T_539; // @[TLB.scala 211:44:freechips.rocketchip.system.DefaultRV32Config.fir@198998.4]
  assign _GEN_25 = 2'h1 == vpn[1:0] ? sectored_entries_6_valid_1 : sectored_entries_6_valid_0; // @[TLB.scala 100:18:freechips.rocketchip.system.DefaultRV32Config.fir@199003.4]
  assign _GEN_26 = 2'h2 == vpn[1:0] ? sectored_entries_6_valid_2 : _GEN_25; // @[TLB.scala 100:18:freechips.rocketchip.system.DefaultRV32Config.fir@199003.4]
  assign _GEN_27 = 2'h3 == vpn[1:0] ? sectored_entries_6_valid_3 : _GEN_26; // @[TLB.scala 100:18:freechips.rocketchip.system.DefaultRV32Config.fir@199003.4]
  assign _T_544 = _GEN_27 & _T_451; // @[TLB.scala 100:18:freechips.rocketchip.system.DefaultRV32Config.fir@199003.4]
  assign hitsVec_6 = vm_enabled & _T_544; // @[TLB.scala 211:44:freechips.rocketchip.system.DefaultRV32Config.fir@199004.4]
  assign _GEN_29 = 2'h1 == vpn[1:0] ? sectored_entries_7_valid_1 : sectored_entries_7_valid_0; // @[TLB.scala 100:18:freechips.rocketchip.system.DefaultRV32Config.fir@199009.4]
  assign _GEN_30 = 2'h2 == vpn[1:0] ? sectored_entries_7_valid_2 : _GEN_29; // @[TLB.scala 100:18:freechips.rocketchip.system.DefaultRV32Config.fir@199009.4]
  assign _GEN_31 = 2'h3 == vpn[1:0] ? sectored_entries_7_valid_3 : _GEN_30; // @[TLB.scala 100:18:freechips.rocketchip.system.DefaultRV32Config.fir@199009.4]
  assign _T_549 = _GEN_31 & _T_457; // @[TLB.scala 100:18:freechips.rocketchip.system.DefaultRV32Config.fir@199009.4]
  assign hitsVec_7 = vm_enabled & _T_549; // @[TLB.scala 211:44:freechips.rocketchip.system.DefaultRV32Config.fir@199010.4]
  assign hitsVec_8 = vm_enabled & superpage_hits_0; // @[TLB.scala 211:44:freechips.rocketchip.system.DefaultRV32Config.fir@199025.4]
  assign hitsVec_9 = vm_enabled & superpage_hits_1; // @[TLB.scala 211:44:freechips.rocketchip.system.DefaultRV32Config.fir@199040.4]
  assign hitsVec_10 = vm_enabled & superpage_hits_2; // @[TLB.scala 211:44:freechips.rocketchip.system.DefaultRV32Config.fir@199055.4]
  assign hitsVec_11 = vm_enabled & superpage_hits_3; // @[TLB.scala 211:44:freechips.rocketchip.system.DefaultRV32Config.fir@199070.4]
  assign _T_610 = special_entry_tag[19:10] == vpn[19:10]; // @[TLB.scala 95:77:freechips.rocketchip.system.DefaultRV32Config.fir@199075.4]
  assign _T_612 = special_entry_valid_0 & _T_610; // @[TLB.scala 95:29:freechips.rocketchip.system.DefaultRV32Config.fir@199077.4]
  assign _T_617 = special_entry_tag[9:0] == vpn[9:0]; // @[TLB.scala 95:77:freechips.rocketchip.system.DefaultRV32Config.fir@199082.4]
  assign _T_618 = _T_26 | _T_617; // @[TLB.scala 95:40:freechips.rocketchip.system.DefaultRV32Config.fir@199083.4]
  assign _T_619 = _T_612 & _T_618; // @[TLB.scala 95:29:freechips.rocketchip.system.DefaultRV32Config.fir@199084.4]
  assign hitsVec_12 = vm_enabled & _T_619; // @[TLB.scala 211:44:freechips.rocketchip.system.DefaultRV32Config.fir@199085.4]
  assign _T_624 = {hitsVec_5,hitsVec_4,hitsVec_3,hitsVec_2,hitsVec_1,hitsVec_0}; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@199090.4]
  assign real_hits = {hitsVec_12,hitsVec_11,hitsVec_10,hitsVec_9,hitsVec_8,hitsVec_7,hitsVec_6,_T_624}; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@199097.4]
  assign _T_631 = ~vm_enabled; // @[TLB.scala 213:18:freechips.rocketchip.system.DefaultRV32Config.fir@199098.4]
  assign hits = {_T_631,hitsVec_12,hitsVec_11,hitsVec_10,hitsVec_9,hitsVec_8,hitsVec_7,hitsVec_6,_T_624}; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@199099.4]
  assign _GEN_33 = 2'h1 == vpn[1:0] ? sectored_entries_0_data_1 : sectored_entries_0_data_0; // @[:freechips.rocketchip.system.DefaultRV32Config.fir@199106.4]
  assign _GEN_34 = 2'h2 == vpn[1:0] ? sectored_entries_0_data_2 : _GEN_33; // @[:freechips.rocketchip.system.DefaultRV32Config.fir@199106.4]
  assign _GEN_35 = 2'h3 == vpn[1:0] ? sectored_entries_0_data_3 : _GEN_34; // @[:freechips.rocketchip.system.DefaultRV32Config.fir@199106.4]
  assign _GEN_37 = 2'h1 == vpn[1:0] ? sectored_entries_1_data_1 : sectored_entries_1_data_0; // @[:freechips.rocketchip.system.DefaultRV32Config.fir@199149.4]
  assign _GEN_38 = 2'h2 == vpn[1:0] ? sectored_entries_1_data_2 : _GEN_37; // @[:freechips.rocketchip.system.DefaultRV32Config.fir@199149.4]
  assign _GEN_39 = 2'h3 == vpn[1:0] ? sectored_entries_1_data_3 : _GEN_38; // @[:freechips.rocketchip.system.DefaultRV32Config.fir@199149.4]
  assign _GEN_41 = 2'h1 == vpn[1:0] ? sectored_entries_2_data_1 : sectored_entries_2_data_0; // @[:freechips.rocketchip.system.DefaultRV32Config.fir@199192.4]
  assign _GEN_42 = 2'h2 == vpn[1:0] ? sectored_entries_2_data_2 : _GEN_41; // @[:freechips.rocketchip.system.DefaultRV32Config.fir@199192.4]
  assign _GEN_43 = 2'h3 == vpn[1:0] ? sectored_entries_2_data_3 : _GEN_42; // @[:freechips.rocketchip.system.DefaultRV32Config.fir@199192.4]
  assign _GEN_45 = 2'h1 == vpn[1:0] ? sectored_entries_3_data_1 : sectored_entries_3_data_0; // @[:freechips.rocketchip.system.DefaultRV32Config.fir@199235.4]
  assign _GEN_46 = 2'h2 == vpn[1:0] ? sectored_entries_3_data_2 : _GEN_45; // @[:freechips.rocketchip.system.DefaultRV32Config.fir@199235.4]
  assign _GEN_47 = 2'h3 == vpn[1:0] ? sectored_entries_3_data_3 : _GEN_46; // @[:freechips.rocketchip.system.DefaultRV32Config.fir@199235.4]
  assign _GEN_49 = 2'h1 == vpn[1:0] ? sectored_entries_4_data_1 : sectored_entries_4_data_0; // @[:freechips.rocketchip.system.DefaultRV32Config.fir@199278.4]
  assign _GEN_50 = 2'h2 == vpn[1:0] ? sectored_entries_4_data_2 : _GEN_49; // @[:freechips.rocketchip.system.DefaultRV32Config.fir@199278.4]
  assign _GEN_51 = 2'h3 == vpn[1:0] ? sectored_entries_4_data_3 : _GEN_50; // @[:freechips.rocketchip.system.DefaultRV32Config.fir@199278.4]
  assign _GEN_53 = 2'h1 == vpn[1:0] ? sectored_entries_5_data_1 : sectored_entries_5_data_0; // @[:freechips.rocketchip.system.DefaultRV32Config.fir@199321.4]
  assign _GEN_54 = 2'h2 == vpn[1:0] ? sectored_entries_5_data_2 : _GEN_53; // @[:freechips.rocketchip.system.DefaultRV32Config.fir@199321.4]
  assign _GEN_55 = 2'h3 == vpn[1:0] ? sectored_entries_5_data_3 : _GEN_54; // @[:freechips.rocketchip.system.DefaultRV32Config.fir@199321.4]
  assign _GEN_57 = 2'h1 == vpn[1:0] ? sectored_entries_6_data_1 : sectored_entries_6_data_0; // @[:freechips.rocketchip.system.DefaultRV32Config.fir@199364.4]
  assign _GEN_58 = 2'h2 == vpn[1:0] ? sectored_entries_6_data_2 : _GEN_57; // @[:freechips.rocketchip.system.DefaultRV32Config.fir@199364.4]
  assign _GEN_59 = 2'h3 == vpn[1:0] ? sectored_entries_6_data_3 : _GEN_58; // @[:freechips.rocketchip.system.DefaultRV32Config.fir@199364.4]
  assign _GEN_61 = 2'h1 == vpn[1:0] ? sectored_entries_7_data_1 : sectored_entries_7_data_0; // @[:freechips.rocketchip.system.DefaultRV32Config.fir@199407.4]
  assign _GEN_62 = 2'h2 == vpn[1:0] ? sectored_entries_7_data_2 : _GEN_61; // @[:freechips.rocketchip.system.DefaultRV32Config.fir@199407.4]
  assign _GEN_63 = 2'h3 == vpn[1:0] ? sectored_entries_7_data_3 : _GEN_62; // @[:freechips.rocketchip.system.DefaultRV32Config.fir@199407.4]
  assign _T_807 = vpn | OptimizationBarrier_9_io_y_ppn; // @[TLB.scala 109:47:freechips.rocketchip.system.DefaultRV32Config.fir@199491.4]
  assign _T_809 = {OptimizationBarrier_9_io_y_ppn[19:10],_T_807[9:0]}; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@199493.4]
  assign _T_832 = vpn | OptimizationBarrier_10_io_y_ppn; // @[TLB.scala 109:47:freechips.rocketchip.system.DefaultRV32Config.fir@199540.4]
  assign _T_834 = {OptimizationBarrier_10_io_y_ppn[19:10],_T_832[9:0]}; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@199542.4]
  assign _T_857 = vpn | OptimizationBarrier_11_io_y_ppn; // @[TLB.scala 109:47:freechips.rocketchip.system.DefaultRV32Config.fir@199589.4]
  assign _T_859 = {OptimizationBarrier_11_io_y_ppn[19:10],_T_857[9:0]}; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@199591.4]
  assign _T_882 = vpn | OptimizationBarrier_12_io_y_ppn; // @[TLB.scala 109:47:freechips.rocketchip.system.DefaultRV32Config.fir@199638.4]
  assign _T_884 = {OptimizationBarrier_12_io_y_ppn[19:10],_T_882[9:0]}; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@199640.4]
  assign _T_907 = _T_28 | OptimizationBarrier_13_io_y_ppn; // @[TLB.scala 109:47:freechips.rocketchip.system.DefaultRV32Config.fir@199687.4]
  assign _T_909 = {OptimizationBarrier_13_io_y_ppn[19:10],_T_907[9:0]}; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@199689.4]
  assign _T_911 = hitsVec_0 ? OptimizationBarrier_1_io_y_ppn : 20'h0; // @[Mux.scala 27:72:freechips.rocketchip.system.DefaultRV32Config.fir@199691.4]
  assign _T_912 = hitsVec_1 ? OptimizationBarrier_2_io_y_ppn : 20'h0; // @[Mux.scala 27:72:freechips.rocketchip.system.DefaultRV32Config.fir@199692.4]
  assign _T_913 = hitsVec_2 ? OptimizationBarrier_3_io_y_ppn : 20'h0; // @[Mux.scala 27:72:freechips.rocketchip.system.DefaultRV32Config.fir@199693.4]
  assign _T_914 = hitsVec_3 ? OptimizationBarrier_4_io_y_ppn : 20'h0; // @[Mux.scala 27:72:freechips.rocketchip.system.DefaultRV32Config.fir@199694.4]
  assign _T_915 = hitsVec_4 ? OptimizationBarrier_5_io_y_ppn : 20'h0; // @[Mux.scala 27:72:freechips.rocketchip.system.DefaultRV32Config.fir@199695.4]
  assign _T_916 = hitsVec_5 ? OptimizationBarrier_6_io_y_ppn : 20'h0; // @[Mux.scala 27:72:freechips.rocketchip.system.DefaultRV32Config.fir@199696.4]
  assign _T_917 = hitsVec_6 ? OptimizationBarrier_7_io_y_ppn : 20'h0; // @[Mux.scala 27:72:freechips.rocketchip.system.DefaultRV32Config.fir@199697.4]
  assign _T_918 = hitsVec_7 ? OptimizationBarrier_8_io_y_ppn : 20'h0; // @[Mux.scala 27:72:freechips.rocketchip.system.DefaultRV32Config.fir@199698.4]
  assign _T_919 = hitsVec_8 ? _T_809 : 20'h0; // @[Mux.scala 27:72:freechips.rocketchip.system.DefaultRV32Config.fir@199699.4]
  assign _T_920 = hitsVec_9 ? _T_834 : 20'h0; // @[Mux.scala 27:72:freechips.rocketchip.system.DefaultRV32Config.fir@199700.4]
  assign _T_921 = hitsVec_10 ? _T_859 : 20'h0; // @[Mux.scala 27:72:freechips.rocketchip.system.DefaultRV32Config.fir@199701.4]
  assign _T_922 = hitsVec_11 ? _T_884 : 20'h0; // @[Mux.scala 27:72:freechips.rocketchip.system.DefaultRV32Config.fir@199702.4]
  assign _T_923 = hitsVec_12 ? _T_909 : 20'h0; // @[Mux.scala 27:72:freechips.rocketchip.system.DefaultRV32Config.fir@199703.4]
  assign _T_924 = _T_631 ? vpn : 20'h0; // @[Mux.scala 27:72:freechips.rocketchip.system.DefaultRV32Config.fir@199704.4]
  assign _T_925 = _T_911 | _T_912; // @[Mux.scala 27:72:freechips.rocketchip.system.DefaultRV32Config.fir@199705.4]
  assign _T_926 = _T_925 | _T_913; // @[Mux.scala 27:72:freechips.rocketchip.system.DefaultRV32Config.fir@199706.4]
  assign _T_927 = _T_926 | _T_914; // @[Mux.scala 27:72:freechips.rocketchip.system.DefaultRV32Config.fir@199707.4]
  assign _T_928 = _T_927 | _T_915; // @[Mux.scala 27:72:freechips.rocketchip.system.DefaultRV32Config.fir@199708.4]
  assign _T_929 = _T_928 | _T_916; // @[Mux.scala 27:72:freechips.rocketchip.system.DefaultRV32Config.fir@199709.4]
  assign _T_930 = _T_929 | _T_917; // @[Mux.scala 27:72:freechips.rocketchip.system.DefaultRV32Config.fir@199710.4]
  assign _T_931 = _T_930 | _T_918; // @[Mux.scala 27:72:freechips.rocketchip.system.DefaultRV32Config.fir@199711.4]
  assign _T_932 = _T_931 | _T_919; // @[Mux.scala 27:72:freechips.rocketchip.system.DefaultRV32Config.fir@199712.4]
  assign _T_933 = _T_932 | _T_920; // @[Mux.scala 27:72:freechips.rocketchip.system.DefaultRV32Config.fir@199713.4]
  assign _T_934 = _T_933 | _T_921; // @[Mux.scala 27:72:freechips.rocketchip.system.DefaultRV32Config.fir@199714.4]
  assign _T_935 = _T_934 | _T_922; // @[Mux.scala 27:72:freechips.rocketchip.system.DefaultRV32Config.fir@199715.4]
  assign _T_936 = _T_935 | _T_923; // @[Mux.scala 27:72:freechips.rocketchip.system.DefaultRV32Config.fir@199716.4]
  assign ppn = _T_936 | _T_924; // @[Mux.scala 27:72:freechips.rocketchip.system.DefaultRV32Config.fir@199717.4]
  assign _T_938 = ~invalidate_refill; // @[TLB.scala 217:22:freechips.rocketchip.system.DefaultRV32Config.fir@199720.4]
  assign _T_939 = io_ptw_resp_valid & _T_938; // @[TLB.scala 217:19:freechips.rocketchip.system.DefaultRV32Config.fir@199721.4]
  assign _T_941 = io_ptw_resp_bits_pte_g & io_ptw_resp_bits_pte_v; // @[TLB.scala 223:25:freechips.rocketchip.system.DefaultRV32Config.fir@199728.6]
  assign _T_942 = ~io_ptw_resp_bits_pte_w; // @[PTW.scala 69:47:freechips.rocketchip.system.DefaultRV32Config.fir@199731.6]
  assign _T_943 = io_ptw_resp_bits_pte_x & _T_942; // @[PTW.scala 69:44:freechips.rocketchip.system.DefaultRV32Config.fir@199732.6]
  assign _T_944 = io_ptw_resp_bits_pte_r | _T_943; // @[PTW.scala 69:38:freechips.rocketchip.system.DefaultRV32Config.fir@199733.6]
  assign _T_945 = io_ptw_resp_bits_pte_v & _T_944; // @[PTW.scala 69:32:freechips.rocketchip.system.DefaultRV32Config.fir@199734.6]
  assign _T_946 = _T_945 & io_ptw_resp_bits_pte_a; // @[PTW.scala 69:52:freechips.rocketchip.system.DefaultRV32Config.fir@199735.6]
  assign _T_947 = _T_946 & io_ptw_resp_bits_pte_r; // @[PTW.scala 73:35:freechips.rocketchip.system.DefaultRV32Config.fir@199736.6]
  assign _T_953 = _T_946 & io_ptw_resp_bits_pte_w; // @[PTW.scala 74:35:freechips.rocketchip.system.DefaultRV32Config.fir@199743.6]
  assign _T_954 = _T_953 & io_ptw_resp_bits_pte_d; // @[PTW.scala 74:40:freechips.rocketchip.system.DefaultRV32Config.fir@199744.6]
  assign _T_960 = _T_946 & io_ptw_resp_bits_pte_x; // @[PTW.scala 75:35:freechips.rocketchip.system.DefaultRV32Config.fir@199751.6]
  assign _T_961 = ~io_ptw_resp_bits_homogeneous; // @[TLB.scala 237:37:freechips.rocketchip.system.DefaultRV32Config.fir@199761.6]
  assign _T_970 = {prot_x,prot_r,_T_232,prot_al,prot_al,prot_eff,cacheable,1'h0}; // @[TLB.scala 123:24:freechips.rocketchip.system.DefaultRV32Config.fir@199774.8]
  assign _T_978 = {refill_ppn,io_ptw_resp_bits_pte_u,_T_941,io_ptw_resp_bits_ae,_T_954,_T_960,_T_947,prot_w,_T_970}; // @[TLB.scala 123:24:freechips.rocketchip.system.DefaultRV32Config.fir@199782.8]
  assign _T_979 = io_ptw_resp_bits_level < 1'h1; // @[TLB.scala 239:40:freechips.rocketchip.system.DefaultRV32Config.fir@199786.8]
  assign _T_980 = r_superpage_repl_addr == 2'h0; // @[TLB.scala 240:82:freechips.rocketchip.system.DefaultRV32Config.fir@199788.10]
  assign _GEN_66 = _T_980 | superpage_entries_0_valid_0; // @[TLB.scala 240:89:freechips.rocketchip.system.DefaultRV32Config.fir@199789.10]
  assign _T_996 = r_superpage_repl_addr == 2'h1; // @[TLB.scala 240:82:freechips.rocketchip.system.DefaultRV32Config.fir@199810.10]
  assign _GEN_70 = _T_996 | superpage_entries_1_valid_0; // @[TLB.scala 240:89:freechips.rocketchip.system.DefaultRV32Config.fir@199811.10]
  assign _T_1012 = r_superpage_repl_addr == 2'h2; // @[TLB.scala 240:82:freechips.rocketchip.system.DefaultRV32Config.fir@199832.10]
  assign _GEN_74 = _T_1012 | superpage_entries_2_valid_0; // @[TLB.scala 240:89:freechips.rocketchip.system.DefaultRV32Config.fir@199833.10]
  assign _T_1028 = r_superpage_repl_addr == 2'h3; // @[TLB.scala 240:82:freechips.rocketchip.system.DefaultRV32Config.fir@199854.10]
  assign _GEN_78 = _T_1028 | superpage_entries_3_valid_0; // @[TLB.scala 240:89:freechips.rocketchip.system.DefaultRV32Config.fir@199855.10]
  assign _T_1044 = r_sectored_hit ? r_sectored_hit_addr : r_sectored_repl_addr; // @[TLB.scala 244:22:freechips.rocketchip.system.DefaultRV32Config.fir@199878.10]
  assign _T_1045 = _T_1044 == 3'h0; // @[TLB.scala 245:65:freechips.rocketchip.system.DefaultRV32Config.fir@199879.10]
  assign _T_1046 = ~r_sectored_hit; // @[TLB.scala 246:15:freechips.rocketchip.system.DefaultRV32Config.fir@199881.12]
  assign _GEN_80 = _T_1046 ? 1'h0 : sectored_entries_0_valid_0; // @[TLB.scala 246:32:freechips.rocketchip.system.DefaultRV32Config.fir@199882.12]
  assign _GEN_81 = _T_1046 ? 1'h0 : sectored_entries_0_valid_1; // @[TLB.scala 246:32:freechips.rocketchip.system.DefaultRV32Config.fir@199882.12]
  assign _GEN_82 = _T_1046 ? 1'h0 : sectored_entries_0_valid_2; // @[TLB.scala 246:32:freechips.rocketchip.system.DefaultRV32Config.fir@199882.12]
  assign _GEN_83 = _T_1046 ? 1'h0 : sectored_entries_0_valid_3; // @[TLB.scala 246:32:freechips.rocketchip.system.DefaultRV32Config.fir@199882.12]
  assign _GEN_950 = 2'h0 == r_refill_tag[1:0]; // @[TLB.scala 122:16:freechips.rocketchip.system.DefaultRV32Config.fir@199891.12]
  assign _GEN_84 = _GEN_950 | _GEN_80; // @[TLB.scala 122:16:freechips.rocketchip.system.DefaultRV32Config.fir@199891.12]
  assign _GEN_951 = 2'h1 == r_refill_tag[1:0]; // @[TLB.scala 122:16:freechips.rocketchip.system.DefaultRV32Config.fir@199891.12]
  assign _GEN_85 = _GEN_951 | _GEN_81; // @[TLB.scala 122:16:freechips.rocketchip.system.DefaultRV32Config.fir@199891.12]
  assign _GEN_952 = 2'h2 == r_refill_tag[1:0]; // @[TLB.scala 122:16:freechips.rocketchip.system.DefaultRV32Config.fir@199891.12]
  assign _GEN_86 = _GEN_952 | _GEN_82; // @[TLB.scala 122:16:freechips.rocketchip.system.DefaultRV32Config.fir@199891.12]
  assign _GEN_953 = 2'h3 == r_refill_tag[1:0]; // @[TLB.scala 122:16:freechips.rocketchip.system.DefaultRV32Config.fir@199891.12]
  assign _GEN_87 = _GEN_953 | _GEN_83; // @[TLB.scala 122:16:freechips.rocketchip.system.DefaultRV32Config.fir@199891.12]
  assign _GEN_92 = _T_1045 ? _GEN_84 : sectored_entries_0_valid_0; // @[TLB.scala 245:72:freechips.rocketchip.system.DefaultRV32Config.fir@199880.10]
  assign _GEN_93 = _T_1045 ? _GEN_85 : sectored_entries_0_valid_1; // @[TLB.scala 245:72:freechips.rocketchip.system.DefaultRV32Config.fir@199880.10]
  assign _GEN_94 = _T_1045 ? _GEN_86 : sectored_entries_0_valid_2; // @[TLB.scala 245:72:freechips.rocketchip.system.DefaultRV32Config.fir@199880.10]
  assign _GEN_95 = _T_1045 ? _GEN_87 : sectored_entries_0_valid_3; // @[TLB.scala 245:72:freechips.rocketchip.system.DefaultRV32Config.fir@199880.10]
  assign _T_1063 = _T_1044 == 3'h1; // @[TLB.scala 245:65:freechips.rocketchip.system.DefaultRV32Config.fir@199909.10]
  assign _GEN_102 = _T_1046 ? 1'h0 : sectored_entries_1_valid_0; // @[TLB.scala 246:32:freechips.rocketchip.system.DefaultRV32Config.fir@199912.12]
  assign _GEN_103 = _T_1046 ? 1'h0 : sectored_entries_1_valid_1; // @[TLB.scala 246:32:freechips.rocketchip.system.DefaultRV32Config.fir@199912.12]
  assign _GEN_104 = _T_1046 ? 1'h0 : sectored_entries_1_valid_2; // @[TLB.scala 246:32:freechips.rocketchip.system.DefaultRV32Config.fir@199912.12]
  assign _GEN_105 = _T_1046 ? 1'h0 : sectored_entries_1_valid_3; // @[TLB.scala 246:32:freechips.rocketchip.system.DefaultRV32Config.fir@199912.12]
  assign _GEN_106 = _GEN_950 | _GEN_102; // @[TLB.scala 122:16:freechips.rocketchip.system.DefaultRV32Config.fir@199921.12]
  assign _GEN_107 = _GEN_951 | _GEN_103; // @[TLB.scala 122:16:freechips.rocketchip.system.DefaultRV32Config.fir@199921.12]
  assign _GEN_108 = _GEN_952 | _GEN_104; // @[TLB.scala 122:16:freechips.rocketchip.system.DefaultRV32Config.fir@199921.12]
  assign _GEN_109 = _GEN_953 | _GEN_105; // @[TLB.scala 122:16:freechips.rocketchip.system.DefaultRV32Config.fir@199921.12]
  assign _GEN_114 = _T_1063 ? _GEN_106 : sectored_entries_1_valid_0; // @[TLB.scala 245:72:freechips.rocketchip.system.DefaultRV32Config.fir@199910.10]
  assign _GEN_115 = _T_1063 ? _GEN_107 : sectored_entries_1_valid_1; // @[TLB.scala 245:72:freechips.rocketchip.system.DefaultRV32Config.fir@199910.10]
  assign _GEN_116 = _T_1063 ? _GEN_108 : sectored_entries_1_valid_2; // @[TLB.scala 245:72:freechips.rocketchip.system.DefaultRV32Config.fir@199910.10]
  assign _GEN_117 = _T_1063 ? _GEN_109 : sectored_entries_1_valid_3; // @[TLB.scala 245:72:freechips.rocketchip.system.DefaultRV32Config.fir@199910.10]
  assign _T_1081 = _T_1044 == 3'h2; // @[TLB.scala 245:65:freechips.rocketchip.system.DefaultRV32Config.fir@199939.10]
  assign _GEN_124 = _T_1046 ? 1'h0 : sectored_entries_2_valid_0; // @[TLB.scala 246:32:freechips.rocketchip.system.DefaultRV32Config.fir@199942.12]
  assign _GEN_125 = _T_1046 ? 1'h0 : sectored_entries_2_valid_1; // @[TLB.scala 246:32:freechips.rocketchip.system.DefaultRV32Config.fir@199942.12]
  assign _GEN_126 = _T_1046 ? 1'h0 : sectored_entries_2_valid_2; // @[TLB.scala 246:32:freechips.rocketchip.system.DefaultRV32Config.fir@199942.12]
  assign _GEN_127 = _T_1046 ? 1'h0 : sectored_entries_2_valid_3; // @[TLB.scala 246:32:freechips.rocketchip.system.DefaultRV32Config.fir@199942.12]
  assign _GEN_128 = _GEN_950 | _GEN_124; // @[TLB.scala 122:16:freechips.rocketchip.system.DefaultRV32Config.fir@199951.12]
  assign _GEN_129 = _GEN_951 | _GEN_125; // @[TLB.scala 122:16:freechips.rocketchip.system.DefaultRV32Config.fir@199951.12]
  assign _GEN_130 = _GEN_952 | _GEN_126; // @[TLB.scala 122:16:freechips.rocketchip.system.DefaultRV32Config.fir@199951.12]
  assign _GEN_131 = _GEN_953 | _GEN_127; // @[TLB.scala 122:16:freechips.rocketchip.system.DefaultRV32Config.fir@199951.12]
  assign _GEN_136 = _T_1081 ? _GEN_128 : sectored_entries_2_valid_0; // @[TLB.scala 245:72:freechips.rocketchip.system.DefaultRV32Config.fir@199940.10]
  assign _GEN_137 = _T_1081 ? _GEN_129 : sectored_entries_2_valid_1; // @[TLB.scala 245:72:freechips.rocketchip.system.DefaultRV32Config.fir@199940.10]
  assign _GEN_138 = _T_1081 ? _GEN_130 : sectored_entries_2_valid_2; // @[TLB.scala 245:72:freechips.rocketchip.system.DefaultRV32Config.fir@199940.10]
  assign _GEN_139 = _T_1081 ? _GEN_131 : sectored_entries_2_valid_3; // @[TLB.scala 245:72:freechips.rocketchip.system.DefaultRV32Config.fir@199940.10]
  assign _T_1099 = _T_1044 == 3'h3; // @[TLB.scala 245:65:freechips.rocketchip.system.DefaultRV32Config.fir@199969.10]
  assign _GEN_146 = _T_1046 ? 1'h0 : sectored_entries_3_valid_0; // @[TLB.scala 246:32:freechips.rocketchip.system.DefaultRV32Config.fir@199972.12]
  assign _GEN_147 = _T_1046 ? 1'h0 : sectored_entries_3_valid_1; // @[TLB.scala 246:32:freechips.rocketchip.system.DefaultRV32Config.fir@199972.12]
  assign _GEN_148 = _T_1046 ? 1'h0 : sectored_entries_3_valid_2; // @[TLB.scala 246:32:freechips.rocketchip.system.DefaultRV32Config.fir@199972.12]
  assign _GEN_149 = _T_1046 ? 1'h0 : sectored_entries_3_valid_3; // @[TLB.scala 246:32:freechips.rocketchip.system.DefaultRV32Config.fir@199972.12]
  assign _GEN_150 = _GEN_950 | _GEN_146; // @[TLB.scala 122:16:freechips.rocketchip.system.DefaultRV32Config.fir@199981.12]
  assign _GEN_151 = _GEN_951 | _GEN_147; // @[TLB.scala 122:16:freechips.rocketchip.system.DefaultRV32Config.fir@199981.12]
  assign _GEN_152 = _GEN_952 | _GEN_148; // @[TLB.scala 122:16:freechips.rocketchip.system.DefaultRV32Config.fir@199981.12]
  assign _GEN_153 = _GEN_953 | _GEN_149; // @[TLB.scala 122:16:freechips.rocketchip.system.DefaultRV32Config.fir@199981.12]
  assign _GEN_158 = _T_1099 ? _GEN_150 : sectored_entries_3_valid_0; // @[TLB.scala 245:72:freechips.rocketchip.system.DefaultRV32Config.fir@199970.10]
  assign _GEN_159 = _T_1099 ? _GEN_151 : sectored_entries_3_valid_1; // @[TLB.scala 245:72:freechips.rocketchip.system.DefaultRV32Config.fir@199970.10]
  assign _GEN_160 = _T_1099 ? _GEN_152 : sectored_entries_3_valid_2; // @[TLB.scala 245:72:freechips.rocketchip.system.DefaultRV32Config.fir@199970.10]
  assign _GEN_161 = _T_1099 ? _GEN_153 : sectored_entries_3_valid_3; // @[TLB.scala 245:72:freechips.rocketchip.system.DefaultRV32Config.fir@199970.10]
  assign _T_1117 = _T_1044 == 3'h4; // @[TLB.scala 245:65:freechips.rocketchip.system.DefaultRV32Config.fir@199999.10]
  assign _GEN_168 = _T_1046 ? 1'h0 : sectored_entries_4_valid_0; // @[TLB.scala 246:32:freechips.rocketchip.system.DefaultRV32Config.fir@200002.12]
  assign _GEN_169 = _T_1046 ? 1'h0 : sectored_entries_4_valid_1; // @[TLB.scala 246:32:freechips.rocketchip.system.DefaultRV32Config.fir@200002.12]
  assign _GEN_170 = _T_1046 ? 1'h0 : sectored_entries_4_valid_2; // @[TLB.scala 246:32:freechips.rocketchip.system.DefaultRV32Config.fir@200002.12]
  assign _GEN_171 = _T_1046 ? 1'h0 : sectored_entries_4_valid_3; // @[TLB.scala 246:32:freechips.rocketchip.system.DefaultRV32Config.fir@200002.12]
  assign _GEN_172 = _GEN_950 | _GEN_168; // @[TLB.scala 122:16:freechips.rocketchip.system.DefaultRV32Config.fir@200011.12]
  assign _GEN_173 = _GEN_951 | _GEN_169; // @[TLB.scala 122:16:freechips.rocketchip.system.DefaultRV32Config.fir@200011.12]
  assign _GEN_174 = _GEN_952 | _GEN_170; // @[TLB.scala 122:16:freechips.rocketchip.system.DefaultRV32Config.fir@200011.12]
  assign _GEN_175 = _GEN_953 | _GEN_171; // @[TLB.scala 122:16:freechips.rocketchip.system.DefaultRV32Config.fir@200011.12]
  assign _GEN_180 = _T_1117 ? _GEN_172 : sectored_entries_4_valid_0; // @[TLB.scala 245:72:freechips.rocketchip.system.DefaultRV32Config.fir@200000.10]
  assign _GEN_181 = _T_1117 ? _GEN_173 : sectored_entries_4_valid_1; // @[TLB.scala 245:72:freechips.rocketchip.system.DefaultRV32Config.fir@200000.10]
  assign _GEN_182 = _T_1117 ? _GEN_174 : sectored_entries_4_valid_2; // @[TLB.scala 245:72:freechips.rocketchip.system.DefaultRV32Config.fir@200000.10]
  assign _GEN_183 = _T_1117 ? _GEN_175 : sectored_entries_4_valid_3; // @[TLB.scala 245:72:freechips.rocketchip.system.DefaultRV32Config.fir@200000.10]
  assign _T_1135 = _T_1044 == 3'h5; // @[TLB.scala 245:65:freechips.rocketchip.system.DefaultRV32Config.fir@200029.10]
  assign _GEN_190 = _T_1046 ? 1'h0 : sectored_entries_5_valid_0; // @[TLB.scala 246:32:freechips.rocketchip.system.DefaultRV32Config.fir@200032.12]
  assign _GEN_191 = _T_1046 ? 1'h0 : sectored_entries_5_valid_1; // @[TLB.scala 246:32:freechips.rocketchip.system.DefaultRV32Config.fir@200032.12]
  assign _GEN_192 = _T_1046 ? 1'h0 : sectored_entries_5_valid_2; // @[TLB.scala 246:32:freechips.rocketchip.system.DefaultRV32Config.fir@200032.12]
  assign _GEN_193 = _T_1046 ? 1'h0 : sectored_entries_5_valid_3; // @[TLB.scala 246:32:freechips.rocketchip.system.DefaultRV32Config.fir@200032.12]
  assign _GEN_194 = _GEN_950 | _GEN_190; // @[TLB.scala 122:16:freechips.rocketchip.system.DefaultRV32Config.fir@200041.12]
  assign _GEN_195 = _GEN_951 | _GEN_191; // @[TLB.scala 122:16:freechips.rocketchip.system.DefaultRV32Config.fir@200041.12]
  assign _GEN_196 = _GEN_952 | _GEN_192; // @[TLB.scala 122:16:freechips.rocketchip.system.DefaultRV32Config.fir@200041.12]
  assign _GEN_197 = _GEN_953 | _GEN_193; // @[TLB.scala 122:16:freechips.rocketchip.system.DefaultRV32Config.fir@200041.12]
  assign _GEN_202 = _T_1135 ? _GEN_194 : sectored_entries_5_valid_0; // @[TLB.scala 245:72:freechips.rocketchip.system.DefaultRV32Config.fir@200030.10]
  assign _GEN_203 = _T_1135 ? _GEN_195 : sectored_entries_5_valid_1; // @[TLB.scala 245:72:freechips.rocketchip.system.DefaultRV32Config.fir@200030.10]
  assign _GEN_204 = _T_1135 ? _GEN_196 : sectored_entries_5_valid_2; // @[TLB.scala 245:72:freechips.rocketchip.system.DefaultRV32Config.fir@200030.10]
  assign _GEN_205 = _T_1135 ? _GEN_197 : sectored_entries_5_valid_3; // @[TLB.scala 245:72:freechips.rocketchip.system.DefaultRV32Config.fir@200030.10]
  assign _T_1153 = _T_1044 == 3'h6; // @[TLB.scala 245:65:freechips.rocketchip.system.DefaultRV32Config.fir@200059.10]
  assign _GEN_212 = _T_1046 ? 1'h0 : sectored_entries_6_valid_0; // @[TLB.scala 246:32:freechips.rocketchip.system.DefaultRV32Config.fir@200062.12]
  assign _GEN_213 = _T_1046 ? 1'h0 : sectored_entries_6_valid_1; // @[TLB.scala 246:32:freechips.rocketchip.system.DefaultRV32Config.fir@200062.12]
  assign _GEN_214 = _T_1046 ? 1'h0 : sectored_entries_6_valid_2; // @[TLB.scala 246:32:freechips.rocketchip.system.DefaultRV32Config.fir@200062.12]
  assign _GEN_215 = _T_1046 ? 1'h0 : sectored_entries_6_valid_3; // @[TLB.scala 246:32:freechips.rocketchip.system.DefaultRV32Config.fir@200062.12]
  assign _GEN_216 = _GEN_950 | _GEN_212; // @[TLB.scala 122:16:freechips.rocketchip.system.DefaultRV32Config.fir@200071.12]
  assign _GEN_217 = _GEN_951 | _GEN_213; // @[TLB.scala 122:16:freechips.rocketchip.system.DefaultRV32Config.fir@200071.12]
  assign _GEN_218 = _GEN_952 | _GEN_214; // @[TLB.scala 122:16:freechips.rocketchip.system.DefaultRV32Config.fir@200071.12]
  assign _GEN_219 = _GEN_953 | _GEN_215; // @[TLB.scala 122:16:freechips.rocketchip.system.DefaultRV32Config.fir@200071.12]
  assign _GEN_224 = _T_1153 ? _GEN_216 : sectored_entries_6_valid_0; // @[TLB.scala 245:72:freechips.rocketchip.system.DefaultRV32Config.fir@200060.10]
  assign _GEN_225 = _T_1153 ? _GEN_217 : sectored_entries_6_valid_1; // @[TLB.scala 245:72:freechips.rocketchip.system.DefaultRV32Config.fir@200060.10]
  assign _GEN_226 = _T_1153 ? _GEN_218 : sectored_entries_6_valid_2; // @[TLB.scala 245:72:freechips.rocketchip.system.DefaultRV32Config.fir@200060.10]
  assign _GEN_227 = _T_1153 ? _GEN_219 : sectored_entries_6_valid_3; // @[TLB.scala 245:72:freechips.rocketchip.system.DefaultRV32Config.fir@200060.10]
  assign _T_1171 = _T_1044 == 3'h7; // @[TLB.scala 245:65:freechips.rocketchip.system.DefaultRV32Config.fir@200089.10]
  assign _GEN_234 = _T_1046 ? 1'h0 : sectored_entries_7_valid_0; // @[TLB.scala 246:32:freechips.rocketchip.system.DefaultRV32Config.fir@200092.12]
  assign _GEN_235 = _T_1046 ? 1'h0 : sectored_entries_7_valid_1; // @[TLB.scala 246:32:freechips.rocketchip.system.DefaultRV32Config.fir@200092.12]
  assign _GEN_236 = _T_1046 ? 1'h0 : sectored_entries_7_valid_2; // @[TLB.scala 246:32:freechips.rocketchip.system.DefaultRV32Config.fir@200092.12]
  assign _GEN_237 = _T_1046 ? 1'h0 : sectored_entries_7_valid_3; // @[TLB.scala 246:32:freechips.rocketchip.system.DefaultRV32Config.fir@200092.12]
  assign _GEN_238 = _GEN_950 | _GEN_234; // @[TLB.scala 122:16:freechips.rocketchip.system.DefaultRV32Config.fir@200101.12]
  assign _GEN_239 = _GEN_951 | _GEN_235; // @[TLB.scala 122:16:freechips.rocketchip.system.DefaultRV32Config.fir@200101.12]
  assign _GEN_240 = _GEN_952 | _GEN_236; // @[TLB.scala 122:16:freechips.rocketchip.system.DefaultRV32Config.fir@200101.12]
  assign _GEN_241 = _GEN_953 | _GEN_237; // @[TLB.scala 122:16:freechips.rocketchip.system.DefaultRV32Config.fir@200101.12]
  assign _GEN_246 = _T_1171 ? _GEN_238 : sectored_entries_7_valid_0; // @[TLB.scala 245:72:freechips.rocketchip.system.DefaultRV32Config.fir@200090.10]
  assign _GEN_247 = _T_1171 ? _GEN_239 : sectored_entries_7_valid_1; // @[TLB.scala 245:72:freechips.rocketchip.system.DefaultRV32Config.fir@200090.10]
  assign _GEN_248 = _T_1171 ? _GEN_240 : sectored_entries_7_valid_2; // @[TLB.scala 245:72:freechips.rocketchip.system.DefaultRV32Config.fir@200090.10]
  assign _GEN_249 = _T_1171 ? _GEN_241 : sectored_entries_7_valid_3; // @[TLB.scala 245:72:freechips.rocketchip.system.DefaultRV32Config.fir@200090.10]
  assign _GEN_258 = _T_979 ? _GEN_66 : superpage_entries_0_valid_0; // @[TLB.scala 239:54:freechips.rocketchip.system.DefaultRV32Config.fir@199787.8]
  assign _GEN_262 = _T_979 ? _GEN_70 : superpage_entries_1_valid_0; // @[TLB.scala 239:54:freechips.rocketchip.system.DefaultRV32Config.fir@199787.8]
  assign _GEN_266 = _T_979 ? _GEN_74 : superpage_entries_2_valid_0; // @[TLB.scala 239:54:freechips.rocketchip.system.DefaultRV32Config.fir@199787.8]
  assign _GEN_270 = _T_979 ? _GEN_78 : superpage_entries_3_valid_0; // @[TLB.scala 239:54:freechips.rocketchip.system.DefaultRV32Config.fir@199787.8]
  assign _GEN_272 = _T_979 ? sectored_entries_0_valid_0 : _GEN_92; // @[TLB.scala 239:54:freechips.rocketchip.system.DefaultRV32Config.fir@199787.8]
  assign _GEN_273 = _T_979 ? sectored_entries_0_valid_1 : _GEN_93; // @[TLB.scala 239:54:freechips.rocketchip.system.DefaultRV32Config.fir@199787.8]
  assign _GEN_274 = _T_979 ? sectored_entries_0_valid_2 : _GEN_94; // @[TLB.scala 239:54:freechips.rocketchip.system.DefaultRV32Config.fir@199787.8]
  assign _GEN_275 = _T_979 ? sectored_entries_0_valid_3 : _GEN_95; // @[TLB.scala 239:54:freechips.rocketchip.system.DefaultRV32Config.fir@199787.8]
  assign _GEN_282 = _T_979 ? sectored_entries_1_valid_0 : _GEN_114; // @[TLB.scala 239:54:freechips.rocketchip.system.DefaultRV32Config.fir@199787.8]
  assign _GEN_283 = _T_979 ? sectored_entries_1_valid_1 : _GEN_115; // @[TLB.scala 239:54:freechips.rocketchip.system.DefaultRV32Config.fir@199787.8]
  assign _GEN_284 = _T_979 ? sectored_entries_1_valid_2 : _GEN_116; // @[TLB.scala 239:54:freechips.rocketchip.system.DefaultRV32Config.fir@199787.8]
  assign _GEN_285 = _T_979 ? sectored_entries_1_valid_3 : _GEN_117; // @[TLB.scala 239:54:freechips.rocketchip.system.DefaultRV32Config.fir@199787.8]
  assign _GEN_292 = _T_979 ? sectored_entries_2_valid_0 : _GEN_136; // @[TLB.scala 239:54:freechips.rocketchip.system.DefaultRV32Config.fir@199787.8]
  assign _GEN_293 = _T_979 ? sectored_entries_2_valid_1 : _GEN_137; // @[TLB.scala 239:54:freechips.rocketchip.system.DefaultRV32Config.fir@199787.8]
  assign _GEN_294 = _T_979 ? sectored_entries_2_valid_2 : _GEN_138; // @[TLB.scala 239:54:freechips.rocketchip.system.DefaultRV32Config.fir@199787.8]
  assign _GEN_295 = _T_979 ? sectored_entries_2_valid_3 : _GEN_139; // @[TLB.scala 239:54:freechips.rocketchip.system.DefaultRV32Config.fir@199787.8]
  assign _GEN_302 = _T_979 ? sectored_entries_3_valid_0 : _GEN_158; // @[TLB.scala 239:54:freechips.rocketchip.system.DefaultRV32Config.fir@199787.8]
  assign _GEN_303 = _T_979 ? sectored_entries_3_valid_1 : _GEN_159; // @[TLB.scala 239:54:freechips.rocketchip.system.DefaultRV32Config.fir@199787.8]
  assign _GEN_304 = _T_979 ? sectored_entries_3_valid_2 : _GEN_160; // @[TLB.scala 239:54:freechips.rocketchip.system.DefaultRV32Config.fir@199787.8]
  assign _GEN_305 = _T_979 ? sectored_entries_3_valid_3 : _GEN_161; // @[TLB.scala 239:54:freechips.rocketchip.system.DefaultRV32Config.fir@199787.8]
  assign _GEN_312 = _T_979 ? sectored_entries_4_valid_0 : _GEN_180; // @[TLB.scala 239:54:freechips.rocketchip.system.DefaultRV32Config.fir@199787.8]
  assign _GEN_313 = _T_979 ? sectored_entries_4_valid_1 : _GEN_181; // @[TLB.scala 239:54:freechips.rocketchip.system.DefaultRV32Config.fir@199787.8]
  assign _GEN_314 = _T_979 ? sectored_entries_4_valid_2 : _GEN_182; // @[TLB.scala 239:54:freechips.rocketchip.system.DefaultRV32Config.fir@199787.8]
  assign _GEN_315 = _T_979 ? sectored_entries_4_valid_3 : _GEN_183; // @[TLB.scala 239:54:freechips.rocketchip.system.DefaultRV32Config.fir@199787.8]
  assign _GEN_322 = _T_979 ? sectored_entries_5_valid_0 : _GEN_202; // @[TLB.scala 239:54:freechips.rocketchip.system.DefaultRV32Config.fir@199787.8]
  assign _GEN_323 = _T_979 ? sectored_entries_5_valid_1 : _GEN_203; // @[TLB.scala 239:54:freechips.rocketchip.system.DefaultRV32Config.fir@199787.8]
  assign _GEN_324 = _T_979 ? sectored_entries_5_valid_2 : _GEN_204; // @[TLB.scala 239:54:freechips.rocketchip.system.DefaultRV32Config.fir@199787.8]
  assign _GEN_325 = _T_979 ? sectored_entries_5_valid_3 : _GEN_205; // @[TLB.scala 239:54:freechips.rocketchip.system.DefaultRV32Config.fir@199787.8]
  assign _GEN_332 = _T_979 ? sectored_entries_6_valid_0 : _GEN_224; // @[TLB.scala 239:54:freechips.rocketchip.system.DefaultRV32Config.fir@199787.8]
  assign _GEN_333 = _T_979 ? sectored_entries_6_valid_1 : _GEN_225; // @[TLB.scala 239:54:freechips.rocketchip.system.DefaultRV32Config.fir@199787.8]
  assign _GEN_334 = _T_979 ? sectored_entries_6_valid_2 : _GEN_226; // @[TLB.scala 239:54:freechips.rocketchip.system.DefaultRV32Config.fir@199787.8]
  assign _GEN_335 = _T_979 ? sectored_entries_6_valid_3 : _GEN_227; // @[TLB.scala 239:54:freechips.rocketchip.system.DefaultRV32Config.fir@199787.8]
  assign _GEN_342 = _T_979 ? sectored_entries_7_valid_0 : _GEN_246; // @[TLB.scala 239:54:freechips.rocketchip.system.DefaultRV32Config.fir@199787.8]
  assign _GEN_343 = _T_979 ? sectored_entries_7_valid_1 : _GEN_247; // @[TLB.scala 239:54:freechips.rocketchip.system.DefaultRV32Config.fir@199787.8]
  assign _GEN_344 = _T_979 ? sectored_entries_7_valid_2 : _GEN_248; // @[TLB.scala 239:54:freechips.rocketchip.system.DefaultRV32Config.fir@199787.8]
  assign _GEN_345 = _T_979 ? sectored_entries_7_valid_3 : _GEN_249; // @[TLB.scala 239:54:freechips.rocketchip.system.DefaultRV32Config.fir@199787.8]
  assign _GEN_354 = _T_961 | special_entry_valid_0; // @[TLB.scala 237:68:freechips.rocketchip.system.DefaultRV32Config.fir@199763.6]
  assign _GEN_358 = _T_961 ? superpage_entries_0_valid_0 : _GEN_258; // @[TLB.scala 237:68:freechips.rocketchip.system.DefaultRV32Config.fir@199763.6]
  assign _GEN_362 = _T_961 ? superpage_entries_1_valid_0 : _GEN_262; // @[TLB.scala 237:68:freechips.rocketchip.system.DefaultRV32Config.fir@199763.6]
  assign _GEN_366 = _T_961 ? superpage_entries_2_valid_0 : _GEN_266; // @[TLB.scala 237:68:freechips.rocketchip.system.DefaultRV32Config.fir@199763.6]
  assign _GEN_370 = _T_961 ? superpage_entries_3_valid_0 : _GEN_270; // @[TLB.scala 237:68:freechips.rocketchip.system.DefaultRV32Config.fir@199763.6]
  assign _GEN_372 = _T_961 ? sectored_entries_0_valid_0 : _GEN_272; // @[TLB.scala 237:68:freechips.rocketchip.system.DefaultRV32Config.fir@199763.6]
  assign _GEN_373 = _T_961 ? sectored_entries_0_valid_1 : _GEN_273; // @[TLB.scala 237:68:freechips.rocketchip.system.DefaultRV32Config.fir@199763.6]
  assign _GEN_374 = _T_961 ? sectored_entries_0_valid_2 : _GEN_274; // @[TLB.scala 237:68:freechips.rocketchip.system.DefaultRV32Config.fir@199763.6]
  assign _GEN_375 = _T_961 ? sectored_entries_0_valid_3 : _GEN_275; // @[TLB.scala 237:68:freechips.rocketchip.system.DefaultRV32Config.fir@199763.6]
  assign _GEN_382 = _T_961 ? sectored_entries_1_valid_0 : _GEN_282; // @[TLB.scala 237:68:freechips.rocketchip.system.DefaultRV32Config.fir@199763.6]
  assign _GEN_383 = _T_961 ? sectored_entries_1_valid_1 : _GEN_283; // @[TLB.scala 237:68:freechips.rocketchip.system.DefaultRV32Config.fir@199763.6]
  assign _GEN_384 = _T_961 ? sectored_entries_1_valid_2 : _GEN_284; // @[TLB.scala 237:68:freechips.rocketchip.system.DefaultRV32Config.fir@199763.6]
  assign _GEN_385 = _T_961 ? sectored_entries_1_valid_3 : _GEN_285; // @[TLB.scala 237:68:freechips.rocketchip.system.DefaultRV32Config.fir@199763.6]
  assign _GEN_392 = _T_961 ? sectored_entries_2_valid_0 : _GEN_292; // @[TLB.scala 237:68:freechips.rocketchip.system.DefaultRV32Config.fir@199763.6]
  assign _GEN_393 = _T_961 ? sectored_entries_2_valid_1 : _GEN_293; // @[TLB.scala 237:68:freechips.rocketchip.system.DefaultRV32Config.fir@199763.6]
  assign _GEN_394 = _T_961 ? sectored_entries_2_valid_2 : _GEN_294; // @[TLB.scala 237:68:freechips.rocketchip.system.DefaultRV32Config.fir@199763.6]
  assign _GEN_395 = _T_961 ? sectored_entries_2_valid_3 : _GEN_295; // @[TLB.scala 237:68:freechips.rocketchip.system.DefaultRV32Config.fir@199763.6]
  assign _GEN_402 = _T_961 ? sectored_entries_3_valid_0 : _GEN_302; // @[TLB.scala 237:68:freechips.rocketchip.system.DefaultRV32Config.fir@199763.6]
  assign _GEN_403 = _T_961 ? sectored_entries_3_valid_1 : _GEN_303; // @[TLB.scala 237:68:freechips.rocketchip.system.DefaultRV32Config.fir@199763.6]
  assign _GEN_404 = _T_961 ? sectored_entries_3_valid_2 : _GEN_304; // @[TLB.scala 237:68:freechips.rocketchip.system.DefaultRV32Config.fir@199763.6]
  assign _GEN_405 = _T_961 ? sectored_entries_3_valid_3 : _GEN_305; // @[TLB.scala 237:68:freechips.rocketchip.system.DefaultRV32Config.fir@199763.6]
  assign _GEN_412 = _T_961 ? sectored_entries_4_valid_0 : _GEN_312; // @[TLB.scala 237:68:freechips.rocketchip.system.DefaultRV32Config.fir@199763.6]
  assign _GEN_413 = _T_961 ? sectored_entries_4_valid_1 : _GEN_313; // @[TLB.scala 237:68:freechips.rocketchip.system.DefaultRV32Config.fir@199763.6]
  assign _GEN_414 = _T_961 ? sectored_entries_4_valid_2 : _GEN_314; // @[TLB.scala 237:68:freechips.rocketchip.system.DefaultRV32Config.fir@199763.6]
  assign _GEN_415 = _T_961 ? sectored_entries_4_valid_3 : _GEN_315; // @[TLB.scala 237:68:freechips.rocketchip.system.DefaultRV32Config.fir@199763.6]
  assign _GEN_422 = _T_961 ? sectored_entries_5_valid_0 : _GEN_322; // @[TLB.scala 237:68:freechips.rocketchip.system.DefaultRV32Config.fir@199763.6]
  assign _GEN_423 = _T_961 ? sectored_entries_5_valid_1 : _GEN_323; // @[TLB.scala 237:68:freechips.rocketchip.system.DefaultRV32Config.fir@199763.6]
  assign _GEN_424 = _T_961 ? sectored_entries_5_valid_2 : _GEN_324; // @[TLB.scala 237:68:freechips.rocketchip.system.DefaultRV32Config.fir@199763.6]
  assign _GEN_425 = _T_961 ? sectored_entries_5_valid_3 : _GEN_325; // @[TLB.scala 237:68:freechips.rocketchip.system.DefaultRV32Config.fir@199763.6]
  assign _GEN_432 = _T_961 ? sectored_entries_6_valid_0 : _GEN_332; // @[TLB.scala 237:68:freechips.rocketchip.system.DefaultRV32Config.fir@199763.6]
  assign _GEN_433 = _T_961 ? sectored_entries_6_valid_1 : _GEN_333; // @[TLB.scala 237:68:freechips.rocketchip.system.DefaultRV32Config.fir@199763.6]
  assign _GEN_434 = _T_961 ? sectored_entries_6_valid_2 : _GEN_334; // @[TLB.scala 237:68:freechips.rocketchip.system.DefaultRV32Config.fir@199763.6]
  assign _GEN_435 = _T_961 ? sectored_entries_6_valid_3 : _GEN_335; // @[TLB.scala 237:68:freechips.rocketchip.system.DefaultRV32Config.fir@199763.6]
  assign _GEN_442 = _T_961 ? sectored_entries_7_valid_0 : _GEN_342; // @[TLB.scala 237:68:freechips.rocketchip.system.DefaultRV32Config.fir@199763.6]
  assign _GEN_443 = _T_961 ? sectored_entries_7_valid_1 : _GEN_343; // @[TLB.scala 237:68:freechips.rocketchip.system.DefaultRV32Config.fir@199763.6]
  assign _GEN_444 = _T_961 ? sectored_entries_7_valid_2 : _GEN_344; // @[TLB.scala 237:68:freechips.rocketchip.system.DefaultRV32Config.fir@199763.6]
  assign _GEN_445 = _T_961 ? sectored_entries_7_valid_3 : _GEN_345; // @[TLB.scala 237:68:freechips.rocketchip.system.DefaultRV32Config.fir@199763.6]
  assign _GEN_454 = _T_939 ? _GEN_354 : special_entry_valid_0; // @[TLB.scala 217:42:freechips.rocketchip.system.DefaultRV32Config.fir@199722.4]
  assign _GEN_458 = _T_939 ? _GEN_358 : superpage_entries_0_valid_0; // @[TLB.scala 217:42:freechips.rocketchip.system.DefaultRV32Config.fir@199722.4]
  assign _GEN_462 = _T_939 ? _GEN_362 : superpage_entries_1_valid_0; // @[TLB.scala 217:42:freechips.rocketchip.system.DefaultRV32Config.fir@199722.4]
  assign _GEN_466 = _T_939 ? _GEN_366 : superpage_entries_2_valid_0; // @[TLB.scala 217:42:freechips.rocketchip.system.DefaultRV32Config.fir@199722.4]
  assign _GEN_470 = _T_939 ? _GEN_370 : superpage_entries_3_valid_0; // @[TLB.scala 217:42:freechips.rocketchip.system.DefaultRV32Config.fir@199722.4]
  assign _GEN_472 = _T_939 ? _GEN_372 : sectored_entries_0_valid_0; // @[TLB.scala 217:42:freechips.rocketchip.system.DefaultRV32Config.fir@199722.4]
  assign _GEN_473 = _T_939 ? _GEN_373 : sectored_entries_0_valid_1; // @[TLB.scala 217:42:freechips.rocketchip.system.DefaultRV32Config.fir@199722.4]
  assign _GEN_474 = _T_939 ? _GEN_374 : sectored_entries_0_valid_2; // @[TLB.scala 217:42:freechips.rocketchip.system.DefaultRV32Config.fir@199722.4]
  assign _GEN_475 = _T_939 ? _GEN_375 : sectored_entries_0_valid_3; // @[TLB.scala 217:42:freechips.rocketchip.system.DefaultRV32Config.fir@199722.4]
  assign _GEN_482 = _T_939 ? _GEN_382 : sectored_entries_1_valid_0; // @[TLB.scala 217:42:freechips.rocketchip.system.DefaultRV32Config.fir@199722.4]
  assign _GEN_483 = _T_939 ? _GEN_383 : sectored_entries_1_valid_1; // @[TLB.scala 217:42:freechips.rocketchip.system.DefaultRV32Config.fir@199722.4]
  assign _GEN_484 = _T_939 ? _GEN_384 : sectored_entries_1_valid_2; // @[TLB.scala 217:42:freechips.rocketchip.system.DefaultRV32Config.fir@199722.4]
  assign _GEN_485 = _T_939 ? _GEN_385 : sectored_entries_1_valid_3; // @[TLB.scala 217:42:freechips.rocketchip.system.DefaultRV32Config.fir@199722.4]
  assign _GEN_492 = _T_939 ? _GEN_392 : sectored_entries_2_valid_0; // @[TLB.scala 217:42:freechips.rocketchip.system.DefaultRV32Config.fir@199722.4]
  assign _GEN_493 = _T_939 ? _GEN_393 : sectored_entries_2_valid_1; // @[TLB.scala 217:42:freechips.rocketchip.system.DefaultRV32Config.fir@199722.4]
  assign _GEN_494 = _T_939 ? _GEN_394 : sectored_entries_2_valid_2; // @[TLB.scala 217:42:freechips.rocketchip.system.DefaultRV32Config.fir@199722.4]
  assign _GEN_495 = _T_939 ? _GEN_395 : sectored_entries_2_valid_3; // @[TLB.scala 217:42:freechips.rocketchip.system.DefaultRV32Config.fir@199722.4]
  assign _GEN_502 = _T_939 ? _GEN_402 : sectored_entries_3_valid_0; // @[TLB.scala 217:42:freechips.rocketchip.system.DefaultRV32Config.fir@199722.4]
  assign _GEN_503 = _T_939 ? _GEN_403 : sectored_entries_3_valid_1; // @[TLB.scala 217:42:freechips.rocketchip.system.DefaultRV32Config.fir@199722.4]
  assign _GEN_504 = _T_939 ? _GEN_404 : sectored_entries_3_valid_2; // @[TLB.scala 217:42:freechips.rocketchip.system.DefaultRV32Config.fir@199722.4]
  assign _GEN_505 = _T_939 ? _GEN_405 : sectored_entries_3_valid_3; // @[TLB.scala 217:42:freechips.rocketchip.system.DefaultRV32Config.fir@199722.4]
  assign _GEN_512 = _T_939 ? _GEN_412 : sectored_entries_4_valid_0; // @[TLB.scala 217:42:freechips.rocketchip.system.DefaultRV32Config.fir@199722.4]
  assign _GEN_513 = _T_939 ? _GEN_413 : sectored_entries_4_valid_1; // @[TLB.scala 217:42:freechips.rocketchip.system.DefaultRV32Config.fir@199722.4]
  assign _GEN_514 = _T_939 ? _GEN_414 : sectored_entries_4_valid_2; // @[TLB.scala 217:42:freechips.rocketchip.system.DefaultRV32Config.fir@199722.4]
  assign _GEN_515 = _T_939 ? _GEN_415 : sectored_entries_4_valid_3; // @[TLB.scala 217:42:freechips.rocketchip.system.DefaultRV32Config.fir@199722.4]
  assign _GEN_522 = _T_939 ? _GEN_422 : sectored_entries_5_valid_0; // @[TLB.scala 217:42:freechips.rocketchip.system.DefaultRV32Config.fir@199722.4]
  assign _GEN_523 = _T_939 ? _GEN_423 : sectored_entries_5_valid_1; // @[TLB.scala 217:42:freechips.rocketchip.system.DefaultRV32Config.fir@199722.4]
  assign _GEN_524 = _T_939 ? _GEN_424 : sectored_entries_5_valid_2; // @[TLB.scala 217:42:freechips.rocketchip.system.DefaultRV32Config.fir@199722.4]
  assign _GEN_525 = _T_939 ? _GEN_425 : sectored_entries_5_valid_3; // @[TLB.scala 217:42:freechips.rocketchip.system.DefaultRV32Config.fir@199722.4]
  assign _GEN_532 = _T_939 ? _GEN_432 : sectored_entries_6_valid_0; // @[TLB.scala 217:42:freechips.rocketchip.system.DefaultRV32Config.fir@199722.4]
  assign _GEN_533 = _T_939 ? _GEN_433 : sectored_entries_6_valid_1; // @[TLB.scala 217:42:freechips.rocketchip.system.DefaultRV32Config.fir@199722.4]
  assign _GEN_534 = _T_939 ? _GEN_434 : sectored_entries_6_valid_2; // @[TLB.scala 217:42:freechips.rocketchip.system.DefaultRV32Config.fir@199722.4]
  assign _GEN_535 = _T_939 ? _GEN_435 : sectored_entries_6_valid_3; // @[TLB.scala 217:42:freechips.rocketchip.system.DefaultRV32Config.fir@199722.4]
  assign _GEN_542 = _T_939 ? _GEN_442 : sectored_entries_7_valid_0; // @[TLB.scala 217:42:freechips.rocketchip.system.DefaultRV32Config.fir@199722.4]
  assign _GEN_543 = _T_939 ? _GEN_443 : sectored_entries_7_valid_1; // @[TLB.scala 217:42:freechips.rocketchip.system.DefaultRV32Config.fir@199722.4]
  assign _GEN_544 = _T_939 ? _GEN_444 : sectored_entries_7_valid_2; // @[TLB.scala 217:42:freechips.rocketchip.system.DefaultRV32Config.fir@199722.4]
  assign _GEN_545 = _T_939 ? _GEN_445 : sectored_entries_7_valid_3; // @[TLB.scala 217:42:freechips.rocketchip.system.DefaultRV32Config.fir@199722.4]
  assign _T_1659 = {OptimizationBarrier_19_io_y_ae,OptimizationBarrier_18_io_y_ae,OptimizationBarrier_17_io_y_ae,OptimizationBarrier_16_io_y_ae,OptimizationBarrier_15_io_y_ae,OptimizationBarrier_14_io_y_ae}; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@201191.4]
  assign ptw_ae_array = {1'h0,OptimizationBarrier_26_io_y_ae,OptimizationBarrier_25_io_y_ae,OptimizationBarrier_24_io_y_ae,OptimizationBarrier_23_io_y_ae,OptimizationBarrier_22_io_y_ae,OptimizationBarrier_21_io_y_ae,OptimizationBarrier_20_io_y_ae,_T_1659}; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@201199.4]
  assign _T_1673 = {OptimizationBarrier_19_io_y_u,OptimizationBarrier_18_io_y_u,OptimizationBarrier_17_io_y_u,OptimizationBarrier_16_io_y_u,OptimizationBarrier_15_io_y_u,OptimizationBarrier_14_io_y_u}; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@201206.4]
  assign _T_1680 = {OptimizationBarrier_26_io_y_u,OptimizationBarrier_25_io_y_u,OptimizationBarrier_24_io_y_u,OptimizationBarrier_23_io_y_u,OptimizationBarrier_22_io_y_u,OptimizationBarrier_21_io_y_u,OptimizationBarrier_20_io_y_u,_T_1673}; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@201213.4]
  assign _T_1694 = ~_T_1680; // @[TLB.scala 256:98:freechips.rocketchip.system.DefaultRV32Config.fir@201227.4]
  assign priv_x_ok = priv_s ? _T_1694 : _T_1680; // @[TLB.scala 257:22:freechips.rocketchip.system.DefaultRV32Config.fir@201255.4]
  assign _T_1737 = {OptimizationBarrier_19_io_y_sx,OptimizationBarrier_18_io_y_sx,OptimizationBarrier_17_io_y_sx,OptimizationBarrier_16_io_y_sx,OptimizationBarrier_15_io_y_sx,OptimizationBarrier_14_io_y_sx}; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@201272.4]
  assign _T_1744 = {OptimizationBarrier_26_io_y_sx,OptimizationBarrier_25_io_y_sx,OptimizationBarrier_24_io_y_sx,OptimizationBarrier_23_io_y_sx,OptimizationBarrier_22_io_y_sx,OptimizationBarrier_21_io_y_sx,OptimizationBarrier_20_io_y_sx,_T_1737}; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@201279.4]
  assign _T_1773 = priv_x_ok & _T_1744; // @[TLB.scala 260:39:freechips.rocketchip.system.DefaultRV32Config.fir@201310.4]
  assign x_array = {1'h1,_T_1773}; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@201311.4]
  assign _T_1788 = ~ptw_ae_array; // @[TLB.scala 261:89:freechips.rocketchip.system.DefaultRV32Config.fir@201326.4]
  assign _T_1805 = prot_x ? 2'h3 : 2'h0; // @[Bitwise.scala 72:12:freechips.rocketchip.system.DefaultRV32Config.fir@201345.4]
  assign _T_1810 = {OptimizationBarrier_32_io_y_px,OptimizationBarrier_31_io_y_px,OptimizationBarrier_30_io_y_px,OptimizationBarrier_29_io_y_px,OptimizationBarrier_28_io_y_px,OptimizationBarrier_27_io_y_px}; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@201350.4]
  assign _T_1817 = {_T_1805,OptimizationBarrier_38_io_y_px,OptimizationBarrier_37_io_y_px,OptimizationBarrier_36_io_y_px,OptimizationBarrier_35_io_y_px,OptimizationBarrier_34_io_y_px,OptimizationBarrier_33_io_y_px,_T_1810}; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@201357.4]
  assign px_array = _T_1817 & _T_1788; // @[TLB.scala 263:87:freechips.rocketchip.system.DefaultRV32Config.fir@201359.4]
  assign _T_1833 = cacheable ? 2'h3 : 2'h0; // @[Bitwise.scala 72:12:freechips.rocketchip.system.DefaultRV32Config.fir@201375.4]
  assign _T_1838 = {OptimizationBarrier_32_io_y_c,OptimizationBarrier_31_io_y_c,OptimizationBarrier_30_io_y_c,OptimizationBarrier_29_io_y_c,OptimizationBarrier_28_io_y_c,OptimizationBarrier_27_io_y_c}; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@201380.4]
  assign c_array = {_T_1833,OptimizationBarrier_38_io_y_c,OptimizationBarrier_37_io_y_c,OptimizationBarrier_36_io_y_c,OptimizationBarrier_35_io_y_c,OptimizationBarrier_34_io_y_c,OptimizationBarrier_33_io_y_c,_T_1838}; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@201387.4]
  assign _T_2003 = x_array | ptw_ae_array; // @[TLB.scala 313:33:freechips.rocketchip.system.DefaultRV32Config.fir@201570.4]
  assign pf_inst_array = ~_T_2003; // @[TLB.scala 313:23:freechips.rocketchip.system.DefaultRV32Config.fir@201571.4]
  assign tlb_hit = |real_hits; // @[TLB.scala 315:27:freechips.rocketchip.system.DefaultRV32Config.fir@201572.4]
  assign _T_2006 = ~tlb_hit; // @[TLB.scala 316:43:freechips.rocketchip.system.DefaultRV32Config.fir@201575.4]
  assign tlb_miss = vm_enabled & _T_2006; // @[TLB.scala 316:40:freechips.rocketchip.system.DefaultRV32Config.fir@201576.4]
  assign _T_2009 = io_req_valid & vm_enabled; // @[TLB.scala 320:22:freechips.rocketchip.system.DefaultRV32Config.fir@201579.4]
  assign _T_2010 = sector_hits_0 | sector_hits_1; // @[package.scala 64:59:freechips.rocketchip.system.DefaultRV32Config.fir@201581.6]
  assign _T_2011 = _T_2010 | sector_hits_2; // @[package.scala 64:59:freechips.rocketchip.system.DefaultRV32Config.fir@201582.6]
  assign _T_2012 = _T_2011 | sector_hits_3; // @[package.scala 64:59:freechips.rocketchip.system.DefaultRV32Config.fir@201583.6]
  assign _T_2013 = _T_2012 | sector_hits_4; // @[package.scala 64:59:freechips.rocketchip.system.DefaultRV32Config.fir@201584.6]
  assign _T_2014 = _T_2013 | sector_hits_5; // @[package.scala 64:59:freechips.rocketchip.system.DefaultRV32Config.fir@201585.6]
  assign _T_2015 = _T_2014 | sector_hits_6; // @[package.scala 64:59:freechips.rocketchip.system.DefaultRV32Config.fir@201586.6]
  assign _T_2016 = _T_2015 | sector_hits_7; // @[package.scala 64:59:freechips.rocketchip.system.DefaultRV32Config.fir@201587.6]
  assign _T_2023 = {sector_hits_7,sector_hits_6,sector_hits_5,sector_hits_4,sector_hits_3,sector_hits_2,sector_hits_1,sector_hits_0}; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@201595.8]
  assign _T_2026 = |_T_2023[7:4]; // @[OneHot.scala 32:14:freechips.rocketchip.system.DefaultRV32Config.fir@201598.8]
  assign _T_2027 = _T_2023[7:4] | _T_2023[3:0]; // @[OneHot.scala 32:28:freechips.rocketchip.system.DefaultRV32Config.fir@201599.8]
  assign _T_2030 = |_T_2027[3:2]; // @[OneHot.scala 32:14:freechips.rocketchip.system.DefaultRV32Config.fir@201602.8]
  assign _T_2031 = _T_2027[3:2] | _T_2027[1:0]; // @[OneHot.scala 32:28:freechips.rocketchip.system.DefaultRV32Config.fir@201603.8]
  assign _T_2034 = {_T_2026,_T_2030,_T_2031[1]}; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@201606.8]
  assign _T_2037 = ~_T_2034[2]; // @[Replacement.scala 186:33:freechips.rocketchip.system.DefaultRV32Config.fir@201609.8]
  assign _T_2042 = ~_T_2034[1]; // @[Replacement.scala 186:33:freechips.rocketchip.system.DefaultRV32Config.fir@201614.8]
  assign _T_2047 = ~_T_2034[0]; // @[Replacement.scala 208:7:freechips.rocketchip.system.DefaultRV32Config.fir@201619.8]
  assign _T_2048 = _T_2042 ? _T_2007[4] : _T_2047; // @[Replacement.scala 193:16:freechips.rocketchip.system.DefaultRV32Config.fir@201620.8]
  assign _T_2052 = _T_2042 ? _T_2047 : _T_2007[3]; // @[Replacement.scala 196:16:freechips.rocketchip.system.DefaultRV32Config.fir@201624.8]
  assign _T_2054 = {_T_2042,_T_2048,_T_2052}; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@201626.8]
  assign _T_2055 = _T_2037 ? _T_2007[5:3] : _T_2054; // @[Replacement.scala 193:16:freechips.rocketchip.system.DefaultRV32Config.fir@201627.8]
  assign _T_2064 = _T_2042 ? _T_2007[1] : _T_2047; // @[Replacement.scala 193:16:freechips.rocketchip.system.DefaultRV32Config.fir@201636.8]
  assign _T_2068 = _T_2042 ? _T_2047 : _T_2007[0]; // @[Replacement.scala 196:16:freechips.rocketchip.system.DefaultRV32Config.fir@201640.8]
  assign _T_2070 = {_T_2042,_T_2064,_T_2068}; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@201642.8]
  assign _T_2071 = _T_2037 ? _T_2070 : _T_2007[2:0]; // @[Replacement.scala 196:16:freechips.rocketchip.system.DefaultRV32Config.fir@201643.8]
  assign _T_2073 = {_T_2037,_T_2055,_T_2071}; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@201645.8]
  assign _T_2074 = superpage_hits_0 | superpage_hits_1; // @[package.scala 64:59:freechips.rocketchip.system.DefaultRV32Config.fir@201648.6]
  assign _T_2075 = _T_2074 | superpage_hits_2; // @[package.scala 64:59:freechips.rocketchip.system.DefaultRV32Config.fir@201649.6]
  assign _T_2076 = _T_2075 | superpage_hits_3; // @[package.scala 64:59:freechips.rocketchip.system.DefaultRV32Config.fir@201650.6]
  assign _T_2079 = {superpage_hits_3,superpage_hits_2,superpage_hits_1,superpage_hits_0}; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@201654.8]
  assign _T_2082 = |_T_2079[3:2]; // @[OneHot.scala 32:14:freechips.rocketchip.system.DefaultRV32Config.fir@201657.8]
  assign _T_2083 = _T_2079[3:2] | _T_2079[1:0]; // @[OneHot.scala 32:28:freechips.rocketchip.system.DefaultRV32Config.fir@201658.8]
  assign _T_2085 = {_T_2082,_T_2083[1]}; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@201660.8]
  assign _T_2088 = ~_T_2085[1]; // @[Replacement.scala 186:33:freechips.rocketchip.system.DefaultRV32Config.fir@201663.8]
  assign _T_2093 = ~_T_2085[0]; // @[Replacement.scala 208:7:freechips.rocketchip.system.DefaultRV32Config.fir@201668.8]
  assign _T_2094 = _T_2088 ? _T_2008[1] : _T_2093; // @[Replacement.scala 193:16:freechips.rocketchip.system.DefaultRV32Config.fir@201669.8]
  assign _T_2098 = _T_2088 ? _T_2093 : _T_2008[0]; // @[Replacement.scala 196:16:freechips.rocketchip.system.DefaultRV32Config.fir@201673.8]
  assign _T_2100 = {_T_2088,_T_2094,_T_2098}; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@201675.8]
  assign _T_2110 = real_hits[1] | real_hits[2]; // @[Misc.scala 182:16:freechips.rocketchip.system.DefaultRV32Config.fir@201688.4]
  assign _T_2112 = real_hits[1] & real_hits[2]; // @[Misc.scala 182:61:freechips.rocketchip.system.DefaultRV32Config.fir@201690.4]
  assign _T_2114 = real_hits[0] | _T_2110; // @[Misc.scala 182:16:freechips.rocketchip.system.DefaultRV32Config.fir@201692.4]
  assign _T_2116 = real_hits[0] & _T_2110; // @[Misc.scala 182:61:freechips.rocketchip.system.DefaultRV32Config.fir@201694.4]
  assign _T_2117 = _T_2112 | _T_2116; // @[Misc.scala 182:49:freechips.rocketchip.system.DefaultRV32Config.fir@201695.4]
  assign _T_2126 = real_hits[4] | real_hits[5]; // @[Misc.scala 182:16:freechips.rocketchip.system.DefaultRV32Config.fir@201704.4]
  assign _T_2128 = real_hits[4] & real_hits[5]; // @[Misc.scala 182:61:freechips.rocketchip.system.DefaultRV32Config.fir@201706.4]
  assign _T_2130 = real_hits[3] | _T_2126; // @[Misc.scala 182:16:freechips.rocketchip.system.DefaultRV32Config.fir@201708.4]
  assign _T_2132 = real_hits[3] & _T_2126; // @[Misc.scala 182:61:freechips.rocketchip.system.DefaultRV32Config.fir@201710.4]
  assign _T_2133 = _T_2128 | _T_2132; // @[Misc.scala 182:49:freechips.rocketchip.system.DefaultRV32Config.fir@201711.4]
  assign _T_2134 = _T_2114 | _T_2130; // @[Misc.scala 182:16:freechips.rocketchip.system.DefaultRV32Config.fir@201712.4]
  assign _T_2135 = _T_2117 | _T_2133; // @[Misc.scala 182:37:freechips.rocketchip.system.DefaultRV32Config.fir@201713.4]
  assign _T_2136 = _T_2114 & _T_2130; // @[Misc.scala 182:61:freechips.rocketchip.system.DefaultRV32Config.fir@201714.4]
  assign _T_2137 = _T_2135 | _T_2136; // @[Misc.scala 182:49:freechips.rocketchip.system.DefaultRV32Config.fir@201715.4]
  assign _T_2147 = real_hits[7] | real_hits[8]; // @[Misc.scala 182:16:freechips.rocketchip.system.DefaultRV32Config.fir@201725.4]
  assign _T_2149 = real_hits[7] & real_hits[8]; // @[Misc.scala 182:61:freechips.rocketchip.system.DefaultRV32Config.fir@201727.4]
  assign _T_2151 = real_hits[6] | _T_2147; // @[Misc.scala 182:16:freechips.rocketchip.system.DefaultRV32Config.fir@201729.4]
  assign _T_2153 = real_hits[6] & _T_2147; // @[Misc.scala 182:61:freechips.rocketchip.system.DefaultRV32Config.fir@201731.4]
  assign _T_2154 = _T_2149 | _T_2153; // @[Misc.scala 182:49:freechips.rocketchip.system.DefaultRV32Config.fir@201732.4]
  assign _T_2161 = real_hits[9] | real_hits[10]; // @[Misc.scala 182:16:freechips.rocketchip.system.DefaultRV32Config.fir@201739.4]
  assign _T_2163 = real_hits[9] & real_hits[10]; // @[Misc.scala 182:61:freechips.rocketchip.system.DefaultRV32Config.fir@201741.4]
  assign _T_2170 = real_hits[11] | real_hits[12]; // @[Misc.scala 182:16:freechips.rocketchip.system.DefaultRV32Config.fir@201748.4]
  assign _T_2172 = real_hits[11] & real_hits[12]; // @[Misc.scala 182:61:freechips.rocketchip.system.DefaultRV32Config.fir@201750.4]
  assign _T_2174 = _T_2161 | _T_2170; // @[Misc.scala 182:16:freechips.rocketchip.system.DefaultRV32Config.fir@201752.4]
  assign _T_2175 = _T_2163 | _T_2172; // @[Misc.scala 182:37:freechips.rocketchip.system.DefaultRV32Config.fir@201753.4]
  assign _T_2176 = _T_2161 & _T_2170; // @[Misc.scala 182:61:freechips.rocketchip.system.DefaultRV32Config.fir@201754.4]
  assign _T_2177 = _T_2175 | _T_2176; // @[Misc.scala 182:49:freechips.rocketchip.system.DefaultRV32Config.fir@201755.4]
  assign _T_2178 = _T_2151 | _T_2174; // @[Misc.scala 182:16:freechips.rocketchip.system.DefaultRV32Config.fir@201756.4]
  assign _T_2179 = _T_2154 | _T_2177; // @[Misc.scala 182:37:freechips.rocketchip.system.DefaultRV32Config.fir@201757.4]
  assign _T_2180 = _T_2151 & _T_2174; // @[Misc.scala 182:61:freechips.rocketchip.system.DefaultRV32Config.fir@201758.4]
  assign _T_2181 = _T_2179 | _T_2180; // @[Misc.scala 182:49:freechips.rocketchip.system.DefaultRV32Config.fir@201759.4]
  assign _T_2183 = _T_2137 | _T_2181; // @[Misc.scala 182:37:freechips.rocketchip.system.DefaultRV32Config.fir@201761.4]
  assign _T_2184 = _T_2134 & _T_2178; // @[Misc.scala 182:61:freechips.rocketchip.system.DefaultRV32Config.fir@201762.4]
  assign multipleHits = _T_2183 | _T_2184; // @[Misc.scala 182:49:freechips.rocketchip.system.DefaultRV32Config.fir@201763.4]
  assign _T_2194 = pf_inst_array & hits; // @[TLB.scala 335:47:freechips.rocketchip.system.DefaultRV32Config.fir@201776.4]
  assign _T_2201 = ~px_array; // @[TLB.scala 338:23:freechips.rocketchip.system.DefaultRV32Config.fir@201786.4]
  assign _T_2202 = _T_2201 & hits; // @[TLB.scala 338:33:freechips.rocketchip.system.DefaultRV32Config.fir@201787.4]
  assign _T_2208 = c_array & hits; // @[TLB.scala 342:33:freechips.rocketchip.system.DefaultRV32Config.fir@201797.4]
  assign _T_2215 = io_ptw_resp_valid | tlb_miss; // @[TLB.scala 345:29:freechips.rocketchip.system.DefaultRV32Config.fir@201807.4]
  assign _T_2221 = io_req_ready & io_req_valid; // @[Decoupled.scala 40:37:freechips.rocketchip.system.DefaultRV32Config.fir@201818.4]
  assign _T_2222 = _T_2221 & tlb_miss; // @[TLB.scala 354:25:freechips.rocketchip.system.DefaultRV32Config.fir@201819.4]
  assign _T_2228 = _T_2008[2] ? _T_2008[1] : _T_2008[0]; // @[Replacement.scala 240:16:freechips.rocketchip.system.DefaultRV32Config.fir@201828.6]
  assign _T_2229 = {_T_2008[2],_T_2228}; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@201829.6]
  assign _T_2232 = {superpage_entries_3_valid_0,superpage_entries_2_valid_0,superpage_entries_1_valid_0,superpage_entries_0_valid_0}; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@201832.6]
  assign _T_2233 = &_T_2232; // @[TLB.scala 402:16:freechips.rocketchip.system.DefaultRV32Config.fir@201833.6]
  assign _T_2234 = ~_T_2232; // @[TLB.scala 402:43:freechips.rocketchip.system.DefaultRV32Config.fir@201834.6]
  assign _T_2251 = _T_2007[5] ? _T_2007[4] : _T_2007[3]; // @[Replacement.scala 240:16:freechips.rocketchip.system.DefaultRV32Config.fir@201852.6]
  assign _T_2252 = {_T_2007[5],_T_2251}; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@201853.6]
  assign _T_2258 = _T_2007[2] ? _T_2007[1] : _T_2007[0]; // @[Replacement.scala 240:16:freechips.rocketchip.system.DefaultRV32Config.fir@201859.6]
  assign _T_2259 = {_T_2007[2],_T_2258}; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@201860.6]
  assign _T_2260 = _T_2007[6] ? _T_2252 : _T_2259; // @[Replacement.scala 240:16:freechips.rocketchip.system.DefaultRV32Config.fir@201861.6]
  assign _T_2261 = {_T_2007[6],_T_2260}; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@201862.6]
  assign _T_2292 = {_T_454,_T_448,_T_442,_T_436,_T_430,_T_424,_T_418,_T_412}; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@201893.6]
  assign _T_2293 = &_T_2292; // @[TLB.scala 402:16:freechips.rocketchip.system.DefaultRV32Config.fir@201894.6]
  assign _T_2294 = ~_T_2292; // @[TLB.scala 402:43:freechips.rocketchip.system.DefaultRV32Config.fir@201895.6]
  assign _T_2338 = state == 2'h2; // @[TLB.scala 368:17:freechips.rocketchip.system.DefaultRV32Config.fir@201954.4]
  assign _T_2339 = _T_2338 & io_sfence_valid; // @[TLB.scala 368:28:freechips.rocketchip.system.DefaultRV32Config.fir@201955.4]
  assign _T_2340 = ~io_sfence_bits_rs1; // @[TLB.scala 376:14:freechips.rocketchip.system.DefaultRV32Config.fir@201963.6]
  assign _T_2342 = io_sfence_bits_addr[31:12] == vpn; // @[TLB.scala 376:72:freechips.rocketchip.system.DefaultRV32Config.fir@201965.6]
  assign _T_2343 = _T_2340 | _T_2342; // @[TLB.scala 376:34:freechips.rocketchip.system.DefaultRV32Config.fir@201966.6]
  assign _T_2345 = _T_2343 | reset; // @[TLB.scala 376:13:freechips.rocketchip.system.DefaultRV32Config.fir@201968.6]
  assign _T_2346 = ~_T_2345; // @[TLB.scala 376:13:freechips.rocketchip.system.DefaultRV32Config.fir@201969.6]
  assign _T_2353 = _T_413[19:10] == 10'h0; // @[TLB.scala 135:61:freechips.rocketchip.system.DefaultRV32Config.fir@201984.8]
  assign _T_2498 = ~sectored_entries_0_data_0[13]; // @[TLB.scala 143:13:freechips.rocketchip.system.DefaultRV32Config.fir@202298.10]
  assign _GEN_648 = _T_2498 ? 1'h0 : _GEN_472; // @[TLB.scala 143:19:freechips.rocketchip.system.DefaultRV32Config.fir@202299.10]
  assign _T_2499 = ~sectored_entries_0_data_1[13]; // @[TLB.scala 143:13:freechips.rocketchip.system.DefaultRV32Config.fir@202302.10]
  assign _GEN_649 = _T_2499 ? 1'h0 : _GEN_473; // @[TLB.scala 143:19:freechips.rocketchip.system.DefaultRV32Config.fir@202303.10]
  assign _T_2500 = ~sectored_entries_0_data_2[13]; // @[TLB.scala 143:13:freechips.rocketchip.system.DefaultRV32Config.fir@202306.10]
  assign _GEN_650 = _T_2500 ? 1'h0 : _GEN_474; // @[TLB.scala 143:19:freechips.rocketchip.system.DefaultRV32Config.fir@202307.10]
  assign _T_2501 = ~sectored_entries_0_data_3[13]; // @[TLB.scala 143:13:freechips.rocketchip.system.DefaultRV32Config.fir@202310.10]
  assign _GEN_651 = _T_2501 ? 1'h0 : _GEN_475; // @[TLB.scala 143:19:freechips.rocketchip.system.DefaultRV32Config.fir@202311.10]
  assign _GEN_652 = io_sfence_bits_rs2 & _GEN_648; // @[TLB.scala 379:40:freechips.rocketchip.system.DefaultRV32Config.fir@202149.8]
  assign _GEN_653 = io_sfence_bits_rs2 & _GEN_649; // @[TLB.scala 379:40:freechips.rocketchip.system.DefaultRV32Config.fir@202149.8]
  assign _GEN_654 = io_sfence_bits_rs2 & _GEN_650; // @[TLB.scala 379:40:freechips.rocketchip.system.DefaultRV32Config.fir@202149.8]
  assign _GEN_655 = io_sfence_bits_rs2 & _GEN_651; // @[TLB.scala 379:40:freechips.rocketchip.system.DefaultRV32Config.fir@202149.8]
  assign _T_2508 = _T_419[19:10] == 10'h0; // @[TLB.scala 135:61:freechips.rocketchip.system.DefaultRV32Config.fir@202331.8]
  assign _T_2653 = ~sectored_entries_1_data_0[13]; // @[TLB.scala 143:13:freechips.rocketchip.system.DefaultRV32Config.fir@202645.10]
  assign _GEN_676 = _T_2653 ? 1'h0 : _GEN_482; // @[TLB.scala 143:19:freechips.rocketchip.system.DefaultRV32Config.fir@202646.10]
  assign _T_2654 = ~sectored_entries_1_data_1[13]; // @[TLB.scala 143:13:freechips.rocketchip.system.DefaultRV32Config.fir@202649.10]
  assign _GEN_677 = _T_2654 ? 1'h0 : _GEN_483; // @[TLB.scala 143:19:freechips.rocketchip.system.DefaultRV32Config.fir@202650.10]
  assign _T_2655 = ~sectored_entries_1_data_2[13]; // @[TLB.scala 143:13:freechips.rocketchip.system.DefaultRV32Config.fir@202653.10]
  assign _GEN_678 = _T_2655 ? 1'h0 : _GEN_484; // @[TLB.scala 143:19:freechips.rocketchip.system.DefaultRV32Config.fir@202654.10]
  assign _T_2656 = ~sectored_entries_1_data_3[13]; // @[TLB.scala 143:13:freechips.rocketchip.system.DefaultRV32Config.fir@202657.10]
  assign _GEN_679 = _T_2656 ? 1'h0 : _GEN_485; // @[TLB.scala 143:19:freechips.rocketchip.system.DefaultRV32Config.fir@202658.10]
  assign _GEN_680 = io_sfence_bits_rs2 & _GEN_676; // @[TLB.scala 379:40:freechips.rocketchip.system.DefaultRV32Config.fir@202496.8]
  assign _GEN_681 = io_sfence_bits_rs2 & _GEN_677; // @[TLB.scala 379:40:freechips.rocketchip.system.DefaultRV32Config.fir@202496.8]
  assign _GEN_682 = io_sfence_bits_rs2 & _GEN_678; // @[TLB.scala 379:40:freechips.rocketchip.system.DefaultRV32Config.fir@202496.8]
  assign _GEN_683 = io_sfence_bits_rs2 & _GEN_679; // @[TLB.scala 379:40:freechips.rocketchip.system.DefaultRV32Config.fir@202496.8]
  assign _T_2663 = _T_425[19:10] == 10'h0; // @[TLB.scala 135:61:freechips.rocketchip.system.DefaultRV32Config.fir@202678.8]
  assign _T_2808 = ~sectored_entries_2_data_0[13]; // @[TLB.scala 143:13:freechips.rocketchip.system.DefaultRV32Config.fir@202992.10]
  assign _GEN_704 = _T_2808 ? 1'h0 : _GEN_492; // @[TLB.scala 143:19:freechips.rocketchip.system.DefaultRV32Config.fir@202993.10]
  assign _T_2809 = ~sectored_entries_2_data_1[13]; // @[TLB.scala 143:13:freechips.rocketchip.system.DefaultRV32Config.fir@202996.10]
  assign _GEN_705 = _T_2809 ? 1'h0 : _GEN_493; // @[TLB.scala 143:19:freechips.rocketchip.system.DefaultRV32Config.fir@202997.10]
  assign _T_2810 = ~sectored_entries_2_data_2[13]; // @[TLB.scala 143:13:freechips.rocketchip.system.DefaultRV32Config.fir@203000.10]
  assign _GEN_706 = _T_2810 ? 1'h0 : _GEN_494; // @[TLB.scala 143:19:freechips.rocketchip.system.DefaultRV32Config.fir@203001.10]
  assign _T_2811 = ~sectored_entries_2_data_3[13]; // @[TLB.scala 143:13:freechips.rocketchip.system.DefaultRV32Config.fir@203004.10]
  assign _GEN_707 = _T_2811 ? 1'h0 : _GEN_495; // @[TLB.scala 143:19:freechips.rocketchip.system.DefaultRV32Config.fir@203005.10]
  assign _GEN_708 = io_sfence_bits_rs2 & _GEN_704; // @[TLB.scala 379:40:freechips.rocketchip.system.DefaultRV32Config.fir@202843.8]
  assign _GEN_709 = io_sfence_bits_rs2 & _GEN_705; // @[TLB.scala 379:40:freechips.rocketchip.system.DefaultRV32Config.fir@202843.8]
  assign _GEN_710 = io_sfence_bits_rs2 & _GEN_706; // @[TLB.scala 379:40:freechips.rocketchip.system.DefaultRV32Config.fir@202843.8]
  assign _GEN_711 = io_sfence_bits_rs2 & _GEN_707; // @[TLB.scala 379:40:freechips.rocketchip.system.DefaultRV32Config.fir@202843.8]
  assign _T_2818 = _T_431[19:10] == 10'h0; // @[TLB.scala 135:61:freechips.rocketchip.system.DefaultRV32Config.fir@203025.8]
  assign _T_2963 = ~sectored_entries_3_data_0[13]; // @[TLB.scala 143:13:freechips.rocketchip.system.DefaultRV32Config.fir@203339.10]
  assign _GEN_732 = _T_2963 ? 1'h0 : _GEN_502; // @[TLB.scala 143:19:freechips.rocketchip.system.DefaultRV32Config.fir@203340.10]
  assign _T_2964 = ~sectored_entries_3_data_1[13]; // @[TLB.scala 143:13:freechips.rocketchip.system.DefaultRV32Config.fir@203343.10]
  assign _GEN_733 = _T_2964 ? 1'h0 : _GEN_503; // @[TLB.scala 143:19:freechips.rocketchip.system.DefaultRV32Config.fir@203344.10]
  assign _T_2965 = ~sectored_entries_3_data_2[13]; // @[TLB.scala 143:13:freechips.rocketchip.system.DefaultRV32Config.fir@203347.10]
  assign _GEN_734 = _T_2965 ? 1'h0 : _GEN_504; // @[TLB.scala 143:19:freechips.rocketchip.system.DefaultRV32Config.fir@203348.10]
  assign _T_2966 = ~sectored_entries_3_data_3[13]; // @[TLB.scala 143:13:freechips.rocketchip.system.DefaultRV32Config.fir@203351.10]
  assign _GEN_735 = _T_2966 ? 1'h0 : _GEN_505; // @[TLB.scala 143:19:freechips.rocketchip.system.DefaultRV32Config.fir@203352.10]
  assign _GEN_736 = io_sfence_bits_rs2 & _GEN_732; // @[TLB.scala 379:40:freechips.rocketchip.system.DefaultRV32Config.fir@203190.8]
  assign _GEN_737 = io_sfence_bits_rs2 & _GEN_733; // @[TLB.scala 379:40:freechips.rocketchip.system.DefaultRV32Config.fir@203190.8]
  assign _GEN_738 = io_sfence_bits_rs2 & _GEN_734; // @[TLB.scala 379:40:freechips.rocketchip.system.DefaultRV32Config.fir@203190.8]
  assign _GEN_739 = io_sfence_bits_rs2 & _GEN_735; // @[TLB.scala 379:40:freechips.rocketchip.system.DefaultRV32Config.fir@203190.8]
  assign _T_2973 = _T_437[19:10] == 10'h0; // @[TLB.scala 135:61:freechips.rocketchip.system.DefaultRV32Config.fir@203372.8]
  assign _T_3118 = ~sectored_entries_4_data_0[13]; // @[TLB.scala 143:13:freechips.rocketchip.system.DefaultRV32Config.fir@203686.10]
  assign _GEN_760 = _T_3118 ? 1'h0 : _GEN_512; // @[TLB.scala 143:19:freechips.rocketchip.system.DefaultRV32Config.fir@203687.10]
  assign _T_3119 = ~sectored_entries_4_data_1[13]; // @[TLB.scala 143:13:freechips.rocketchip.system.DefaultRV32Config.fir@203690.10]
  assign _GEN_761 = _T_3119 ? 1'h0 : _GEN_513; // @[TLB.scala 143:19:freechips.rocketchip.system.DefaultRV32Config.fir@203691.10]
  assign _T_3120 = ~sectored_entries_4_data_2[13]; // @[TLB.scala 143:13:freechips.rocketchip.system.DefaultRV32Config.fir@203694.10]
  assign _GEN_762 = _T_3120 ? 1'h0 : _GEN_514; // @[TLB.scala 143:19:freechips.rocketchip.system.DefaultRV32Config.fir@203695.10]
  assign _T_3121 = ~sectored_entries_4_data_3[13]; // @[TLB.scala 143:13:freechips.rocketchip.system.DefaultRV32Config.fir@203698.10]
  assign _GEN_763 = _T_3121 ? 1'h0 : _GEN_515; // @[TLB.scala 143:19:freechips.rocketchip.system.DefaultRV32Config.fir@203699.10]
  assign _GEN_764 = io_sfence_bits_rs2 & _GEN_760; // @[TLB.scala 379:40:freechips.rocketchip.system.DefaultRV32Config.fir@203537.8]
  assign _GEN_765 = io_sfence_bits_rs2 & _GEN_761; // @[TLB.scala 379:40:freechips.rocketchip.system.DefaultRV32Config.fir@203537.8]
  assign _GEN_766 = io_sfence_bits_rs2 & _GEN_762; // @[TLB.scala 379:40:freechips.rocketchip.system.DefaultRV32Config.fir@203537.8]
  assign _GEN_767 = io_sfence_bits_rs2 & _GEN_763; // @[TLB.scala 379:40:freechips.rocketchip.system.DefaultRV32Config.fir@203537.8]
  assign _T_3128 = _T_443[19:10] == 10'h0; // @[TLB.scala 135:61:freechips.rocketchip.system.DefaultRV32Config.fir@203719.8]
  assign _T_3273 = ~sectored_entries_5_data_0[13]; // @[TLB.scala 143:13:freechips.rocketchip.system.DefaultRV32Config.fir@204033.10]
  assign _GEN_788 = _T_3273 ? 1'h0 : _GEN_522; // @[TLB.scala 143:19:freechips.rocketchip.system.DefaultRV32Config.fir@204034.10]
  assign _T_3274 = ~sectored_entries_5_data_1[13]; // @[TLB.scala 143:13:freechips.rocketchip.system.DefaultRV32Config.fir@204037.10]
  assign _GEN_789 = _T_3274 ? 1'h0 : _GEN_523; // @[TLB.scala 143:19:freechips.rocketchip.system.DefaultRV32Config.fir@204038.10]
  assign _T_3275 = ~sectored_entries_5_data_2[13]; // @[TLB.scala 143:13:freechips.rocketchip.system.DefaultRV32Config.fir@204041.10]
  assign _GEN_790 = _T_3275 ? 1'h0 : _GEN_524; // @[TLB.scala 143:19:freechips.rocketchip.system.DefaultRV32Config.fir@204042.10]
  assign _T_3276 = ~sectored_entries_5_data_3[13]; // @[TLB.scala 143:13:freechips.rocketchip.system.DefaultRV32Config.fir@204045.10]
  assign _GEN_791 = _T_3276 ? 1'h0 : _GEN_525; // @[TLB.scala 143:19:freechips.rocketchip.system.DefaultRV32Config.fir@204046.10]
  assign _GEN_792 = io_sfence_bits_rs2 & _GEN_788; // @[TLB.scala 379:40:freechips.rocketchip.system.DefaultRV32Config.fir@203884.8]
  assign _GEN_793 = io_sfence_bits_rs2 & _GEN_789; // @[TLB.scala 379:40:freechips.rocketchip.system.DefaultRV32Config.fir@203884.8]
  assign _GEN_794 = io_sfence_bits_rs2 & _GEN_790; // @[TLB.scala 379:40:freechips.rocketchip.system.DefaultRV32Config.fir@203884.8]
  assign _GEN_795 = io_sfence_bits_rs2 & _GEN_791; // @[TLB.scala 379:40:freechips.rocketchip.system.DefaultRV32Config.fir@203884.8]
  assign _T_3283 = _T_449[19:10] == 10'h0; // @[TLB.scala 135:61:freechips.rocketchip.system.DefaultRV32Config.fir@204066.8]
  assign _T_3428 = ~sectored_entries_6_data_0[13]; // @[TLB.scala 143:13:freechips.rocketchip.system.DefaultRV32Config.fir@204380.10]
  assign _GEN_816 = _T_3428 ? 1'h0 : _GEN_532; // @[TLB.scala 143:19:freechips.rocketchip.system.DefaultRV32Config.fir@204381.10]
  assign _T_3429 = ~sectored_entries_6_data_1[13]; // @[TLB.scala 143:13:freechips.rocketchip.system.DefaultRV32Config.fir@204384.10]
  assign _GEN_817 = _T_3429 ? 1'h0 : _GEN_533; // @[TLB.scala 143:19:freechips.rocketchip.system.DefaultRV32Config.fir@204385.10]
  assign _T_3430 = ~sectored_entries_6_data_2[13]; // @[TLB.scala 143:13:freechips.rocketchip.system.DefaultRV32Config.fir@204388.10]
  assign _GEN_818 = _T_3430 ? 1'h0 : _GEN_534; // @[TLB.scala 143:19:freechips.rocketchip.system.DefaultRV32Config.fir@204389.10]
  assign _T_3431 = ~sectored_entries_6_data_3[13]; // @[TLB.scala 143:13:freechips.rocketchip.system.DefaultRV32Config.fir@204392.10]
  assign _GEN_819 = _T_3431 ? 1'h0 : _GEN_535; // @[TLB.scala 143:19:freechips.rocketchip.system.DefaultRV32Config.fir@204393.10]
  assign _GEN_820 = io_sfence_bits_rs2 & _GEN_816; // @[TLB.scala 379:40:freechips.rocketchip.system.DefaultRV32Config.fir@204231.8]
  assign _GEN_821 = io_sfence_bits_rs2 & _GEN_817; // @[TLB.scala 379:40:freechips.rocketchip.system.DefaultRV32Config.fir@204231.8]
  assign _GEN_822 = io_sfence_bits_rs2 & _GEN_818; // @[TLB.scala 379:40:freechips.rocketchip.system.DefaultRV32Config.fir@204231.8]
  assign _GEN_823 = io_sfence_bits_rs2 & _GEN_819; // @[TLB.scala 379:40:freechips.rocketchip.system.DefaultRV32Config.fir@204231.8]
  assign _T_3438 = _T_455[19:10] == 10'h0; // @[TLB.scala 135:61:freechips.rocketchip.system.DefaultRV32Config.fir@204413.8]
  assign _T_3583 = ~sectored_entries_7_data_0[13]; // @[TLB.scala 143:13:freechips.rocketchip.system.DefaultRV32Config.fir@204727.10]
  assign _GEN_844 = _T_3583 ? 1'h0 : _GEN_542; // @[TLB.scala 143:19:freechips.rocketchip.system.DefaultRV32Config.fir@204728.10]
  assign _T_3584 = ~sectored_entries_7_data_1[13]; // @[TLB.scala 143:13:freechips.rocketchip.system.DefaultRV32Config.fir@204731.10]
  assign _GEN_845 = _T_3584 ? 1'h0 : _GEN_543; // @[TLB.scala 143:19:freechips.rocketchip.system.DefaultRV32Config.fir@204732.10]
  assign _T_3585 = ~sectored_entries_7_data_2[13]; // @[TLB.scala 143:13:freechips.rocketchip.system.DefaultRV32Config.fir@204735.10]
  assign _GEN_846 = _T_3585 ? 1'h0 : _GEN_544; // @[TLB.scala 143:19:freechips.rocketchip.system.DefaultRV32Config.fir@204736.10]
  assign _T_3586 = ~sectored_entries_7_data_3[13]; // @[TLB.scala 143:13:freechips.rocketchip.system.DefaultRV32Config.fir@204739.10]
  assign _GEN_847 = _T_3586 ? 1'h0 : _GEN_545; // @[TLB.scala 143:19:freechips.rocketchip.system.DefaultRV32Config.fir@204740.10]
  assign _GEN_848 = io_sfence_bits_rs2 & _GEN_844; // @[TLB.scala 379:40:freechips.rocketchip.system.DefaultRV32Config.fir@204578.8]
  assign _GEN_849 = io_sfence_bits_rs2 & _GEN_845; // @[TLB.scala 379:40:freechips.rocketchip.system.DefaultRV32Config.fir@204578.8]
  assign _GEN_850 = io_sfence_bits_rs2 & _GEN_846; // @[TLB.scala 379:40:freechips.rocketchip.system.DefaultRV32Config.fir@204578.8]
  assign _GEN_851 = io_sfence_bits_rs2 & _GEN_847; // @[TLB.scala 379:40:freechips.rocketchip.system.DefaultRV32Config.fir@204578.8]
  assign _T_3619 = ~superpage_entries_0_data_0[13]; // @[TLB.scala 143:13:freechips.rocketchip.system.DefaultRV32Config.fir@204808.10]
  assign _GEN_857 = _T_3619 ? 1'h0 : _GEN_458; // @[TLB.scala 143:19:freechips.rocketchip.system.DefaultRV32Config.fir@204809.10]
  assign _GEN_858 = io_sfence_bits_rs2 & _GEN_857; // @[TLB.scala 379:40:freechips.rocketchip.system.DefaultRV32Config.fir@204770.8]
  assign _T_3652 = ~superpage_entries_1_data_0[13]; // @[TLB.scala 143:13:freechips.rocketchip.system.DefaultRV32Config.fir@204874.10]
  assign _GEN_861 = _T_3652 ? 1'h0 : _GEN_462; // @[TLB.scala 143:19:freechips.rocketchip.system.DefaultRV32Config.fir@204875.10]
  assign _GEN_862 = io_sfence_bits_rs2 & _GEN_861; // @[TLB.scala 379:40:freechips.rocketchip.system.DefaultRV32Config.fir@204836.8]
  assign _T_3685 = ~superpage_entries_2_data_0[13]; // @[TLB.scala 143:13:freechips.rocketchip.system.DefaultRV32Config.fir@204940.10]
  assign _GEN_865 = _T_3685 ? 1'h0 : _GEN_466; // @[TLB.scala 143:19:freechips.rocketchip.system.DefaultRV32Config.fir@204941.10]
  assign _GEN_866 = io_sfence_bits_rs2 & _GEN_865; // @[TLB.scala 379:40:freechips.rocketchip.system.DefaultRV32Config.fir@204902.8]
  assign _T_3718 = ~superpage_entries_3_data_0[13]; // @[TLB.scala 143:13:freechips.rocketchip.system.DefaultRV32Config.fir@205006.10]
  assign _GEN_869 = _T_3718 ? 1'h0 : _GEN_470; // @[TLB.scala 143:19:freechips.rocketchip.system.DefaultRV32Config.fir@205007.10]
  assign _GEN_870 = io_sfence_bits_rs2 & _GEN_869; // @[TLB.scala 379:40:freechips.rocketchip.system.DefaultRV32Config.fir@204968.8]
  assign _T_3751 = ~special_entry_data_0[13]; // @[TLB.scala 143:13:freechips.rocketchip.system.DefaultRV32Config.fir@205072.10]
  assign _GEN_873 = _T_3751 ? 1'h0 : _GEN_454; // @[TLB.scala 143:19:freechips.rocketchip.system.DefaultRV32Config.fir@205073.10]
  assign _GEN_874 = io_sfence_bits_rs2 & _GEN_873; // @[TLB.scala 379:40:freechips.rocketchip.system.DefaultRV32Config.fir@205034.8]
  assign _T_3753 = multipleHits | reset; // @[TLB.scala 383:24:freechips.rocketchip.system.DefaultRV32Config.fir@205082.4]
  assign io_req_ready = state == 2'h0; // @[TLB.scala 332:16:freechips.rocketchip.system.DefaultRV32Config.fir@201765.4]
  assign io_resp_miss = _T_2215 | multipleHits; // @[TLB.scala 345:16:freechips.rocketchip.system.DefaultRV32Config.fir@201809.4]
  assign io_resp_paddr = {ppn,io_req_bits_vaddr[11:0]}; // @[TLB.scala 346:17:freechips.rocketchip.system.DefaultRV32Config.fir@201812.4]
  assign io_resp_pf_inst = |_T_2194; // @[TLB.scala 335:19:freechips.rocketchip.system.DefaultRV32Config.fir@201779.4]
  assign io_resp_ae_inst = |_T_2202; // @[TLB.scala 338:19:freechips.rocketchip.system.DefaultRV32Config.fir@201789.4]
  assign io_resp_cacheable = |_T_2208; // @[TLB.scala 342:21:freechips.rocketchip.system.DefaultRV32Config.fir@201799.4]
  assign io_ptw_req_valid = state == 2'h1; // @[TLB.scala 348:20:freechips.rocketchip.system.DefaultRV32Config.fir@201814.4]
  assign io_ptw_req_bits_valid = ~io_kill; // @[TLB.scala 349:25:freechips.rocketchip.system.DefaultRV32Config.fir@201816.4]
  assign io_ptw_req_bits_bits_addr = r_refill_tag; // @[TLB.scala 350:29:freechips.rocketchip.system.DefaultRV32Config.fir@201817.4]
  assign OptimizationBarrier_io_x_ppn = special_entry_data_0[34:15]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@198421.4]
  assign OptimizationBarrier_io_x_u = special_entry_data_0[14]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@198421.4]
  assign OptimizationBarrier_io_x_ae = special_entry_data_0[12]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@198421.4]
  assign OptimizationBarrier_io_x_sw = special_entry_data_0[11]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@198421.4]
  assign OptimizationBarrier_io_x_sx = special_entry_data_0[10]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@198421.4]
  assign OptimizationBarrier_io_x_sr = special_entry_data_0[9]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@198421.4]
  assign OptimizationBarrier_io_x_pw = special_entry_data_0[8]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@198421.4]
  assign OptimizationBarrier_io_x_px = special_entry_data_0[7]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@198421.4]
  assign OptimizationBarrier_io_x_pr = special_entry_data_0[6]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@198421.4]
  assign OptimizationBarrier_io_x_ppp = special_entry_data_0[5]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@198421.4]
  assign OptimizationBarrier_io_x_pal = special_entry_data_0[4]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@198421.4]
  assign OptimizationBarrier_io_x_paa = special_entry_data_0[3]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@198421.4]
  assign OptimizationBarrier_io_x_eff = special_entry_data_0[2]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@198421.4]
  assign OptimizationBarrier_io_x_c = special_entry_data_0[1]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@198421.4]
  assign pmp_io_prv = mpu_priv[1:0]; // @[TLB.scala 194:14:freechips.rocketchip.system.DefaultRV32Config.fir@198452.4]
  assign pmp_io_pmp_0_cfg_l = io_ptw_pmp_0_cfg_l; // @[TLB.scala 193:14:freechips.rocketchip.system.DefaultRV32Config.fir@198444.4]
  assign pmp_io_pmp_0_cfg_a = io_ptw_pmp_0_cfg_a; // @[TLB.scala 193:14:freechips.rocketchip.system.DefaultRV32Config.fir@198444.4]
  assign pmp_io_pmp_0_cfg_x = io_ptw_pmp_0_cfg_x; // @[TLB.scala 193:14:freechips.rocketchip.system.DefaultRV32Config.fir@198444.4]
  assign pmp_io_pmp_0_cfg_w = io_ptw_pmp_0_cfg_w; // @[TLB.scala 193:14:freechips.rocketchip.system.DefaultRV32Config.fir@198444.4]
  assign pmp_io_pmp_0_cfg_r = io_ptw_pmp_0_cfg_r; // @[TLB.scala 193:14:freechips.rocketchip.system.DefaultRV32Config.fir@198444.4]
  assign pmp_io_pmp_0_addr = io_ptw_pmp_0_addr; // @[TLB.scala 193:14:freechips.rocketchip.system.DefaultRV32Config.fir@198444.4]
  assign pmp_io_pmp_0_mask = io_ptw_pmp_0_mask; // @[TLB.scala 193:14:freechips.rocketchip.system.DefaultRV32Config.fir@198444.4]
  assign pmp_io_pmp_1_cfg_l = io_ptw_pmp_1_cfg_l; // @[TLB.scala 193:14:freechips.rocketchip.system.DefaultRV32Config.fir@198445.4]
  assign pmp_io_pmp_1_cfg_a = io_ptw_pmp_1_cfg_a; // @[TLB.scala 193:14:freechips.rocketchip.system.DefaultRV32Config.fir@198445.4]
  assign pmp_io_pmp_1_cfg_x = io_ptw_pmp_1_cfg_x; // @[TLB.scala 193:14:freechips.rocketchip.system.DefaultRV32Config.fir@198445.4]
  assign pmp_io_pmp_1_cfg_w = io_ptw_pmp_1_cfg_w; // @[TLB.scala 193:14:freechips.rocketchip.system.DefaultRV32Config.fir@198445.4]
  assign pmp_io_pmp_1_cfg_r = io_ptw_pmp_1_cfg_r; // @[TLB.scala 193:14:freechips.rocketchip.system.DefaultRV32Config.fir@198445.4]
  assign pmp_io_pmp_1_addr = io_ptw_pmp_1_addr; // @[TLB.scala 193:14:freechips.rocketchip.system.DefaultRV32Config.fir@198445.4]
  assign pmp_io_pmp_1_mask = io_ptw_pmp_1_mask; // @[TLB.scala 193:14:freechips.rocketchip.system.DefaultRV32Config.fir@198445.4]
  assign pmp_io_pmp_2_cfg_l = io_ptw_pmp_2_cfg_l; // @[TLB.scala 193:14:freechips.rocketchip.system.DefaultRV32Config.fir@198446.4]
  assign pmp_io_pmp_2_cfg_a = io_ptw_pmp_2_cfg_a; // @[TLB.scala 193:14:freechips.rocketchip.system.DefaultRV32Config.fir@198446.4]
  assign pmp_io_pmp_2_cfg_x = io_ptw_pmp_2_cfg_x; // @[TLB.scala 193:14:freechips.rocketchip.system.DefaultRV32Config.fir@198446.4]
  assign pmp_io_pmp_2_cfg_w = io_ptw_pmp_2_cfg_w; // @[TLB.scala 193:14:freechips.rocketchip.system.DefaultRV32Config.fir@198446.4]
  assign pmp_io_pmp_2_cfg_r = io_ptw_pmp_2_cfg_r; // @[TLB.scala 193:14:freechips.rocketchip.system.DefaultRV32Config.fir@198446.4]
  assign pmp_io_pmp_2_addr = io_ptw_pmp_2_addr; // @[TLB.scala 193:14:freechips.rocketchip.system.DefaultRV32Config.fir@198446.4]
  assign pmp_io_pmp_2_mask = io_ptw_pmp_2_mask; // @[TLB.scala 193:14:freechips.rocketchip.system.DefaultRV32Config.fir@198446.4]
  assign pmp_io_pmp_3_cfg_l = io_ptw_pmp_3_cfg_l; // @[TLB.scala 193:14:freechips.rocketchip.system.DefaultRV32Config.fir@198447.4]
  assign pmp_io_pmp_3_cfg_a = io_ptw_pmp_3_cfg_a; // @[TLB.scala 193:14:freechips.rocketchip.system.DefaultRV32Config.fir@198447.4]
  assign pmp_io_pmp_3_cfg_x = io_ptw_pmp_3_cfg_x; // @[TLB.scala 193:14:freechips.rocketchip.system.DefaultRV32Config.fir@198447.4]
  assign pmp_io_pmp_3_cfg_w = io_ptw_pmp_3_cfg_w; // @[TLB.scala 193:14:freechips.rocketchip.system.DefaultRV32Config.fir@198447.4]
  assign pmp_io_pmp_3_cfg_r = io_ptw_pmp_3_cfg_r; // @[TLB.scala 193:14:freechips.rocketchip.system.DefaultRV32Config.fir@198447.4]
  assign pmp_io_pmp_3_addr = io_ptw_pmp_3_addr; // @[TLB.scala 193:14:freechips.rocketchip.system.DefaultRV32Config.fir@198447.4]
  assign pmp_io_pmp_3_mask = io_ptw_pmp_3_mask; // @[TLB.scala 193:14:freechips.rocketchip.system.DefaultRV32Config.fir@198447.4]
  assign pmp_io_pmp_4_cfg_l = io_ptw_pmp_4_cfg_l; // @[TLB.scala 193:14:freechips.rocketchip.system.DefaultRV32Config.fir@198448.4]
  assign pmp_io_pmp_4_cfg_a = io_ptw_pmp_4_cfg_a; // @[TLB.scala 193:14:freechips.rocketchip.system.DefaultRV32Config.fir@198448.4]
  assign pmp_io_pmp_4_cfg_x = io_ptw_pmp_4_cfg_x; // @[TLB.scala 193:14:freechips.rocketchip.system.DefaultRV32Config.fir@198448.4]
  assign pmp_io_pmp_4_cfg_w = io_ptw_pmp_4_cfg_w; // @[TLB.scala 193:14:freechips.rocketchip.system.DefaultRV32Config.fir@198448.4]
  assign pmp_io_pmp_4_cfg_r = io_ptw_pmp_4_cfg_r; // @[TLB.scala 193:14:freechips.rocketchip.system.DefaultRV32Config.fir@198448.4]
  assign pmp_io_pmp_4_addr = io_ptw_pmp_4_addr; // @[TLB.scala 193:14:freechips.rocketchip.system.DefaultRV32Config.fir@198448.4]
  assign pmp_io_pmp_4_mask = io_ptw_pmp_4_mask; // @[TLB.scala 193:14:freechips.rocketchip.system.DefaultRV32Config.fir@198448.4]
  assign pmp_io_pmp_5_cfg_l = io_ptw_pmp_5_cfg_l; // @[TLB.scala 193:14:freechips.rocketchip.system.DefaultRV32Config.fir@198449.4]
  assign pmp_io_pmp_5_cfg_a = io_ptw_pmp_5_cfg_a; // @[TLB.scala 193:14:freechips.rocketchip.system.DefaultRV32Config.fir@198449.4]
  assign pmp_io_pmp_5_cfg_x = io_ptw_pmp_5_cfg_x; // @[TLB.scala 193:14:freechips.rocketchip.system.DefaultRV32Config.fir@198449.4]
  assign pmp_io_pmp_5_cfg_w = io_ptw_pmp_5_cfg_w; // @[TLB.scala 193:14:freechips.rocketchip.system.DefaultRV32Config.fir@198449.4]
  assign pmp_io_pmp_5_cfg_r = io_ptw_pmp_5_cfg_r; // @[TLB.scala 193:14:freechips.rocketchip.system.DefaultRV32Config.fir@198449.4]
  assign pmp_io_pmp_5_addr = io_ptw_pmp_5_addr; // @[TLB.scala 193:14:freechips.rocketchip.system.DefaultRV32Config.fir@198449.4]
  assign pmp_io_pmp_5_mask = io_ptw_pmp_5_mask; // @[TLB.scala 193:14:freechips.rocketchip.system.DefaultRV32Config.fir@198449.4]
  assign pmp_io_pmp_6_cfg_l = io_ptw_pmp_6_cfg_l; // @[TLB.scala 193:14:freechips.rocketchip.system.DefaultRV32Config.fir@198450.4]
  assign pmp_io_pmp_6_cfg_a = io_ptw_pmp_6_cfg_a; // @[TLB.scala 193:14:freechips.rocketchip.system.DefaultRV32Config.fir@198450.4]
  assign pmp_io_pmp_6_cfg_x = io_ptw_pmp_6_cfg_x; // @[TLB.scala 193:14:freechips.rocketchip.system.DefaultRV32Config.fir@198450.4]
  assign pmp_io_pmp_6_cfg_w = io_ptw_pmp_6_cfg_w; // @[TLB.scala 193:14:freechips.rocketchip.system.DefaultRV32Config.fir@198450.4]
  assign pmp_io_pmp_6_cfg_r = io_ptw_pmp_6_cfg_r; // @[TLB.scala 193:14:freechips.rocketchip.system.DefaultRV32Config.fir@198450.4]
  assign pmp_io_pmp_6_addr = io_ptw_pmp_6_addr; // @[TLB.scala 193:14:freechips.rocketchip.system.DefaultRV32Config.fir@198450.4]
  assign pmp_io_pmp_6_mask = io_ptw_pmp_6_mask; // @[TLB.scala 193:14:freechips.rocketchip.system.DefaultRV32Config.fir@198450.4]
  assign pmp_io_pmp_7_cfg_l = io_ptw_pmp_7_cfg_l; // @[TLB.scala 193:14:freechips.rocketchip.system.DefaultRV32Config.fir@198451.4]
  assign pmp_io_pmp_7_cfg_a = io_ptw_pmp_7_cfg_a; // @[TLB.scala 193:14:freechips.rocketchip.system.DefaultRV32Config.fir@198451.4]
  assign pmp_io_pmp_7_cfg_x = io_ptw_pmp_7_cfg_x; // @[TLB.scala 193:14:freechips.rocketchip.system.DefaultRV32Config.fir@198451.4]
  assign pmp_io_pmp_7_cfg_w = io_ptw_pmp_7_cfg_w; // @[TLB.scala 193:14:freechips.rocketchip.system.DefaultRV32Config.fir@198451.4]
  assign pmp_io_pmp_7_cfg_r = io_ptw_pmp_7_cfg_r; // @[TLB.scala 193:14:freechips.rocketchip.system.DefaultRV32Config.fir@198451.4]
  assign pmp_io_pmp_7_addr = io_ptw_pmp_7_addr; // @[TLB.scala 193:14:freechips.rocketchip.system.DefaultRV32Config.fir@198451.4]
  assign pmp_io_pmp_7_mask = io_ptw_pmp_7_mask; // @[TLB.scala 193:14:freechips.rocketchip.system.DefaultRV32Config.fir@198451.4]
  assign pmp_io_addr = {mpu_ppn,io_req_bits_vaddr[11:0]}; // @[TLB.scala 191:15:freechips.rocketchip.system.DefaultRV32Config.fir@198442.4]
  assign OptimizationBarrier_1_io_x_ppn = _GEN_35[34:15]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@199143.4]
  assign OptimizationBarrier_1_io_x_u = _GEN_35[14]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@199143.4]
  assign OptimizationBarrier_1_io_x_ae = _GEN_35[12]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@199143.4]
  assign OptimizationBarrier_1_io_x_sw = _GEN_35[11]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@199143.4]
  assign OptimizationBarrier_1_io_x_sx = _GEN_35[10]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@199143.4]
  assign OptimizationBarrier_1_io_x_sr = _GEN_35[9]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@199143.4]
  assign OptimizationBarrier_1_io_x_pw = _GEN_35[8]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@199143.4]
  assign OptimizationBarrier_1_io_x_px = _GEN_35[7]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@199143.4]
  assign OptimizationBarrier_1_io_x_pr = _GEN_35[6]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@199143.4]
  assign OptimizationBarrier_1_io_x_ppp = _GEN_35[5]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@199143.4]
  assign OptimizationBarrier_1_io_x_pal = _GEN_35[4]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@199143.4]
  assign OptimizationBarrier_1_io_x_paa = _GEN_35[3]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@199143.4]
  assign OptimizationBarrier_1_io_x_eff = _GEN_35[2]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@199143.4]
  assign OptimizationBarrier_1_io_x_c = _GEN_35[1]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@199143.4]
  assign OptimizationBarrier_2_io_x_ppn = _GEN_39[34:15]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@199186.4]
  assign OptimizationBarrier_2_io_x_u = _GEN_39[14]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@199186.4]
  assign OptimizationBarrier_2_io_x_ae = _GEN_39[12]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@199186.4]
  assign OptimizationBarrier_2_io_x_sw = _GEN_39[11]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@199186.4]
  assign OptimizationBarrier_2_io_x_sx = _GEN_39[10]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@199186.4]
  assign OptimizationBarrier_2_io_x_sr = _GEN_39[9]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@199186.4]
  assign OptimizationBarrier_2_io_x_pw = _GEN_39[8]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@199186.4]
  assign OptimizationBarrier_2_io_x_px = _GEN_39[7]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@199186.4]
  assign OptimizationBarrier_2_io_x_pr = _GEN_39[6]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@199186.4]
  assign OptimizationBarrier_2_io_x_ppp = _GEN_39[5]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@199186.4]
  assign OptimizationBarrier_2_io_x_pal = _GEN_39[4]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@199186.4]
  assign OptimizationBarrier_2_io_x_paa = _GEN_39[3]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@199186.4]
  assign OptimizationBarrier_2_io_x_eff = _GEN_39[2]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@199186.4]
  assign OptimizationBarrier_2_io_x_c = _GEN_39[1]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@199186.4]
  assign OptimizationBarrier_3_io_x_ppn = _GEN_43[34:15]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@199229.4]
  assign OptimizationBarrier_3_io_x_u = _GEN_43[14]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@199229.4]
  assign OptimizationBarrier_3_io_x_ae = _GEN_43[12]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@199229.4]
  assign OptimizationBarrier_3_io_x_sw = _GEN_43[11]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@199229.4]
  assign OptimizationBarrier_3_io_x_sx = _GEN_43[10]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@199229.4]
  assign OptimizationBarrier_3_io_x_sr = _GEN_43[9]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@199229.4]
  assign OptimizationBarrier_3_io_x_pw = _GEN_43[8]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@199229.4]
  assign OptimizationBarrier_3_io_x_px = _GEN_43[7]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@199229.4]
  assign OptimizationBarrier_3_io_x_pr = _GEN_43[6]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@199229.4]
  assign OptimizationBarrier_3_io_x_ppp = _GEN_43[5]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@199229.4]
  assign OptimizationBarrier_3_io_x_pal = _GEN_43[4]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@199229.4]
  assign OptimizationBarrier_3_io_x_paa = _GEN_43[3]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@199229.4]
  assign OptimizationBarrier_3_io_x_eff = _GEN_43[2]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@199229.4]
  assign OptimizationBarrier_3_io_x_c = _GEN_43[1]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@199229.4]
  assign OptimizationBarrier_4_io_x_ppn = _GEN_47[34:15]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@199272.4]
  assign OptimizationBarrier_4_io_x_u = _GEN_47[14]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@199272.4]
  assign OptimizationBarrier_4_io_x_ae = _GEN_47[12]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@199272.4]
  assign OptimizationBarrier_4_io_x_sw = _GEN_47[11]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@199272.4]
  assign OptimizationBarrier_4_io_x_sx = _GEN_47[10]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@199272.4]
  assign OptimizationBarrier_4_io_x_sr = _GEN_47[9]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@199272.4]
  assign OptimizationBarrier_4_io_x_pw = _GEN_47[8]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@199272.4]
  assign OptimizationBarrier_4_io_x_px = _GEN_47[7]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@199272.4]
  assign OptimizationBarrier_4_io_x_pr = _GEN_47[6]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@199272.4]
  assign OptimizationBarrier_4_io_x_ppp = _GEN_47[5]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@199272.4]
  assign OptimizationBarrier_4_io_x_pal = _GEN_47[4]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@199272.4]
  assign OptimizationBarrier_4_io_x_paa = _GEN_47[3]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@199272.4]
  assign OptimizationBarrier_4_io_x_eff = _GEN_47[2]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@199272.4]
  assign OptimizationBarrier_4_io_x_c = _GEN_47[1]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@199272.4]
  assign OptimizationBarrier_5_io_x_ppn = _GEN_51[34:15]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@199315.4]
  assign OptimizationBarrier_5_io_x_u = _GEN_51[14]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@199315.4]
  assign OptimizationBarrier_5_io_x_ae = _GEN_51[12]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@199315.4]
  assign OptimizationBarrier_5_io_x_sw = _GEN_51[11]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@199315.4]
  assign OptimizationBarrier_5_io_x_sx = _GEN_51[10]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@199315.4]
  assign OptimizationBarrier_5_io_x_sr = _GEN_51[9]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@199315.4]
  assign OptimizationBarrier_5_io_x_pw = _GEN_51[8]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@199315.4]
  assign OptimizationBarrier_5_io_x_px = _GEN_51[7]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@199315.4]
  assign OptimizationBarrier_5_io_x_pr = _GEN_51[6]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@199315.4]
  assign OptimizationBarrier_5_io_x_ppp = _GEN_51[5]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@199315.4]
  assign OptimizationBarrier_5_io_x_pal = _GEN_51[4]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@199315.4]
  assign OptimizationBarrier_5_io_x_paa = _GEN_51[3]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@199315.4]
  assign OptimizationBarrier_5_io_x_eff = _GEN_51[2]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@199315.4]
  assign OptimizationBarrier_5_io_x_c = _GEN_51[1]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@199315.4]
  assign OptimizationBarrier_6_io_x_ppn = _GEN_55[34:15]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@199358.4]
  assign OptimizationBarrier_6_io_x_u = _GEN_55[14]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@199358.4]
  assign OptimizationBarrier_6_io_x_ae = _GEN_55[12]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@199358.4]
  assign OptimizationBarrier_6_io_x_sw = _GEN_55[11]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@199358.4]
  assign OptimizationBarrier_6_io_x_sx = _GEN_55[10]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@199358.4]
  assign OptimizationBarrier_6_io_x_sr = _GEN_55[9]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@199358.4]
  assign OptimizationBarrier_6_io_x_pw = _GEN_55[8]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@199358.4]
  assign OptimizationBarrier_6_io_x_px = _GEN_55[7]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@199358.4]
  assign OptimizationBarrier_6_io_x_pr = _GEN_55[6]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@199358.4]
  assign OptimizationBarrier_6_io_x_ppp = _GEN_55[5]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@199358.4]
  assign OptimizationBarrier_6_io_x_pal = _GEN_55[4]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@199358.4]
  assign OptimizationBarrier_6_io_x_paa = _GEN_55[3]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@199358.4]
  assign OptimizationBarrier_6_io_x_eff = _GEN_55[2]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@199358.4]
  assign OptimizationBarrier_6_io_x_c = _GEN_55[1]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@199358.4]
  assign OptimizationBarrier_7_io_x_ppn = _GEN_59[34:15]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@199401.4]
  assign OptimizationBarrier_7_io_x_u = _GEN_59[14]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@199401.4]
  assign OptimizationBarrier_7_io_x_ae = _GEN_59[12]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@199401.4]
  assign OptimizationBarrier_7_io_x_sw = _GEN_59[11]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@199401.4]
  assign OptimizationBarrier_7_io_x_sx = _GEN_59[10]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@199401.4]
  assign OptimizationBarrier_7_io_x_sr = _GEN_59[9]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@199401.4]
  assign OptimizationBarrier_7_io_x_pw = _GEN_59[8]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@199401.4]
  assign OptimizationBarrier_7_io_x_px = _GEN_59[7]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@199401.4]
  assign OptimizationBarrier_7_io_x_pr = _GEN_59[6]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@199401.4]
  assign OptimizationBarrier_7_io_x_ppp = _GEN_59[5]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@199401.4]
  assign OptimizationBarrier_7_io_x_pal = _GEN_59[4]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@199401.4]
  assign OptimizationBarrier_7_io_x_paa = _GEN_59[3]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@199401.4]
  assign OptimizationBarrier_7_io_x_eff = _GEN_59[2]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@199401.4]
  assign OptimizationBarrier_7_io_x_c = _GEN_59[1]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@199401.4]
  assign OptimizationBarrier_8_io_x_ppn = _GEN_63[34:15]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@199444.4]
  assign OptimizationBarrier_8_io_x_u = _GEN_63[14]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@199444.4]
  assign OptimizationBarrier_8_io_x_ae = _GEN_63[12]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@199444.4]
  assign OptimizationBarrier_8_io_x_sw = _GEN_63[11]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@199444.4]
  assign OptimizationBarrier_8_io_x_sx = _GEN_63[10]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@199444.4]
  assign OptimizationBarrier_8_io_x_sr = _GEN_63[9]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@199444.4]
  assign OptimizationBarrier_8_io_x_pw = _GEN_63[8]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@199444.4]
  assign OptimizationBarrier_8_io_x_px = _GEN_63[7]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@199444.4]
  assign OptimizationBarrier_8_io_x_pr = _GEN_63[6]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@199444.4]
  assign OptimizationBarrier_8_io_x_ppp = _GEN_63[5]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@199444.4]
  assign OptimizationBarrier_8_io_x_pal = _GEN_63[4]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@199444.4]
  assign OptimizationBarrier_8_io_x_paa = _GEN_63[3]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@199444.4]
  assign OptimizationBarrier_8_io_x_eff = _GEN_63[2]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@199444.4]
  assign OptimizationBarrier_8_io_x_c = _GEN_63[1]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@199444.4]
  assign OptimizationBarrier_9_io_x_ppn = superpage_entries_0_data_0[34:15]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@199486.4]
  assign OptimizationBarrier_9_io_x_u = superpage_entries_0_data_0[14]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@199486.4]
  assign OptimizationBarrier_9_io_x_ae = superpage_entries_0_data_0[12]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@199486.4]
  assign OptimizationBarrier_9_io_x_sw = superpage_entries_0_data_0[11]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@199486.4]
  assign OptimizationBarrier_9_io_x_sx = superpage_entries_0_data_0[10]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@199486.4]
  assign OptimizationBarrier_9_io_x_sr = superpage_entries_0_data_0[9]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@199486.4]
  assign OptimizationBarrier_9_io_x_pw = superpage_entries_0_data_0[8]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@199486.4]
  assign OptimizationBarrier_9_io_x_px = superpage_entries_0_data_0[7]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@199486.4]
  assign OptimizationBarrier_9_io_x_pr = superpage_entries_0_data_0[6]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@199486.4]
  assign OptimizationBarrier_9_io_x_ppp = superpage_entries_0_data_0[5]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@199486.4]
  assign OptimizationBarrier_9_io_x_pal = superpage_entries_0_data_0[4]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@199486.4]
  assign OptimizationBarrier_9_io_x_paa = superpage_entries_0_data_0[3]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@199486.4]
  assign OptimizationBarrier_9_io_x_eff = superpage_entries_0_data_0[2]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@199486.4]
  assign OptimizationBarrier_9_io_x_c = superpage_entries_0_data_0[1]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@199486.4]
  assign OptimizationBarrier_10_io_x_ppn = superpage_entries_1_data_0[34:15]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@199535.4]
  assign OptimizationBarrier_10_io_x_u = superpage_entries_1_data_0[14]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@199535.4]
  assign OptimizationBarrier_10_io_x_ae = superpage_entries_1_data_0[12]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@199535.4]
  assign OptimizationBarrier_10_io_x_sw = superpage_entries_1_data_0[11]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@199535.4]
  assign OptimizationBarrier_10_io_x_sx = superpage_entries_1_data_0[10]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@199535.4]
  assign OptimizationBarrier_10_io_x_sr = superpage_entries_1_data_0[9]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@199535.4]
  assign OptimizationBarrier_10_io_x_pw = superpage_entries_1_data_0[8]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@199535.4]
  assign OptimizationBarrier_10_io_x_px = superpage_entries_1_data_0[7]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@199535.4]
  assign OptimizationBarrier_10_io_x_pr = superpage_entries_1_data_0[6]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@199535.4]
  assign OptimizationBarrier_10_io_x_ppp = superpage_entries_1_data_0[5]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@199535.4]
  assign OptimizationBarrier_10_io_x_pal = superpage_entries_1_data_0[4]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@199535.4]
  assign OptimizationBarrier_10_io_x_paa = superpage_entries_1_data_0[3]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@199535.4]
  assign OptimizationBarrier_10_io_x_eff = superpage_entries_1_data_0[2]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@199535.4]
  assign OptimizationBarrier_10_io_x_c = superpage_entries_1_data_0[1]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@199535.4]
  assign OptimizationBarrier_11_io_x_ppn = superpage_entries_2_data_0[34:15]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@199584.4]
  assign OptimizationBarrier_11_io_x_u = superpage_entries_2_data_0[14]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@199584.4]
  assign OptimizationBarrier_11_io_x_ae = superpage_entries_2_data_0[12]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@199584.4]
  assign OptimizationBarrier_11_io_x_sw = superpage_entries_2_data_0[11]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@199584.4]
  assign OptimizationBarrier_11_io_x_sx = superpage_entries_2_data_0[10]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@199584.4]
  assign OptimizationBarrier_11_io_x_sr = superpage_entries_2_data_0[9]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@199584.4]
  assign OptimizationBarrier_11_io_x_pw = superpage_entries_2_data_0[8]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@199584.4]
  assign OptimizationBarrier_11_io_x_px = superpage_entries_2_data_0[7]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@199584.4]
  assign OptimizationBarrier_11_io_x_pr = superpage_entries_2_data_0[6]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@199584.4]
  assign OptimizationBarrier_11_io_x_ppp = superpage_entries_2_data_0[5]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@199584.4]
  assign OptimizationBarrier_11_io_x_pal = superpage_entries_2_data_0[4]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@199584.4]
  assign OptimizationBarrier_11_io_x_paa = superpage_entries_2_data_0[3]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@199584.4]
  assign OptimizationBarrier_11_io_x_eff = superpage_entries_2_data_0[2]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@199584.4]
  assign OptimizationBarrier_11_io_x_c = superpage_entries_2_data_0[1]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@199584.4]
  assign OptimizationBarrier_12_io_x_ppn = superpage_entries_3_data_0[34:15]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@199633.4]
  assign OptimizationBarrier_12_io_x_u = superpage_entries_3_data_0[14]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@199633.4]
  assign OptimizationBarrier_12_io_x_ae = superpage_entries_3_data_0[12]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@199633.4]
  assign OptimizationBarrier_12_io_x_sw = superpage_entries_3_data_0[11]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@199633.4]
  assign OptimizationBarrier_12_io_x_sx = superpage_entries_3_data_0[10]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@199633.4]
  assign OptimizationBarrier_12_io_x_sr = superpage_entries_3_data_0[9]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@199633.4]
  assign OptimizationBarrier_12_io_x_pw = superpage_entries_3_data_0[8]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@199633.4]
  assign OptimizationBarrier_12_io_x_px = superpage_entries_3_data_0[7]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@199633.4]
  assign OptimizationBarrier_12_io_x_pr = superpage_entries_3_data_0[6]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@199633.4]
  assign OptimizationBarrier_12_io_x_ppp = superpage_entries_3_data_0[5]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@199633.4]
  assign OptimizationBarrier_12_io_x_pal = superpage_entries_3_data_0[4]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@199633.4]
  assign OptimizationBarrier_12_io_x_paa = superpage_entries_3_data_0[3]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@199633.4]
  assign OptimizationBarrier_12_io_x_eff = superpage_entries_3_data_0[2]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@199633.4]
  assign OptimizationBarrier_12_io_x_c = superpage_entries_3_data_0[1]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@199633.4]
  assign OptimizationBarrier_13_io_x_ppn = special_entry_data_0[34:15]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@199682.4]
  assign OptimizationBarrier_13_io_x_u = special_entry_data_0[14]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@199682.4]
  assign OptimizationBarrier_13_io_x_ae = special_entry_data_0[12]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@199682.4]
  assign OptimizationBarrier_13_io_x_sw = special_entry_data_0[11]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@199682.4]
  assign OptimizationBarrier_13_io_x_sx = special_entry_data_0[10]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@199682.4]
  assign OptimizationBarrier_13_io_x_sr = special_entry_data_0[9]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@199682.4]
  assign OptimizationBarrier_13_io_x_pw = special_entry_data_0[8]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@199682.4]
  assign OptimizationBarrier_13_io_x_px = special_entry_data_0[7]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@199682.4]
  assign OptimizationBarrier_13_io_x_pr = special_entry_data_0[6]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@199682.4]
  assign OptimizationBarrier_13_io_x_ppp = special_entry_data_0[5]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@199682.4]
  assign OptimizationBarrier_13_io_x_pal = special_entry_data_0[4]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@199682.4]
  assign OptimizationBarrier_13_io_x_paa = special_entry_data_0[3]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@199682.4]
  assign OptimizationBarrier_13_io_x_eff = special_entry_data_0[2]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@199682.4]
  assign OptimizationBarrier_13_io_x_c = special_entry_data_0[1]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@199682.4]
  assign OptimizationBarrier_14_io_x_ppn = _GEN_35[34:15]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@200163.4]
  assign OptimizationBarrier_14_io_x_u = _GEN_35[14]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@200163.4]
  assign OptimizationBarrier_14_io_x_ae = _GEN_35[12]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@200163.4]
  assign OptimizationBarrier_14_io_x_sw = _GEN_35[11]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@200163.4]
  assign OptimizationBarrier_14_io_x_sx = _GEN_35[10]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@200163.4]
  assign OptimizationBarrier_14_io_x_sr = _GEN_35[9]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@200163.4]
  assign OptimizationBarrier_14_io_x_pw = _GEN_35[8]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@200163.4]
  assign OptimizationBarrier_14_io_x_px = _GEN_35[7]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@200163.4]
  assign OptimizationBarrier_14_io_x_pr = _GEN_35[6]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@200163.4]
  assign OptimizationBarrier_14_io_x_ppp = _GEN_35[5]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@200163.4]
  assign OptimizationBarrier_14_io_x_pal = _GEN_35[4]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@200163.4]
  assign OptimizationBarrier_14_io_x_paa = _GEN_35[3]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@200163.4]
  assign OptimizationBarrier_14_io_x_eff = _GEN_35[2]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@200163.4]
  assign OptimizationBarrier_14_io_x_c = _GEN_35[1]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@200163.4]
  assign OptimizationBarrier_15_io_x_ppn = _GEN_39[34:15]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@200206.4]
  assign OptimizationBarrier_15_io_x_u = _GEN_39[14]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@200206.4]
  assign OptimizationBarrier_15_io_x_ae = _GEN_39[12]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@200206.4]
  assign OptimizationBarrier_15_io_x_sw = _GEN_39[11]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@200206.4]
  assign OptimizationBarrier_15_io_x_sx = _GEN_39[10]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@200206.4]
  assign OptimizationBarrier_15_io_x_sr = _GEN_39[9]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@200206.4]
  assign OptimizationBarrier_15_io_x_pw = _GEN_39[8]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@200206.4]
  assign OptimizationBarrier_15_io_x_px = _GEN_39[7]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@200206.4]
  assign OptimizationBarrier_15_io_x_pr = _GEN_39[6]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@200206.4]
  assign OptimizationBarrier_15_io_x_ppp = _GEN_39[5]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@200206.4]
  assign OptimizationBarrier_15_io_x_pal = _GEN_39[4]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@200206.4]
  assign OptimizationBarrier_15_io_x_paa = _GEN_39[3]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@200206.4]
  assign OptimizationBarrier_15_io_x_eff = _GEN_39[2]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@200206.4]
  assign OptimizationBarrier_15_io_x_c = _GEN_39[1]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@200206.4]
  assign OptimizationBarrier_16_io_x_ppn = _GEN_43[34:15]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@200249.4]
  assign OptimizationBarrier_16_io_x_u = _GEN_43[14]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@200249.4]
  assign OptimizationBarrier_16_io_x_ae = _GEN_43[12]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@200249.4]
  assign OptimizationBarrier_16_io_x_sw = _GEN_43[11]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@200249.4]
  assign OptimizationBarrier_16_io_x_sx = _GEN_43[10]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@200249.4]
  assign OptimizationBarrier_16_io_x_sr = _GEN_43[9]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@200249.4]
  assign OptimizationBarrier_16_io_x_pw = _GEN_43[8]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@200249.4]
  assign OptimizationBarrier_16_io_x_px = _GEN_43[7]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@200249.4]
  assign OptimizationBarrier_16_io_x_pr = _GEN_43[6]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@200249.4]
  assign OptimizationBarrier_16_io_x_ppp = _GEN_43[5]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@200249.4]
  assign OptimizationBarrier_16_io_x_pal = _GEN_43[4]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@200249.4]
  assign OptimizationBarrier_16_io_x_paa = _GEN_43[3]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@200249.4]
  assign OptimizationBarrier_16_io_x_eff = _GEN_43[2]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@200249.4]
  assign OptimizationBarrier_16_io_x_c = _GEN_43[1]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@200249.4]
  assign OptimizationBarrier_17_io_x_ppn = _GEN_47[34:15]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@200292.4]
  assign OptimizationBarrier_17_io_x_u = _GEN_47[14]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@200292.4]
  assign OptimizationBarrier_17_io_x_ae = _GEN_47[12]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@200292.4]
  assign OptimizationBarrier_17_io_x_sw = _GEN_47[11]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@200292.4]
  assign OptimizationBarrier_17_io_x_sx = _GEN_47[10]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@200292.4]
  assign OptimizationBarrier_17_io_x_sr = _GEN_47[9]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@200292.4]
  assign OptimizationBarrier_17_io_x_pw = _GEN_47[8]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@200292.4]
  assign OptimizationBarrier_17_io_x_px = _GEN_47[7]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@200292.4]
  assign OptimizationBarrier_17_io_x_pr = _GEN_47[6]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@200292.4]
  assign OptimizationBarrier_17_io_x_ppp = _GEN_47[5]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@200292.4]
  assign OptimizationBarrier_17_io_x_pal = _GEN_47[4]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@200292.4]
  assign OptimizationBarrier_17_io_x_paa = _GEN_47[3]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@200292.4]
  assign OptimizationBarrier_17_io_x_eff = _GEN_47[2]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@200292.4]
  assign OptimizationBarrier_17_io_x_c = _GEN_47[1]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@200292.4]
  assign OptimizationBarrier_18_io_x_ppn = _GEN_51[34:15]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@200335.4]
  assign OptimizationBarrier_18_io_x_u = _GEN_51[14]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@200335.4]
  assign OptimizationBarrier_18_io_x_ae = _GEN_51[12]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@200335.4]
  assign OptimizationBarrier_18_io_x_sw = _GEN_51[11]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@200335.4]
  assign OptimizationBarrier_18_io_x_sx = _GEN_51[10]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@200335.4]
  assign OptimizationBarrier_18_io_x_sr = _GEN_51[9]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@200335.4]
  assign OptimizationBarrier_18_io_x_pw = _GEN_51[8]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@200335.4]
  assign OptimizationBarrier_18_io_x_px = _GEN_51[7]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@200335.4]
  assign OptimizationBarrier_18_io_x_pr = _GEN_51[6]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@200335.4]
  assign OptimizationBarrier_18_io_x_ppp = _GEN_51[5]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@200335.4]
  assign OptimizationBarrier_18_io_x_pal = _GEN_51[4]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@200335.4]
  assign OptimizationBarrier_18_io_x_paa = _GEN_51[3]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@200335.4]
  assign OptimizationBarrier_18_io_x_eff = _GEN_51[2]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@200335.4]
  assign OptimizationBarrier_18_io_x_c = _GEN_51[1]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@200335.4]
  assign OptimizationBarrier_19_io_x_ppn = _GEN_55[34:15]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@200378.4]
  assign OptimizationBarrier_19_io_x_u = _GEN_55[14]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@200378.4]
  assign OptimizationBarrier_19_io_x_ae = _GEN_55[12]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@200378.4]
  assign OptimizationBarrier_19_io_x_sw = _GEN_55[11]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@200378.4]
  assign OptimizationBarrier_19_io_x_sx = _GEN_55[10]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@200378.4]
  assign OptimizationBarrier_19_io_x_sr = _GEN_55[9]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@200378.4]
  assign OptimizationBarrier_19_io_x_pw = _GEN_55[8]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@200378.4]
  assign OptimizationBarrier_19_io_x_px = _GEN_55[7]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@200378.4]
  assign OptimizationBarrier_19_io_x_pr = _GEN_55[6]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@200378.4]
  assign OptimizationBarrier_19_io_x_ppp = _GEN_55[5]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@200378.4]
  assign OptimizationBarrier_19_io_x_pal = _GEN_55[4]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@200378.4]
  assign OptimizationBarrier_19_io_x_paa = _GEN_55[3]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@200378.4]
  assign OptimizationBarrier_19_io_x_eff = _GEN_55[2]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@200378.4]
  assign OptimizationBarrier_19_io_x_c = _GEN_55[1]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@200378.4]
  assign OptimizationBarrier_20_io_x_ppn = _GEN_59[34:15]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@200421.4]
  assign OptimizationBarrier_20_io_x_u = _GEN_59[14]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@200421.4]
  assign OptimizationBarrier_20_io_x_ae = _GEN_59[12]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@200421.4]
  assign OptimizationBarrier_20_io_x_sw = _GEN_59[11]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@200421.4]
  assign OptimizationBarrier_20_io_x_sx = _GEN_59[10]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@200421.4]
  assign OptimizationBarrier_20_io_x_sr = _GEN_59[9]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@200421.4]
  assign OptimizationBarrier_20_io_x_pw = _GEN_59[8]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@200421.4]
  assign OptimizationBarrier_20_io_x_px = _GEN_59[7]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@200421.4]
  assign OptimizationBarrier_20_io_x_pr = _GEN_59[6]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@200421.4]
  assign OptimizationBarrier_20_io_x_ppp = _GEN_59[5]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@200421.4]
  assign OptimizationBarrier_20_io_x_pal = _GEN_59[4]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@200421.4]
  assign OptimizationBarrier_20_io_x_paa = _GEN_59[3]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@200421.4]
  assign OptimizationBarrier_20_io_x_eff = _GEN_59[2]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@200421.4]
  assign OptimizationBarrier_20_io_x_c = _GEN_59[1]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@200421.4]
  assign OptimizationBarrier_21_io_x_ppn = _GEN_63[34:15]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@200464.4]
  assign OptimizationBarrier_21_io_x_u = _GEN_63[14]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@200464.4]
  assign OptimizationBarrier_21_io_x_ae = _GEN_63[12]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@200464.4]
  assign OptimizationBarrier_21_io_x_sw = _GEN_63[11]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@200464.4]
  assign OptimizationBarrier_21_io_x_sx = _GEN_63[10]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@200464.4]
  assign OptimizationBarrier_21_io_x_sr = _GEN_63[9]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@200464.4]
  assign OptimizationBarrier_21_io_x_pw = _GEN_63[8]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@200464.4]
  assign OptimizationBarrier_21_io_x_px = _GEN_63[7]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@200464.4]
  assign OptimizationBarrier_21_io_x_pr = _GEN_63[6]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@200464.4]
  assign OptimizationBarrier_21_io_x_ppp = _GEN_63[5]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@200464.4]
  assign OptimizationBarrier_21_io_x_pal = _GEN_63[4]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@200464.4]
  assign OptimizationBarrier_21_io_x_paa = _GEN_63[3]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@200464.4]
  assign OptimizationBarrier_21_io_x_eff = _GEN_63[2]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@200464.4]
  assign OptimizationBarrier_21_io_x_c = _GEN_63[1]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@200464.4]
  assign OptimizationBarrier_22_io_x_ppn = superpage_entries_0_data_0[34:15]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@200506.4]
  assign OptimizationBarrier_22_io_x_u = superpage_entries_0_data_0[14]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@200506.4]
  assign OptimizationBarrier_22_io_x_ae = superpage_entries_0_data_0[12]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@200506.4]
  assign OptimizationBarrier_22_io_x_sw = superpage_entries_0_data_0[11]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@200506.4]
  assign OptimizationBarrier_22_io_x_sx = superpage_entries_0_data_0[10]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@200506.4]
  assign OptimizationBarrier_22_io_x_sr = superpage_entries_0_data_0[9]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@200506.4]
  assign OptimizationBarrier_22_io_x_pw = superpage_entries_0_data_0[8]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@200506.4]
  assign OptimizationBarrier_22_io_x_px = superpage_entries_0_data_0[7]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@200506.4]
  assign OptimizationBarrier_22_io_x_pr = superpage_entries_0_data_0[6]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@200506.4]
  assign OptimizationBarrier_22_io_x_ppp = superpage_entries_0_data_0[5]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@200506.4]
  assign OptimizationBarrier_22_io_x_pal = superpage_entries_0_data_0[4]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@200506.4]
  assign OptimizationBarrier_22_io_x_paa = superpage_entries_0_data_0[3]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@200506.4]
  assign OptimizationBarrier_22_io_x_eff = superpage_entries_0_data_0[2]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@200506.4]
  assign OptimizationBarrier_22_io_x_c = superpage_entries_0_data_0[1]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@200506.4]
  assign OptimizationBarrier_23_io_x_ppn = superpage_entries_1_data_0[34:15]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@200548.4]
  assign OptimizationBarrier_23_io_x_u = superpage_entries_1_data_0[14]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@200548.4]
  assign OptimizationBarrier_23_io_x_ae = superpage_entries_1_data_0[12]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@200548.4]
  assign OptimizationBarrier_23_io_x_sw = superpage_entries_1_data_0[11]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@200548.4]
  assign OptimizationBarrier_23_io_x_sx = superpage_entries_1_data_0[10]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@200548.4]
  assign OptimizationBarrier_23_io_x_sr = superpage_entries_1_data_0[9]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@200548.4]
  assign OptimizationBarrier_23_io_x_pw = superpage_entries_1_data_0[8]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@200548.4]
  assign OptimizationBarrier_23_io_x_px = superpage_entries_1_data_0[7]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@200548.4]
  assign OptimizationBarrier_23_io_x_pr = superpage_entries_1_data_0[6]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@200548.4]
  assign OptimizationBarrier_23_io_x_ppp = superpage_entries_1_data_0[5]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@200548.4]
  assign OptimizationBarrier_23_io_x_pal = superpage_entries_1_data_0[4]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@200548.4]
  assign OptimizationBarrier_23_io_x_paa = superpage_entries_1_data_0[3]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@200548.4]
  assign OptimizationBarrier_23_io_x_eff = superpage_entries_1_data_0[2]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@200548.4]
  assign OptimizationBarrier_23_io_x_c = superpage_entries_1_data_0[1]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@200548.4]
  assign OptimizationBarrier_24_io_x_ppn = superpage_entries_2_data_0[34:15]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@200590.4]
  assign OptimizationBarrier_24_io_x_u = superpage_entries_2_data_0[14]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@200590.4]
  assign OptimizationBarrier_24_io_x_ae = superpage_entries_2_data_0[12]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@200590.4]
  assign OptimizationBarrier_24_io_x_sw = superpage_entries_2_data_0[11]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@200590.4]
  assign OptimizationBarrier_24_io_x_sx = superpage_entries_2_data_0[10]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@200590.4]
  assign OptimizationBarrier_24_io_x_sr = superpage_entries_2_data_0[9]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@200590.4]
  assign OptimizationBarrier_24_io_x_pw = superpage_entries_2_data_0[8]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@200590.4]
  assign OptimizationBarrier_24_io_x_px = superpage_entries_2_data_0[7]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@200590.4]
  assign OptimizationBarrier_24_io_x_pr = superpage_entries_2_data_0[6]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@200590.4]
  assign OptimizationBarrier_24_io_x_ppp = superpage_entries_2_data_0[5]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@200590.4]
  assign OptimizationBarrier_24_io_x_pal = superpage_entries_2_data_0[4]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@200590.4]
  assign OptimizationBarrier_24_io_x_paa = superpage_entries_2_data_0[3]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@200590.4]
  assign OptimizationBarrier_24_io_x_eff = superpage_entries_2_data_0[2]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@200590.4]
  assign OptimizationBarrier_24_io_x_c = superpage_entries_2_data_0[1]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@200590.4]
  assign OptimizationBarrier_25_io_x_ppn = superpage_entries_3_data_0[34:15]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@200632.4]
  assign OptimizationBarrier_25_io_x_u = superpage_entries_3_data_0[14]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@200632.4]
  assign OptimizationBarrier_25_io_x_ae = superpage_entries_3_data_0[12]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@200632.4]
  assign OptimizationBarrier_25_io_x_sw = superpage_entries_3_data_0[11]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@200632.4]
  assign OptimizationBarrier_25_io_x_sx = superpage_entries_3_data_0[10]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@200632.4]
  assign OptimizationBarrier_25_io_x_sr = superpage_entries_3_data_0[9]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@200632.4]
  assign OptimizationBarrier_25_io_x_pw = superpage_entries_3_data_0[8]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@200632.4]
  assign OptimizationBarrier_25_io_x_px = superpage_entries_3_data_0[7]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@200632.4]
  assign OptimizationBarrier_25_io_x_pr = superpage_entries_3_data_0[6]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@200632.4]
  assign OptimizationBarrier_25_io_x_ppp = superpage_entries_3_data_0[5]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@200632.4]
  assign OptimizationBarrier_25_io_x_pal = superpage_entries_3_data_0[4]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@200632.4]
  assign OptimizationBarrier_25_io_x_paa = superpage_entries_3_data_0[3]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@200632.4]
  assign OptimizationBarrier_25_io_x_eff = superpage_entries_3_data_0[2]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@200632.4]
  assign OptimizationBarrier_25_io_x_c = superpage_entries_3_data_0[1]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@200632.4]
  assign OptimizationBarrier_26_io_x_ppn = special_entry_data_0[34:15]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@200674.4]
  assign OptimizationBarrier_26_io_x_u = special_entry_data_0[14]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@200674.4]
  assign OptimizationBarrier_26_io_x_ae = special_entry_data_0[12]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@200674.4]
  assign OptimizationBarrier_26_io_x_sw = special_entry_data_0[11]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@200674.4]
  assign OptimizationBarrier_26_io_x_sx = special_entry_data_0[10]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@200674.4]
  assign OptimizationBarrier_26_io_x_sr = special_entry_data_0[9]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@200674.4]
  assign OptimizationBarrier_26_io_x_pw = special_entry_data_0[8]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@200674.4]
  assign OptimizationBarrier_26_io_x_px = special_entry_data_0[7]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@200674.4]
  assign OptimizationBarrier_26_io_x_pr = special_entry_data_0[6]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@200674.4]
  assign OptimizationBarrier_26_io_x_ppp = special_entry_data_0[5]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@200674.4]
  assign OptimizationBarrier_26_io_x_pal = special_entry_data_0[4]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@200674.4]
  assign OptimizationBarrier_26_io_x_paa = special_entry_data_0[3]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@200674.4]
  assign OptimizationBarrier_26_io_x_eff = special_entry_data_0[2]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@200674.4]
  assign OptimizationBarrier_26_io_x_c = special_entry_data_0[1]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@200674.4]
  assign OptimizationBarrier_27_io_x_ppn = _GEN_35[34:15]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@200717.4]
  assign OptimizationBarrier_27_io_x_u = _GEN_35[14]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@200717.4]
  assign OptimizationBarrier_27_io_x_ae = _GEN_35[12]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@200717.4]
  assign OptimizationBarrier_27_io_x_sw = _GEN_35[11]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@200717.4]
  assign OptimizationBarrier_27_io_x_sx = _GEN_35[10]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@200717.4]
  assign OptimizationBarrier_27_io_x_sr = _GEN_35[9]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@200717.4]
  assign OptimizationBarrier_27_io_x_pw = _GEN_35[8]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@200717.4]
  assign OptimizationBarrier_27_io_x_px = _GEN_35[7]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@200717.4]
  assign OptimizationBarrier_27_io_x_pr = _GEN_35[6]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@200717.4]
  assign OptimizationBarrier_27_io_x_ppp = _GEN_35[5]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@200717.4]
  assign OptimizationBarrier_27_io_x_pal = _GEN_35[4]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@200717.4]
  assign OptimizationBarrier_27_io_x_paa = _GEN_35[3]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@200717.4]
  assign OptimizationBarrier_27_io_x_eff = _GEN_35[2]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@200717.4]
  assign OptimizationBarrier_27_io_x_c = _GEN_35[1]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@200717.4]
  assign OptimizationBarrier_28_io_x_ppn = _GEN_39[34:15]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@200760.4]
  assign OptimizationBarrier_28_io_x_u = _GEN_39[14]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@200760.4]
  assign OptimizationBarrier_28_io_x_ae = _GEN_39[12]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@200760.4]
  assign OptimizationBarrier_28_io_x_sw = _GEN_39[11]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@200760.4]
  assign OptimizationBarrier_28_io_x_sx = _GEN_39[10]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@200760.4]
  assign OptimizationBarrier_28_io_x_sr = _GEN_39[9]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@200760.4]
  assign OptimizationBarrier_28_io_x_pw = _GEN_39[8]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@200760.4]
  assign OptimizationBarrier_28_io_x_px = _GEN_39[7]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@200760.4]
  assign OptimizationBarrier_28_io_x_pr = _GEN_39[6]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@200760.4]
  assign OptimizationBarrier_28_io_x_ppp = _GEN_39[5]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@200760.4]
  assign OptimizationBarrier_28_io_x_pal = _GEN_39[4]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@200760.4]
  assign OptimizationBarrier_28_io_x_paa = _GEN_39[3]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@200760.4]
  assign OptimizationBarrier_28_io_x_eff = _GEN_39[2]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@200760.4]
  assign OptimizationBarrier_28_io_x_c = _GEN_39[1]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@200760.4]
  assign OptimizationBarrier_29_io_x_ppn = _GEN_43[34:15]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@200803.4]
  assign OptimizationBarrier_29_io_x_u = _GEN_43[14]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@200803.4]
  assign OptimizationBarrier_29_io_x_ae = _GEN_43[12]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@200803.4]
  assign OptimizationBarrier_29_io_x_sw = _GEN_43[11]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@200803.4]
  assign OptimizationBarrier_29_io_x_sx = _GEN_43[10]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@200803.4]
  assign OptimizationBarrier_29_io_x_sr = _GEN_43[9]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@200803.4]
  assign OptimizationBarrier_29_io_x_pw = _GEN_43[8]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@200803.4]
  assign OptimizationBarrier_29_io_x_px = _GEN_43[7]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@200803.4]
  assign OptimizationBarrier_29_io_x_pr = _GEN_43[6]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@200803.4]
  assign OptimizationBarrier_29_io_x_ppp = _GEN_43[5]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@200803.4]
  assign OptimizationBarrier_29_io_x_pal = _GEN_43[4]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@200803.4]
  assign OptimizationBarrier_29_io_x_paa = _GEN_43[3]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@200803.4]
  assign OptimizationBarrier_29_io_x_eff = _GEN_43[2]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@200803.4]
  assign OptimizationBarrier_29_io_x_c = _GEN_43[1]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@200803.4]
  assign OptimizationBarrier_30_io_x_ppn = _GEN_47[34:15]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@200846.4]
  assign OptimizationBarrier_30_io_x_u = _GEN_47[14]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@200846.4]
  assign OptimizationBarrier_30_io_x_ae = _GEN_47[12]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@200846.4]
  assign OptimizationBarrier_30_io_x_sw = _GEN_47[11]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@200846.4]
  assign OptimizationBarrier_30_io_x_sx = _GEN_47[10]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@200846.4]
  assign OptimizationBarrier_30_io_x_sr = _GEN_47[9]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@200846.4]
  assign OptimizationBarrier_30_io_x_pw = _GEN_47[8]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@200846.4]
  assign OptimizationBarrier_30_io_x_px = _GEN_47[7]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@200846.4]
  assign OptimizationBarrier_30_io_x_pr = _GEN_47[6]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@200846.4]
  assign OptimizationBarrier_30_io_x_ppp = _GEN_47[5]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@200846.4]
  assign OptimizationBarrier_30_io_x_pal = _GEN_47[4]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@200846.4]
  assign OptimizationBarrier_30_io_x_paa = _GEN_47[3]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@200846.4]
  assign OptimizationBarrier_30_io_x_eff = _GEN_47[2]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@200846.4]
  assign OptimizationBarrier_30_io_x_c = _GEN_47[1]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@200846.4]
  assign OptimizationBarrier_31_io_x_ppn = _GEN_51[34:15]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@200889.4]
  assign OptimizationBarrier_31_io_x_u = _GEN_51[14]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@200889.4]
  assign OptimizationBarrier_31_io_x_ae = _GEN_51[12]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@200889.4]
  assign OptimizationBarrier_31_io_x_sw = _GEN_51[11]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@200889.4]
  assign OptimizationBarrier_31_io_x_sx = _GEN_51[10]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@200889.4]
  assign OptimizationBarrier_31_io_x_sr = _GEN_51[9]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@200889.4]
  assign OptimizationBarrier_31_io_x_pw = _GEN_51[8]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@200889.4]
  assign OptimizationBarrier_31_io_x_px = _GEN_51[7]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@200889.4]
  assign OptimizationBarrier_31_io_x_pr = _GEN_51[6]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@200889.4]
  assign OptimizationBarrier_31_io_x_ppp = _GEN_51[5]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@200889.4]
  assign OptimizationBarrier_31_io_x_pal = _GEN_51[4]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@200889.4]
  assign OptimizationBarrier_31_io_x_paa = _GEN_51[3]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@200889.4]
  assign OptimizationBarrier_31_io_x_eff = _GEN_51[2]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@200889.4]
  assign OptimizationBarrier_31_io_x_c = _GEN_51[1]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@200889.4]
  assign OptimizationBarrier_32_io_x_ppn = _GEN_55[34:15]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@200932.4]
  assign OptimizationBarrier_32_io_x_u = _GEN_55[14]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@200932.4]
  assign OptimizationBarrier_32_io_x_ae = _GEN_55[12]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@200932.4]
  assign OptimizationBarrier_32_io_x_sw = _GEN_55[11]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@200932.4]
  assign OptimizationBarrier_32_io_x_sx = _GEN_55[10]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@200932.4]
  assign OptimizationBarrier_32_io_x_sr = _GEN_55[9]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@200932.4]
  assign OptimizationBarrier_32_io_x_pw = _GEN_55[8]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@200932.4]
  assign OptimizationBarrier_32_io_x_px = _GEN_55[7]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@200932.4]
  assign OptimizationBarrier_32_io_x_pr = _GEN_55[6]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@200932.4]
  assign OptimizationBarrier_32_io_x_ppp = _GEN_55[5]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@200932.4]
  assign OptimizationBarrier_32_io_x_pal = _GEN_55[4]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@200932.4]
  assign OptimizationBarrier_32_io_x_paa = _GEN_55[3]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@200932.4]
  assign OptimizationBarrier_32_io_x_eff = _GEN_55[2]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@200932.4]
  assign OptimizationBarrier_32_io_x_c = _GEN_55[1]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@200932.4]
  assign OptimizationBarrier_33_io_x_ppn = _GEN_59[34:15]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@200975.4]
  assign OptimizationBarrier_33_io_x_u = _GEN_59[14]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@200975.4]
  assign OptimizationBarrier_33_io_x_ae = _GEN_59[12]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@200975.4]
  assign OptimizationBarrier_33_io_x_sw = _GEN_59[11]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@200975.4]
  assign OptimizationBarrier_33_io_x_sx = _GEN_59[10]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@200975.4]
  assign OptimizationBarrier_33_io_x_sr = _GEN_59[9]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@200975.4]
  assign OptimizationBarrier_33_io_x_pw = _GEN_59[8]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@200975.4]
  assign OptimizationBarrier_33_io_x_px = _GEN_59[7]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@200975.4]
  assign OptimizationBarrier_33_io_x_pr = _GEN_59[6]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@200975.4]
  assign OptimizationBarrier_33_io_x_ppp = _GEN_59[5]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@200975.4]
  assign OptimizationBarrier_33_io_x_pal = _GEN_59[4]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@200975.4]
  assign OptimizationBarrier_33_io_x_paa = _GEN_59[3]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@200975.4]
  assign OptimizationBarrier_33_io_x_eff = _GEN_59[2]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@200975.4]
  assign OptimizationBarrier_33_io_x_c = _GEN_59[1]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@200975.4]
  assign OptimizationBarrier_34_io_x_ppn = _GEN_63[34:15]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@201018.4]
  assign OptimizationBarrier_34_io_x_u = _GEN_63[14]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@201018.4]
  assign OptimizationBarrier_34_io_x_ae = _GEN_63[12]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@201018.4]
  assign OptimizationBarrier_34_io_x_sw = _GEN_63[11]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@201018.4]
  assign OptimizationBarrier_34_io_x_sx = _GEN_63[10]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@201018.4]
  assign OptimizationBarrier_34_io_x_sr = _GEN_63[9]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@201018.4]
  assign OptimizationBarrier_34_io_x_pw = _GEN_63[8]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@201018.4]
  assign OptimizationBarrier_34_io_x_px = _GEN_63[7]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@201018.4]
  assign OptimizationBarrier_34_io_x_pr = _GEN_63[6]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@201018.4]
  assign OptimizationBarrier_34_io_x_ppp = _GEN_63[5]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@201018.4]
  assign OptimizationBarrier_34_io_x_pal = _GEN_63[4]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@201018.4]
  assign OptimizationBarrier_34_io_x_paa = _GEN_63[3]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@201018.4]
  assign OptimizationBarrier_34_io_x_eff = _GEN_63[2]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@201018.4]
  assign OptimizationBarrier_34_io_x_c = _GEN_63[1]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@201018.4]
  assign OptimizationBarrier_35_io_x_ppn = superpage_entries_0_data_0[34:15]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@201060.4]
  assign OptimizationBarrier_35_io_x_u = superpage_entries_0_data_0[14]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@201060.4]
  assign OptimizationBarrier_35_io_x_ae = superpage_entries_0_data_0[12]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@201060.4]
  assign OptimizationBarrier_35_io_x_sw = superpage_entries_0_data_0[11]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@201060.4]
  assign OptimizationBarrier_35_io_x_sx = superpage_entries_0_data_0[10]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@201060.4]
  assign OptimizationBarrier_35_io_x_sr = superpage_entries_0_data_0[9]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@201060.4]
  assign OptimizationBarrier_35_io_x_pw = superpage_entries_0_data_0[8]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@201060.4]
  assign OptimizationBarrier_35_io_x_px = superpage_entries_0_data_0[7]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@201060.4]
  assign OptimizationBarrier_35_io_x_pr = superpage_entries_0_data_0[6]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@201060.4]
  assign OptimizationBarrier_35_io_x_ppp = superpage_entries_0_data_0[5]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@201060.4]
  assign OptimizationBarrier_35_io_x_pal = superpage_entries_0_data_0[4]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@201060.4]
  assign OptimizationBarrier_35_io_x_paa = superpage_entries_0_data_0[3]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@201060.4]
  assign OptimizationBarrier_35_io_x_eff = superpage_entries_0_data_0[2]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@201060.4]
  assign OptimizationBarrier_35_io_x_c = superpage_entries_0_data_0[1]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@201060.4]
  assign OptimizationBarrier_36_io_x_ppn = superpage_entries_1_data_0[34:15]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@201102.4]
  assign OptimizationBarrier_36_io_x_u = superpage_entries_1_data_0[14]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@201102.4]
  assign OptimizationBarrier_36_io_x_ae = superpage_entries_1_data_0[12]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@201102.4]
  assign OptimizationBarrier_36_io_x_sw = superpage_entries_1_data_0[11]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@201102.4]
  assign OptimizationBarrier_36_io_x_sx = superpage_entries_1_data_0[10]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@201102.4]
  assign OptimizationBarrier_36_io_x_sr = superpage_entries_1_data_0[9]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@201102.4]
  assign OptimizationBarrier_36_io_x_pw = superpage_entries_1_data_0[8]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@201102.4]
  assign OptimizationBarrier_36_io_x_px = superpage_entries_1_data_0[7]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@201102.4]
  assign OptimizationBarrier_36_io_x_pr = superpage_entries_1_data_0[6]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@201102.4]
  assign OptimizationBarrier_36_io_x_ppp = superpage_entries_1_data_0[5]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@201102.4]
  assign OptimizationBarrier_36_io_x_pal = superpage_entries_1_data_0[4]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@201102.4]
  assign OptimizationBarrier_36_io_x_paa = superpage_entries_1_data_0[3]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@201102.4]
  assign OptimizationBarrier_36_io_x_eff = superpage_entries_1_data_0[2]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@201102.4]
  assign OptimizationBarrier_36_io_x_c = superpage_entries_1_data_0[1]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@201102.4]
  assign OptimizationBarrier_37_io_x_ppn = superpage_entries_2_data_0[34:15]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@201144.4]
  assign OptimizationBarrier_37_io_x_u = superpage_entries_2_data_0[14]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@201144.4]
  assign OptimizationBarrier_37_io_x_ae = superpage_entries_2_data_0[12]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@201144.4]
  assign OptimizationBarrier_37_io_x_sw = superpage_entries_2_data_0[11]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@201144.4]
  assign OptimizationBarrier_37_io_x_sx = superpage_entries_2_data_0[10]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@201144.4]
  assign OptimizationBarrier_37_io_x_sr = superpage_entries_2_data_0[9]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@201144.4]
  assign OptimizationBarrier_37_io_x_pw = superpage_entries_2_data_0[8]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@201144.4]
  assign OptimizationBarrier_37_io_x_px = superpage_entries_2_data_0[7]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@201144.4]
  assign OptimizationBarrier_37_io_x_pr = superpage_entries_2_data_0[6]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@201144.4]
  assign OptimizationBarrier_37_io_x_ppp = superpage_entries_2_data_0[5]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@201144.4]
  assign OptimizationBarrier_37_io_x_pal = superpage_entries_2_data_0[4]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@201144.4]
  assign OptimizationBarrier_37_io_x_paa = superpage_entries_2_data_0[3]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@201144.4]
  assign OptimizationBarrier_37_io_x_eff = superpage_entries_2_data_0[2]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@201144.4]
  assign OptimizationBarrier_37_io_x_c = superpage_entries_2_data_0[1]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@201144.4]
  assign OptimizationBarrier_38_io_x_ppn = superpage_entries_3_data_0[34:15]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@201186.4]
  assign OptimizationBarrier_38_io_x_u = superpage_entries_3_data_0[14]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@201186.4]
  assign OptimizationBarrier_38_io_x_ae = superpage_entries_3_data_0[12]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@201186.4]
  assign OptimizationBarrier_38_io_x_sw = superpage_entries_3_data_0[11]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@201186.4]
  assign OptimizationBarrier_38_io_x_sx = superpage_entries_3_data_0[10]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@201186.4]
  assign OptimizationBarrier_38_io_x_sr = superpage_entries_3_data_0[9]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@201186.4]
  assign OptimizationBarrier_38_io_x_pw = superpage_entries_3_data_0[8]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@201186.4]
  assign OptimizationBarrier_38_io_x_px = superpage_entries_3_data_0[7]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@201186.4]
  assign OptimizationBarrier_38_io_x_pr = superpage_entries_3_data_0[6]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@201186.4]
  assign OptimizationBarrier_38_io_x_ppp = superpage_entries_3_data_0[5]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@201186.4]
  assign OptimizationBarrier_38_io_x_pal = superpage_entries_3_data_0[4]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@201186.4]
  assign OptimizationBarrier_38_io_x_paa = superpage_entries_3_data_0[3]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@201186.4]
  assign OptimizationBarrier_38_io_x_eff = superpage_entries_3_data_0[2]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@201186.4]
  assign OptimizationBarrier_38_io_x_c = superpage_entries_3_data_0[1]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@201186.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  sectored_entries_0_tag = _RAND_0[19:0];
  _RAND_1 = {2{`RANDOM}};
  sectored_entries_0_data_0 = _RAND_1[34:0];
  _RAND_2 = {2{`RANDOM}};
  sectored_entries_0_data_1 = _RAND_2[34:0];
  _RAND_3 = {2{`RANDOM}};
  sectored_entries_0_data_2 = _RAND_3[34:0];
  _RAND_4 = {2{`RANDOM}};
  sectored_entries_0_data_3 = _RAND_4[34:0];
  _RAND_5 = {1{`RANDOM}};
  sectored_entries_0_valid_0 = _RAND_5[0:0];
  _RAND_6 = {1{`RANDOM}};
  sectored_entries_0_valid_1 = _RAND_6[0:0];
  _RAND_7 = {1{`RANDOM}};
  sectored_entries_0_valid_2 = _RAND_7[0:0];
  _RAND_8 = {1{`RANDOM}};
  sectored_entries_0_valid_3 = _RAND_8[0:0];
  _RAND_9 = {1{`RANDOM}};
  sectored_entries_1_tag = _RAND_9[19:0];
  _RAND_10 = {2{`RANDOM}};
  sectored_entries_1_data_0 = _RAND_10[34:0];
  _RAND_11 = {2{`RANDOM}};
  sectored_entries_1_data_1 = _RAND_11[34:0];
  _RAND_12 = {2{`RANDOM}};
  sectored_entries_1_data_2 = _RAND_12[34:0];
  _RAND_13 = {2{`RANDOM}};
  sectored_entries_1_data_3 = _RAND_13[34:0];
  _RAND_14 = {1{`RANDOM}};
  sectored_entries_1_valid_0 = _RAND_14[0:0];
  _RAND_15 = {1{`RANDOM}};
  sectored_entries_1_valid_1 = _RAND_15[0:0];
  _RAND_16 = {1{`RANDOM}};
  sectored_entries_1_valid_2 = _RAND_16[0:0];
  _RAND_17 = {1{`RANDOM}};
  sectored_entries_1_valid_3 = _RAND_17[0:0];
  _RAND_18 = {1{`RANDOM}};
  sectored_entries_2_tag = _RAND_18[19:0];
  _RAND_19 = {2{`RANDOM}};
  sectored_entries_2_data_0 = _RAND_19[34:0];
  _RAND_20 = {2{`RANDOM}};
  sectored_entries_2_data_1 = _RAND_20[34:0];
  _RAND_21 = {2{`RANDOM}};
  sectored_entries_2_data_2 = _RAND_21[34:0];
  _RAND_22 = {2{`RANDOM}};
  sectored_entries_2_data_3 = _RAND_22[34:0];
  _RAND_23 = {1{`RANDOM}};
  sectored_entries_2_valid_0 = _RAND_23[0:0];
  _RAND_24 = {1{`RANDOM}};
  sectored_entries_2_valid_1 = _RAND_24[0:0];
  _RAND_25 = {1{`RANDOM}};
  sectored_entries_2_valid_2 = _RAND_25[0:0];
  _RAND_26 = {1{`RANDOM}};
  sectored_entries_2_valid_3 = _RAND_26[0:0];
  _RAND_27 = {1{`RANDOM}};
  sectored_entries_3_tag = _RAND_27[19:0];
  _RAND_28 = {2{`RANDOM}};
  sectored_entries_3_data_0 = _RAND_28[34:0];
  _RAND_29 = {2{`RANDOM}};
  sectored_entries_3_data_1 = _RAND_29[34:0];
  _RAND_30 = {2{`RANDOM}};
  sectored_entries_3_data_2 = _RAND_30[34:0];
  _RAND_31 = {2{`RANDOM}};
  sectored_entries_3_data_3 = _RAND_31[34:0];
  _RAND_32 = {1{`RANDOM}};
  sectored_entries_3_valid_0 = _RAND_32[0:0];
  _RAND_33 = {1{`RANDOM}};
  sectored_entries_3_valid_1 = _RAND_33[0:0];
  _RAND_34 = {1{`RANDOM}};
  sectored_entries_3_valid_2 = _RAND_34[0:0];
  _RAND_35 = {1{`RANDOM}};
  sectored_entries_3_valid_3 = _RAND_35[0:0];
  _RAND_36 = {1{`RANDOM}};
  sectored_entries_4_tag = _RAND_36[19:0];
  _RAND_37 = {2{`RANDOM}};
  sectored_entries_4_data_0 = _RAND_37[34:0];
  _RAND_38 = {2{`RANDOM}};
  sectored_entries_4_data_1 = _RAND_38[34:0];
  _RAND_39 = {2{`RANDOM}};
  sectored_entries_4_data_2 = _RAND_39[34:0];
  _RAND_40 = {2{`RANDOM}};
  sectored_entries_4_data_3 = _RAND_40[34:0];
  _RAND_41 = {1{`RANDOM}};
  sectored_entries_4_valid_0 = _RAND_41[0:0];
  _RAND_42 = {1{`RANDOM}};
  sectored_entries_4_valid_1 = _RAND_42[0:0];
  _RAND_43 = {1{`RANDOM}};
  sectored_entries_4_valid_2 = _RAND_43[0:0];
  _RAND_44 = {1{`RANDOM}};
  sectored_entries_4_valid_3 = _RAND_44[0:0];
  _RAND_45 = {1{`RANDOM}};
  sectored_entries_5_tag = _RAND_45[19:0];
  _RAND_46 = {2{`RANDOM}};
  sectored_entries_5_data_0 = _RAND_46[34:0];
  _RAND_47 = {2{`RANDOM}};
  sectored_entries_5_data_1 = _RAND_47[34:0];
  _RAND_48 = {2{`RANDOM}};
  sectored_entries_5_data_2 = _RAND_48[34:0];
  _RAND_49 = {2{`RANDOM}};
  sectored_entries_5_data_3 = _RAND_49[34:0];
  _RAND_50 = {1{`RANDOM}};
  sectored_entries_5_valid_0 = _RAND_50[0:0];
  _RAND_51 = {1{`RANDOM}};
  sectored_entries_5_valid_1 = _RAND_51[0:0];
  _RAND_52 = {1{`RANDOM}};
  sectored_entries_5_valid_2 = _RAND_52[0:0];
  _RAND_53 = {1{`RANDOM}};
  sectored_entries_5_valid_3 = _RAND_53[0:0];
  _RAND_54 = {1{`RANDOM}};
  sectored_entries_6_tag = _RAND_54[19:0];
  _RAND_55 = {2{`RANDOM}};
  sectored_entries_6_data_0 = _RAND_55[34:0];
  _RAND_56 = {2{`RANDOM}};
  sectored_entries_6_data_1 = _RAND_56[34:0];
  _RAND_57 = {2{`RANDOM}};
  sectored_entries_6_data_2 = _RAND_57[34:0];
  _RAND_58 = {2{`RANDOM}};
  sectored_entries_6_data_3 = _RAND_58[34:0];
  _RAND_59 = {1{`RANDOM}};
  sectored_entries_6_valid_0 = _RAND_59[0:0];
  _RAND_60 = {1{`RANDOM}};
  sectored_entries_6_valid_1 = _RAND_60[0:0];
  _RAND_61 = {1{`RANDOM}};
  sectored_entries_6_valid_2 = _RAND_61[0:0];
  _RAND_62 = {1{`RANDOM}};
  sectored_entries_6_valid_3 = _RAND_62[0:0];
  _RAND_63 = {1{`RANDOM}};
  sectored_entries_7_tag = _RAND_63[19:0];
  _RAND_64 = {2{`RANDOM}};
  sectored_entries_7_data_0 = _RAND_64[34:0];
  _RAND_65 = {2{`RANDOM}};
  sectored_entries_7_data_1 = _RAND_65[34:0];
  _RAND_66 = {2{`RANDOM}};
  sectored_entries_7_data_2 = _RAND_66[34:0];
  _RAND_67 = {2{`RANDOM}};
  sectored_entries_7_data_3 = _RAND_67[34:0];
  _RAND_68 = {1{`RANDOM}};
  sectored_entries_7_valid_0 = _RAND_68[0:0];
  _RAND_69 = {1{`RANDOM}};
  sectored_entries_7_valid_1 = _RAND_69[0:0];
  _RAND_70 = {1{`RANDOM}};
  sectored_entries_7_valid_2 = _RAND_70[0:0];
  _RAND_71 = {1{`RANDOM}};
  sectored_entries_7_valid_3 = _RAND_71[0:0];
  _RAND_72 = {1{`RANDOM}};
  superpage_entries_0_tag = _RAND_72[19:0];
  _RAND_73 = {2{`RANDOM}};
  superpage_entries_0_data_0 = _RAND_73[34:0];
  _RAND_74 = {1{`RANDOM}};
  superpage_entries_0_valid_0 = _RAND_74[0:0];
  _RAND_75 = {1{`RANDOM}};
  superpage_entries_1_tag = _RAND_75[19:0];
  _RAND_76 = {2{`RANDOM}};
  superpage_entries_1_data_0 = _RAND_76[34:0];
  _RAND_77 = {1{`RANDOM}};
  superpage_entries_1_valid_0 = _RAND_77[0:0];
  _RAND_78 = {1{`RANDOM}};
  superpage_entries_2_tag = _RAND_78[19:0];
  _RAND_79 = {2{`RANDOM}};
  superpage_entries_2_data_0 = _RAND_79[34:0];
  _RAND_80 = {1{`RANDOM}};
  superpage_entries_2_valid_0 = _RAND_80[0:0];
  _RAND_81 = {1{`RANDOM}};
  superpage_entries_3_tag = _RAND_81[19:0];
  _RAND_82 = {2{`RANDOM}};
  superpage_entries_3_data_0 = _RAND_82[34:0];
  _RAND_83 = {1{`RANDOM}};
  superpage_entries_3_valid_0 = _RAND_83[0:0];
  _RAND_84 = {1{`RANDOM}};
  special_entry_level = _RAND_84[0:0];
  _RAND_85 = {1{`RANDOM}};
  special_entry_tag = _RAND_85[19:0];
  _RAND_86 = {2{`RANDOM}};
  special_entry_data_0 = _RAND_86[34:0];
  _RAND_87 = {1{`RANDOM}};
  special_entry_valid_0 = _RAND_87[0:0];
  _RAND_88 = {1{`RANDOM}};
  state = _RAND_88[1:0];
  _RAND_89 = {1{`RANDOM}};
  r_refill_tag = _RAND_89[19:0];
  _RAND_90 = {1{`RANDOM}};
  r_superpage_repl_addr = _RAND_90[1:0];
  _RAND_91 = {1{`RANDOM}};
  r_sectored_repl_addr = _RAND_91[2:0];
  _RAND_92 = {1{`RANDOM}};
  r_sectored_hit_addr = _RAND_92[2:0];
  _RAND_93 = {1{`RANDOM}};
  r_sectored_hit = _RAND_93[0:0];
  _RAND_94 = {1{`RANDOM}};
  _T_2007 = _RAND_94[6:0];
  _RAND_95 = {1{`RANDOM}};
  _T_2008 = _RAND_95[2:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (_T_939) begin
      if (!(_T_961)) begin
        if (!(_T_979)) begin
          if (_T_1045) begin
            sectored_entries_0_tag <= r_refill_tag;
          end
        end
      end
    end
    if (_T_939) begin
      if (!(_T_961)) begin
        if (!(_T_979)) begin
          if (_T_1045) begin
            if (2'h0 == r_refill_tag[1:0]) begin
              sectored_entries_0_data_0 <= _T_978;
            end
          end
        end
      end
    end
    if (_T_939) begin
      if (!(_T_961)) begin
        if (!(_T_979)) begin
          if (_T_1045) begin
            if (2'h1 == r_refill_tag[1:0]) begin
              sectored_entries_0_data_1 <= _T_978;
            end
          end
        end
      end
    end
    if (_T_939) begin
      if (!(_T_961)) begin
        if (!(_T_979)) begin
          if (_T_1045) begin
            if (2'h2 == r_refill_tag[1:0]) begin
              sectored_entries_0_data_2 <= _T_978;
            end
          end
        end
      end
    end
    if (_T_939) begin
      if (!(_T_961)) begin
        if (!(_T_979)) begin
          if (_T_1045) begin
            if (2'h3 == r_refill_tag[1:0]) begin
              sectored_entries_0_data_3 <= _T_978;
            end
          end
        end
      end
    end
    if (_T_3753) begin
      sectored_entries_0_valid_0 <= 1'h0;
    end else if (io_sfence_valid) begin
      if (io_sfence_bits_rs1) begin
        if (_T_2353) begin
          if (sectored_entries_0_data_0[0]) begin
            sectored_entries_0_valid_0 <= 1'h0;
          end else if (_T_415) begin
            if (2'h0 == vpn[1:0]) begin
              sectored_entries_0_valid_0 <= 1'h0;
            end else if (_T_939) begin
              if (!(_T_961)) begin
                if (!(_T_979)) begin
                  if (_T_1045) begin
                    sectored_entries_0_valid_0 <= _GEN_84;
                  end
                end
              end
            end
          end else if (_T_939) begin
            if (!(_T_961)) begin
              if (!(_T_979)) begin
                if (_T_1045) begin
                  sectored_entries_0_valid_0 <= _GEN_84;
                end
              end
            end
          end
        end else if (_T_415) begin
          if (2'h0 == vpn[1:0]) begin
            sectored_entries_0_valid_0 <= 1'h0;
          end else if (_T_939) begin
            if (!(_T_961)) begin
              if (!(_T_979)) begin
                if (_T_1045) begin
                  sectored_entries_0_valid_0 <= _GEN_84;
                end
              end
            end
          end
        end else if (_T_939) begin
          if (!(_T_961)) begin
            if (!(_T_979)) begin
              if (_T_1045) begin
                sectored_entries_0_valid_0 <= _GEN_84;
              end
            end
          end
        end
      end else begin
        sectored_entries_0_valid_0 <= _GEN_652;
      end
    end else begin
      sectored_entries_0_valid_0 <= _GEN_472;
    end
    if (_T_3753) begin
      sectored_entries_0_valid_1 <= 1'h0;
    end else if (io_sfence_valid) begin
      if (io_sfence_bits_rs1) begin
        if (_T_2353) begin
          if (sectored_entries_0_data_1[0]) begin
            sectored_entries_0_valid_1 <= 1'h0;
          end else if (_T_415) begin
            if (2'h1 == vpn[1:0]) begin
              sectored_entries_0_valid_1 <= 1'h0;
            end else if (_T_939) begin
              if (!(_T_961)) begin
                if (!(_T_979)) begin
                  if (_T_1045) begin
                    sectored_entries_0_valid_1 <= _GEN_85;
                  end
                end
              end
            end
          end else if (_T_939) begin
            if (!(_T_961)) begin
              if (!(_T_979)) begin
                if (_T_1045) begin
                  sectored_entries_0_valid_1 <= _GEN_85;
                end
              end
            end
          end
        end else if (_T_415) begin
          if (2'h1 == vpn[1:0]) begin
            sectored_entries_0_valid_1 <= 1'h0;
          end else if (_T_939) begin
            if (!(_T_961)) begin
              if (!(_T_979)) begin
                if (_T_1045) begin
                  sectored_entries_0_valid_1 <= _GEN_85;
                end
              end
            end
          end
        end else if (_T_939) begin
          if (!(_T_961)) begin
            if (!(_T_979)) begin
              if (_T_1045) begin
                sectored_entries_0_valid_1 <= _GEN_85;
              end
            end
          end
        end
      end else begin
        sectored_entries_0_valid_1 <= _GEN_653;
      end
    end else begin
      sectored_entries_0_valid_1 <= _GEN_473;
    end
    if (_T_3753) begin
      sectored_entries_0_valid_2 <= 1'h0;
    end else if (io_sfence_valid) begin
      if (io_sfence_bits_rs1) begin
        if (_T_2353) begin
          if (sectored_entries_0_data_2[0]) begin
            sectored_entries_0_valid_2 <= 1'h0;
          end else if (_T_415) begin
            if (2'h2 == vpn[1:0]) begin
              sectored_entries_0_valid_2 <= 1'h0;
            end else if (_T_939) begin
              if (!(_T_961)) begin
                if (!(_T_979)) begin
                  if (_T_1045) begin
                    sectored_entries_0_valid_2 <= _GEN_86;
                  end
                end
              end
            end
          end else if (_T_939) begin
            if (!(_T_961)) begin
              if (!(_T_979)) begin
                if (_T_1045) begin
                  sectored_entries_0_valid_2 <= _GEN_86;
                end
              end
            end
          end
        end else if (_T_415) begin
          if (2'h2 == vpn[1:0]) begin
            sectored_entries_0_valid_2 <= 1'h0;
          end else if (_T_939) begin
            if (!(_T_961)) begin
              if (!(_T_979)) begin
                if (_T_1045) begin
                  sectored_entries_0_valid_2 <= _GEN_86;
                end
              end
            end
          end
        end else if (_T_939) begin
          if (!(_T_961)) begin
            if (!(_T_979)) begin
              if (_T_1045) begin
                sectored_entries_0_valid_2 <= _GEN_86;
              end
            end
          end
        end
      end else begin
        sectored_entries_0_valid_2 <= _GEN_654;
      end
    end else begin
      sectored_entries_0_valid_2 <= _GEN_474;
    end
    if (_T_3753) begin
      sectored_entries_0_valid_3 <= 1'h0;
    end else if (io_sfence_valid) begin
      if (io_sfence_bits_rs1) begin
        if (_T_2353) begin
          if (sectored_entries_0_data_3[0]) begin
            sectored_entries_0_valid_3 <= 1'h0;
          end else if (_T_415) begin
            if (2'h3 == vpn[1:0]) begin
              sectored_entries_0_valid_3 <= 1'h0;
            end else if (_T_939) begin
              if (!(_T_961)) begin
                if (!(_T_979)) begin
                  if (_T_1045) begin
                    sectored_entries_0_valid_3 <= _GEN_87;
                  end
                end
              end
            end
          end else if (_T_939) begin
            if (!(_T_961)) begin
              if (!(_T_979)) begin
                if (_T_1045) begin
                  sectored_entries_0_valid_3 <= _GEN_87;
                end
              end
            end
          end
        end else if (_T_415) begin
          if (2'h3 == vpn[1:0]) begin
            sectored_entries_0_valid_3 <= 1'h0;
          end else if (_T_939) begin
            if (!(_T_961)) begin
              if (!(_T_979)) begin
                if (_T_1045) begin
                  sectored_entries_0_valid_3 <= _GEN_87;
                end
              end
            end
          end
        end else if (_T_939) begin
          if (!(_T_961)) begin
            if (!(_T_979)) begin
              if (_T_1045) begin
                sectored_entries_0_valid_3 <= _GEN_87;
              end
            end
          end
        end
      end else begin
        sectored_entries_0_valid_3 <= _GEN_655;
      end
    end else begin
      sectored_entries_0_valid_3 <= _GEN_475;
    end
    if (_T_939) begin
      if (!(_T_961)) begin
        if (!(_T_979)) begin
          if (_T_1063) begin
            sectored_entries_1_tag <= r_refill_tag;
          end
        end
      end
    end
    if (_T_939) begin
      if (!(_T_961)) begin
        if (!(_T_979)) begin
          if (_T_1063) begin
            if (2'h0 == r_refill_tag[1:0]) begin
              sectored_entries_1_data_0 <= _T_978;
            end
          end
        end
      end
    end
    if (_T_939) begin
      if (!(_T_961)) begin
        if (!(_T_979)) begin
          if (_T_1063) begin
            if (2'h1 == r_refill_tag[1:0]) begin
              sectored_entries_1_data_1 <= _T_978;
            end
          end
        end
      end
    end
    if (_T_939) begin
      if (!(_T_961)) begin
        if (!(_T_979)) begin
          if (_T_1063) begin
            if (2'h2 == r_refill_tag[1:0]) begin
              sectored_entries_1_data_2 <= _T_978;
            end
          end
        end
      end
    end
    if (_T_939) begin
      if (!(_T_961)) begin
        if (!(_T_979)) begin
          if (_T_1063) begin
            if (2'h3 == r_refill_tag[1:0]) begin
              sectored_entries_1_data_3 <= _T_978;
            end
          end
        end
      end
    end
    if (_T_3753) begin
      sectored_entries_1_valid_0 <= 1'h0;
    end else if (io_sfence_valid) begin
      if (io_sfence_bits_rs1) begin
        if (_T_2508) begin
          if (sectored_entries_1_data_0[0]) begin
            sectored_entries_1_valid_0 <= 1'h0;
          end else if (_T_421) begin
            if (2'h0 == vpn[1:0]) begin
              sectored_entries_1_valid_0 <= 1'h0;
            end else if (_T_939) begin
              if (!(_T_961)) begin
                if (!(_T_979)) begin
                  if (_T_1063) begin
                    sectored_entries_1_valid_0 <= _GEN_106;
                  end
                end
              end
            end
          end else if (_T_939) begin
            if (!(_T_961)) begin
              if (!(_T_979)) begin
                if (_T_1063) begin
                  sectored_entries_1_valid_0 <= _GEN_106;
                end
              end
            end
          end
        end else if (_T_421) begin
          if (2'h0 == vpn[1:0]) begin
            sectored_entries_1_valid_0 <= 1'h0;
          end else if (_T_939) begin
            if (!(_T_961)) begin
              if (!(_T_979)) begin
                if (_T_1063) begin
                  sectored_entries_1_valid_0 <= _GEN_106;
                end
              end
            end
          end
        end else if (_T_939) begin
          if (!(_T_961)) begin
            if (!(_T_979)) begin
              if (_T_1063) begin
                sectored_entries_1_valid_0 <= _GEN_106;
              end
            end
          end
        end
      end else begin
        sectored_entries_1_valid_0 <= _GEN_680;
      end
    end else begin
      sectored_entries_1_valid_0 <= _GEN_482;
    end
    if (_T_3753) begin
      sectored_entries_1_valid_1 <= 1'h0;
    end else if (io_sfence_valid) begin
      if (io_sfence_bits_rs1) begin
        if (_T_2508) begin
          if (sectored_entries_1_data_1[0]) begin
            sectored_entries_1_valid_1 <= 1'h0;
          end else if (_T_421) begin
            if (2'h1 == vpn[1:0]) begin
              sectored_entries_1_valid_1 <= 1'h0;
            end else if (_T_939) begin
              if (!(_T_961)) begin
                if (!(_T_979)) begin
                  if (_T_1063) begin
                    sectored_entries_1_valid_1 <= _GEN_107;
                  end
                end
              end
            end
          end else if (_T_939) begin
            if (!(_T_961)) begin
              if (!(_T_979)) begin
                if (_T_1063) begin
                  sectored_entries_1_valid_1 <= _GEN_107;
                end
              end
            end
          end
        end else if (_T_421) begin
          if (2'h1 == vpn[1:0]) begin
            sectored_entries_1_valid_1 <= 1'h0;
          end else if (_T_939) begin
            if (!(_T_961)) begin
              if (!(_T_979)) begin
                if (_T_1063) begin
                  sectored_entries_1_valid_1 <= _GEN_107;
                end
              end
            end
          end
        end else if (_T_939) begin
          if (!(_T_961)) begin
            if (!(_T_979)) begin
              if (_T_1063) begin
                sectored_entries_1_valid_1 <= _GEN_107;
              end
            end
          end
        end
      end else begin
        sectored_entries_1_valid_1 <= _GEN_681;
      end
    end else begin
      sectored_entries_1_valid_1 <= _GEN_483;
    end
    if (_T_3753) begin
      sectored_entries_1_valid_2 <= 1'h0;
    end else if (io_sfence_valid) begin
      if (io_sfence_bits_rs1) begin
        if (_T_2508) begin
          if (sectored_entries_1_data_2[0]) begin
            sectored_entries_1_valid_2 <= 1'h0;
          end else if (_T_421) begin
            if (2'h2 == vpn[1:0]) begin
              sectored_entries_1_valid_2 <= 1'h0;
            end else if (_T_939) begin
              if (!(_T_961)) begin
                if (!(_T_979)) begin
                  if (_T_1063) begin
                    sectored_entries_1_valid_2 <= _GEN_108;
                  end
                end
              end
            end
          end else if (_T_939) begin
            if (!(_T_961)) begin
              if (!(_T_979)) begin
                if (_T_1063) begin
                  sectored_entries_1_valid_2 <= _GEN_108;
                end
              end
            end
          end
        end else if (_T_421) begin
          if (2'h2 == vpn[1:0]) begin
            sectored_entries_1_valid_2 <= 1'h0;
          end else if (_T_939) begin
            if (!(_T_961)) begin
              if (!(_T_979)) begin
                if (_T_1063) begin
                  sectored_entries_1_valid_2 <= _GEN_108;
                end
              end
            end
          end
        end else if (_T_939) begin
          if (!(_T_961)) begin
            if (!(_T_979)) begin
              if (_T_1063) begin
                sectored_entries_1_valid_2 <= _GEN_108;
              end
            end
          end
        end
      end else begin
        sectored_entries_1_valid_2 <= _GEN_682;
      end
    end else begin
      sectored_entries_1_valid_2 <= _GEN_484;
    end
    if (_T_3753) begin
      sectored_entries_1_valid_3 <= 1'h0;
    end else if (io_sfence_valid) begin
      if (io_sfence_bits_rs1) begin
        if (_T_2508) begin
          if (sectored_entries_1_data_3[0]) begin
            sectored_entries_1_valid_3 <= 1'h0;
          end else if (_T_421) begin
            if (2'h3 == vpn[1:0]) begin
              sectored_entries_1_valid_3 <= 1'h0;
            end else if (_T_939) begin
              if (!(_T_961)) begin
                if (!(_T_979)) begin
                  if (_T_1063) begin
                    sectored_entries_1_valid_3 <= _GEN_109;
                  end
                end
              end
            end
          end else if (_T_939) begin
            if (!(_T_961)) begin
              if (!(_T_979)) begin
                if (_T_1063) begin
                  sectored_entries_1_valid_3 <= _GEN_109;
                end
              end
            end
          end
        end else if (_T_421) begin
          if (2'h3 == vpn[1:0]) begin
            sectored_entries_1_valid_3 <= 1'h0;
          end else if (_T_939) begin
            if (!(_T_961)) begin
              if (!(_T_979)) begin
                if (_T_1063) begin
                  sectored_entries_1_valid_3 <= _GEN_109;
                end
              end
            end
          end
        end else if (_T_939) begin
          if (!(_T_961)) begin
            if (!(_T_979)) begin
              if (_T_1063) begin
                sectored_entries_1_valid_3 <= _GEN_109;
              end
            end
          end
        end
      end else begin
        sectored_entries_1_valid_3 <= _GEN_683;
      end
    end else begin
      sectored_entries_1_valid_3 <= _GEN_485;
    end
    if (_T_939) begin
      if (!(_T_961)) begin
        if (!(_T_979)) begin
          if (_T_1081) begin
            sectored_entries_2_tag <= r_refill_tag;
          end
        end
      end
    end
    if (_T_939) begin
      if (!(_T_961)) begin
        if (!(_T_979)) begin
          if (_T_1081) begin
            if (2'h0 == r_refill_tag[1:0]) begin
              sectored_entries_2_data_0 <= _T_978;
            end
          end
        end
      end
    end
    if (_T_939) begin
      if (!(_T_961)) begin
        if (!(_T_979)) begin
          if (_T_1081) begin
            if (2'h1 == r_refill_tag[1:0]) begin
              sectored_entries_2_data_1 <= _T_978;
            end
          end
        end
      end
    end
    if (_T_939) begin
      if (!(_T_961)) begin
        if (!(_T_979)) begin
          if (_T_1081) begin
            if (2'h2 == r_refill_tag[1:0]) begin
              sectored_entries_2_data_2 <= _T_978;
            end
          end
        end
      end
    end
    if (_T_939) begin
      if (!(_T_961)) begin
        if (!(_T_979)) begin
          if (_T_1081) begin
            if (2'h3 == r_refill_tag[1:0]) begin
              sectored_entries_2_data_3 <= _T_978;
            end
          end
        end
      end
    end
    if (_T_3753) begin
      sectored_entries_2_valid_0 <= 1'h0;
    end else if (io_sfence_valid) begin
      if (io_sfence_bits_rs1) begin
        if (_T_2663) begin
          if (sectored_entries_2_data_0[0]) begin
            sectored_entries_2_valid_0 <= 1'h0;
          end else if (_T_427) begin
            if (2'h0 == vpn[1:0]) begin
              sectored_entries_2_valid_0 <= 1'h0;
            end else if (_T_939) begin
              if (!(_T_961)) begin
                if (!(_T_979)) begin
                  if (_T_1081) begin
                    sectored_entries_2_valid_0 <= _GEN_128;
                  end
                end
              end
            end
          end else if (_T_939) begin
            if (!(_T_961)) begin
              if (!(_T_979)) begin
                if (_T_1081) begin
                  sectored_entries_2_valid_0 <= _GEN_128;
                end
              end
            end
          end
        end else if (_T_427) begin
          if (2'h0 == vpn[1:0]) begin
            sectored_entries_2_valid_0 <= 1'h0;
          end else if (_T_939) begin
            if (!(_T_961)) begin
              if (!(_T_979)) begin
                if (_T_1081) begin
                  sectored_entries_2_valid_0 <= _GEN_128;
                end
              end
            end
          end
        end else if (_T_939) begin
          if (!(_T_961)) begin
            if (!(_T_979)) begin
              if (_T_1081) begin
                sectored_entries_2_valid_0 <= _GEN_128;
              end
            end
          end
        end
      end else begin
        sectored_entries_2_valid_0 <= _GEN_708;
      end
    end else begin
      sectored_entries_2_valid_0 <= _GEN_492;
    end
    if (_T_3753) begin
      sectored_entries_2_valid_1 <= 1'h0;
    end else if (io_sfence_valid) begin
      if (io_sfence_bits_rs1) begin
        if (_T_2663) begin
          if (sectored_entries_2_data_1[0]) begin
            sectored_entries_2_valid_1 <= 1'h0;
          end else if (_T_427) begin
            if (2'h1 == vpn[1:0]) begin
              sectored_entries_2_valid_1 <= 1'h0;
            end else if (_T_939) begin
              if (!(_T_961)) begin
                if (!(_T_979)) begin
                  if (_T_1081) begin
                    sectored_entries_2_valid_1 <= _GEN_129;
                  end
                end
              end
            end
          end else if (_T_939) begin
            if (!(_T_961)) begin
              if (!(_T_979)) begin
                if (_T_1081) begin
                  sectored_entries_2_valid_1 <= _GEN_129;
                end
              end
            end
          end
        end else if (_T_427) begin
          if (2'h1 == vpn[1:0]) begin
            sectored_entries_2_valid_1 <= 1'h0;
          end else if (_T_939) begin
            if (!(_T_961)) begin
              if (!(_T_979)) begin
                if (_T_1081) begin
                  sectored_entries_2_valid_1 <= _GEN_129;
                end
              end
            end
          end
        end else if (_T_939) begin
          if (!(_T_961)) begin
            if (!(_T_979)) begin
              if (_T_1081) begin
                sectored_entries_2_valid_1 <= _GEN_129;
              end
            end
          end
        end
      end else begin
        sectored_entries_2_valid_1 <= _GEN_709;
      end
    end else begin
      sectored_entries_2_valid_1 <= _GEN_493;
    end
    if (_T_3753) begin
      sectored_entries_2_valid_2 <= 1'h0;
    end else if (io_sfence_valid) begin
      if (io_sfence_bits_rs1) begin
        if (_T_2663) begin
          if (sectored_entries_2_data_2[0]) begin
            sectored_entries_2_valid_2 <= 1'h0;
          end else if (_T_427) begin
            if (2'h2 == vpn[1:0]) begin
              sectored_entries_2_valid_2 <= 1'h0;
            end else if (_T_939) begin
              if (!(_T_961)) begin
                if (!(_T_979)) begin
                  if (_T_1081) begin
                    sectored_entries_2_valid_2 <= _GEN_130;
                  end
                end
              end
            end
          end else if (_T_939) begin
            if (!(_T_961)) begin
              if (!(_T_979)) begin
                if (_T_1081) begin
                  sectored_entries_2_valid_2 <= _GEN_130;
                end
              end
            end
          end
        end else if (_T_427) begin
          if (2'h2 == vpn[1:0]) begin
            sectored_entries_2_valid_2 <= 1'h0;
          end else if (_T_939) begin
            if (!(_T_961)) begin
              if (!(_T_979)) begin
                if (_T_1081) begin
                  sectored_entries_2_valid_2 <= _GEN_130;
                end
              end
            end
          end
        end else if (_T_939) begin
          if (!(_T_961)) begin
            if (!(_T_979)) begin
              if (_T_1081) begin
                sectored_entries_2_valid_2 <= _GEN_130;
              end
            end
          end
        end
      end else begin
        sectored_entries_2_valid_2 <= _GEN_710;
      end
    end else begin
      sectored_entries_2_valid_2 <= _GEN_494;
    end
    if (_T_3753) begin
      sectored_entries_2_valid_3 <= 1'h0;
    end else if (io_sfence_valid) begin
      if (io_sfence_bits_rs1) begin
        if (_T_2663) begin
          if (sectored_entries_2_data_3[0]) begin
            sectored_entries_2_valid_3 <= 1'h0;
          end else if (_T_427) begin
            if (2'h3 == vpn[1:0]) begin
              sectored_entries_2_valid_3 <= 1'h0;
            end else if (_T_939) begin
              if (!(_T_961)) begin
                if (!(_T_979)) begin
                  if (_T_1081) begin
                    sectored_entries_2_valid_3 <= _GEN_131;
                  end
                end
              end
            end
          end else if (_T_939) begin
            if (!(_T_961)) begin
              if (!(_T_979)) begin
                if (_T_1081) begin
                  sectored_entries_2_valid_3 <= _GEN_131;
                end
              end
            end
          end
        end else if (_T_427) begin
          if (2'h3 == vpn[1:0]) begin
            sectored_entries_2_valid_3 <= 1'h0;
          end else if (_T_939) begin
            if (!(_T_961)) begin
              if (!(_T_979)) begin
                if (_T_1081) begin
                  sectored_entries_2_valid_3 <= _GEN_131;
                end
              end
            end
          end
        end else if (_T_939) begin
          if (!(_T_961)) begin
            if (!(_T_979)) begin
              if (_T_1081) begin
                sectored_entries_2_valid_3 <= _GEN_131;
              end
            end
          end
        end
      end else begin
        sectored_entries_2_valid_3 <= _GEN_711;
      end
    end else begin
      sectored_entries_2_valid_3 <= _GEN_495;
    end
    if (_T_939) begin
      if (!(_T_961)) begin
        if (!(_T_979)) begin
          if (_T_1099) begin
            sectored_entries_3_tag <= r_refill_tag;
          end
        end
      end
    end
    if (_T_939) begin
      if (!(_T_961)) begin
        if (!(_T_979)) begin
          if (_T_1099) begin
            if (2'h0 == r_refill_tag[1:0]) begin
              sectored_entries_3_data_0 <= _T_978;
            end
          end
        end
      end
    end
    if (_T_939) begin
      if (!(_T_961)) begin
        if (!(_T_979)) begin
          if (_T_1099) begin
            if (2'h1 == r_refill_tag[1:0]) begin
              sectored_entries_3_data_1 <= _T_978;
            end
          end
        end
      end
    end
    if (_T_939) begin
      if (!(_T_961)) begin
        if (!(_T_979)) begin
          if (_T_1099) begin
            if (2'h2 == r_refill_tag[1:0]) begin
              sectored_entries_3_data_2 <= _T_978;
            end
          end
        end
      end
    end
    if (_T_939) begin
      if (!(_T_961)) begin
        if (!(_T_979)) begin
          if (_T_1099) begin
            if (2'h3 == r_refill_tag[1:0]) begin
              sectored_entries_3_data_3 <= _T_978;
            end
          end
        end
      end
    end
    if (_T_3753) begin
      sectored_entries_3_valid_0 <= 1'h0;
    end else if (io_sfence_valid) begin
      if (io_sfence_bits_rs1) begin
        if (_T_2818) begin
          if (sectored_entries_3_data_0[0]) begin
            sectored_entries_3_valid_0 <= 1'h0;
          end else if (_T_433) begin
            if (2'h0 == vpn[1:0]) begin
              sectored_entries_3_valid_0 <= 1'h0;
            end else if (_T_939) begin
              if (!(_T_961)) begin
                if (!(_T_979)) begin
                  if (_T_1099) begin
                    sectored_entries_3_valid_0 <= _GEN_150;
                  end
                end
              end
            end
          end else if (_T_939) begin
            if (!(_T_961)) begin
              if (!(_T_979)) begin
                if (_T_1099) begin
                  sectored_entries_3_valid_0 <= _GEN_150;
                end
              end
            end
          end
        end else if (_T_433) begin
          if (2'h0 == vpn[1:0]) begin
            sectored_entries_3_valid_0 <= 1'h0;
          end else if (_T_939) begin
            if (!(_T_961)) begin
              if (!(_T_979)) begin
                if (_T_1099) begin
                  sectored_entries_3_valid_0 <= _GEN_150;
                end
              end
            end
          end
        end else if (_T_939) begin
          if (!(_T_961)) begin
            if (!(_T_979)) begin
              if (_T_1099) begin
                sectored_entries_3_valid_0 <= _GEN_150;
              end
            end
          end
        end
      end else begin
        sectored_entries_3_valid_0 <= _GEN_736;
      end
    end else begin
      sectored_entries_3_valid_0 <= _GEN_502;
    end
    if (_T_3753) begin
      sectored_entries_3_valid_1 <= 1'h0;
    end else if (io_sfence_valid) begin
      if (io_sfence_bits_rs1) begin
        if (_T_2818) begin
          if (sectored_entries_3_data_1[0]) begin
            sectored_entries_3_valid_1 <= 1'h0;
          end else if (_T_433) begin
            if (2'h1 == vpn[1:0]) begin
              sectored_entries_3_valid_1 <= 1'h0;
            end else if (_T_939) begin
              if (!(_T_961)) begin
                if (!(_T_979)) begin
                  if (_T_1099) begin
                    sectored_entries_3_valid_1 <= _GEN_151;
                  end
                end
              end
            end
          end else if (_T_939) begin
            if (!(_T_961)) begin
              if (!(_T_979)) begin
                if (_T_1099) begin
                  sectored_entries_3_valid_1 <= _GEN_151;
                end
              end
            end
          end
        end else if (_T_433) begin
          if (2'h1 == vpn[1:0]) begin
            sectored_entries_3_valid_1 <= 1'h0;
          end else if (_T_939) begin
            if (!(_T_961)) begin
              if (!(_T_979)) begin
                if (_T_1099) begin
                  sectored_entries_3_valid_1 <= _GEN_151;
                end
              end
            end
          end
        end else if (_T_939) begin
          if (!(_T_961)) begin
            if (!(_T_979)) begin
              if (_T_1099) begin
                sectored_entries_3_valid_1 <= _GEN_151;
              end
            end
          end
        end
      end else begin
        sectored_entries_3_valid_1 <= _GEN_737;
      end
    end else begin
      sectored_entries_3_valid_1 <= _GEN_503;
    end
    if (_T_3753) begin
      sectored_entries_3_valid_2 <= 1'h0;
    end else if (io_sfence_valid) begin
      if (io_sfence_bits_rs1) begin
        if (_T_2818) begin
          if (sectored_entries_3_data_2[0]) begin
            sectored_entries_3_valid_2 <= 1'h0;
          end else if (_T_433) begin
            if (2'h2 == vpn[1:0]) begin
              sectored_entries_3_valid_2 <= 1'h0;
            end else if (_T_939) begin
              if (!(_T_961)) begin
                if (!(_T_979)) begin
                  if (_T_1099) begin
                    sectored_entries_3_valid_2 <= _GEN_152;
                  end
                end
              end
            end
          end else if (_T_939) begin
            if (!(_T_961)) begin
              if (!(_T_979)) begin
                if (_T_1099) begin
                  sectored_entries_3_valid_2 <= _GEN_152;
                end
              end
            end
          end
        end else if (_T_433) begin
          if (2'h2 == vpn[1:0]) begin
            sectored_entries_3_valid_2 <= 1'h0;
          end else if (_T_939) begin
            if (!(_T_961)) begin
              if (!(_T_979)) begin
                if (_T_1099) begin
                  sectored_entries_3_valid_2 <= _GEN_152;
                end
              end
            end
          end
        end else if (_T_939) begin
          if (!(_T_961)) begin
            if (!(_T_979)) begin
              if (_T_1099) begin
                sectored_entries_3_valid_2 <= _GEN_152;
              end
            end
          end
        end
      end else begin
        sectored_entries_3_valid_2 <= _GEN_738;
      end
    end else begin
      sectored_entries_3_valid_2 <= _GEN_504;
    end
    if (_T_3753) begin
      sectored_entries_3_valid_3 <= 1'h0;
    end else if (io_sfence_valid) begin
      if (io_sfence_bits_rs1) begin
        if (_T_2818) begin
          if (sectored_entries_3_data_3[0]) begin
            sectored_entries_3_valid_3 <= 1'h0;
          end else if (_T_433) begin
            if (2'h3 == vpn[1:0]) begin
              sectored_entries_3_valid_3 <= 1'h0;
            end else if (_T_939) begin
              if (!(_T_961)) begin
                if (!(_T_979)) begin
                  if (_T_1099) begin
                    sectored_entries_3_valid_3 <= _GEN_153;
                  end
                end
              end
            end
          end else if (_T_939) begin
            if (!(_T_961)) begin
              if (!(_T_979)) begin
                if (_T_1099) begin
                  sectored_entries_3_valid_3 <= _GEN_153;
                end
              end
            end
          end
        end else if (_T_433) begin
          if (2'h3 == vpn[1:0]) begin
            sectored_entries_3_valid_3 <= 1'h0;
          end else if (_T_939) begin
            if (!(_T_961)) begin
              if (!(_T_979)) begin
                if (_T_1099) begin
                  sectored_entries_3_valid_3 <= _GEN_153;
                end
              end
            end
          end
        end else if (_T_939) begin
          if (!(_T_961)) begin
            if (!(_T_979)) begin
              if (_T_1099) begin
                sectored_entries_3_valid_3 <= _GEN_153;
              end
            end
          end
        end
      end else begin
        sectored_entries_3_valid_3 <= _GEN_739;
      end
    end else begin
      sectored_entries_3_valid_3 <= _GEN_505;
    end
    if (_T_939) begin
      if (!(_T_961)) begin
        if (!(_T_979)) begin
          if (_T_1117) begin
            sectored_entries_4_tag <= r_refill_tag;
          end
        end
      end
    end
    if (_T_939) begin
      if (!(_T_961)) begin
        if (!(_T_979)) begin
          if (_T_1117) begin
            if (2'h0 == r_refill_tag[1:0]) begin
              sectored_entries_4_data_0 <= _T_978;
            end
          end
        end
      end
    end
    if (_T_939) begin
      if (!(_T_961)) begin
        if (!(_T_979)) begin
          if (_T_1117) begin
            if (2'h1 == r_refill_tag[1:0]) begin
              sectored_entries_4_data_1 <= _T_978;
            end
          end
        end
      end
    end
    if (_T_939) begin
      if (!(_T_961)) begin
        if (!(_T_979)) begin
          if (_T_1117) begin
            if (2'h2 == r_refill_tag[1:0]) begin
              sectored_entries_4_data_2 <= _T_978;
            end
          end
        end
      end
    end
    if (_T_939) begin
      if (!(_T_961)) begin
        if (!(_T_979)) begin
          if (_T_1117) begin
            if (2'h3 == r_refill_tag[1:0]) begin
              sectored_entries_4_data_3 <= _T_978;
            end
          end
        end
      end
    end
    if (_T_3753) begin
      sectored_entries_4_valid_0 <= 1'h0;
    end else if (io_sfence_valid) begin
      if (io_sfence_bits_rs1) begin
        if (_T_2973) begin
          if (sectored_entries_4_data_0[0]) begin
            sectored_entries_4_valid_0 <= 1'h0;
          end else if (_T_439) begin
            if (2'h0 == vpn[1:0]) begin
              sectored_entries_4_valid_0 <= 1'h0;
            end else if (_T_939) begin
              if (!(_T_961)) begin
                if (!(_T_979)) begin
                  if (_T_1117) begin
                    sectored_entries_4_valid_0 <= _GEN_172;
                  end
                end
              end
            end
          end else if (_T_939) begin
            if (!(_T_961)) begin
              if (!(_T_979)) begin
                if (_T_1117) begin
                  sectored_entries_4_valid_0 <= _GEN_172;
                end
              end
            end
          end
        end else if (_T_439) begin
          if (2'h0 == vpn[1:0]) begin
            sectored_entries_4_valid_0 <= 1'h0;
          end else if (_T_939) begin
            if (!(_T_961)) begin
              if (!(_T_979)) begin
                if (_T_1117) begin
                  sectored_entries_4_valid_0 <= _GEN_172;
                end
              end
            end
          end
        end else if (_T_939) begin
          if (!(_T_961)) begin
            if (!(_T_979)) begin
              if (_T_1117) begin
                sectored_entries_4_valid_0 <= _GEN_172;
              end
            end
          end
        end
      end else begin
        sectored_entries_4_valid_0 <= _GEN_764;
      end
    end else begin
      sectored_entries_4_valid_0 <= _GEN_512;
    end
    if (_T_3753) begin
      sectored_entries_4_valid_1 <= 1'h0;
    end else if (io_sfence_valid) begin
      if (io_sfence_bits_rs1) begin
        if (_T_2973) begin
          if (sectored_entries_4_data_1[0]) begin
            sectored_entries_4_valid_1 <= 1'h0;
          end else if (_T_439) begin
            if (2'h1 == vpn[1:0]) begin
              sectored_entries_4_valid_1 <= 1'h0;
            end else if (_T_939) begin
              if (!(_T_961)) begin
                if (!(_T_979)) begin
                  if (_T_1117) begin
                    sectored_entries_4_valid_1 <= _GEN_173;
                  end
                end
              end
            end
          end else if (_T_939) begin
            if (!(_T_961)) begin
              if (!(_T_979)) begin
                if (_T_1117) begin
                  sectored_entries_4_valid_1 <= _GEN_173;
                end
              end
            end
          end
        end else if (_T_439) begin
          if (2'h1 == vpn[1:0]) begin
            sectored_entries_4_valid_1 <= 1'h0;
          end else if (_T_939) begin
            if (!(_T_961)) begin
              if (!(_T_979)) begin
                if (_T_1117) begin
                  sectored_entries_4_valid_1 <= _GEN_173;
                end
              end
            end
          end
        end else if (_T_939) begin
          if (!(_T_961)) begin
            if (!(_T_979)) begin
              if (_T_1117) begin
                sectored_entries_4_valid_1 <= _GEN_173;
              end
            end
          end
        end
      end else begin
        sectored_entries_4_valid_1 <= _GEN_765;
      end
    end else begin
      sectored_entries_4_valid_1 <= _GEN_513;
    end
    if (_T_3753) begin
      sectored_entries_4_valid_2 <= 1'h0;
    end else if (io_sfence_valid) begin
      if (io_sfence_bits_rs1) begin
        if (_T_2973) begin
          if (sectored_entries_4_data_2[0]) begin
            sectored_entries_4_valid_2 <= 1'h0;
          end else if (_T_439) begin
            if (2'h2 == vpn[1:0]) begin
              sectored_entries_4_valid_2 <= 1'h0;
            end else if (_T_939) begin
              if (!(_T_961)) begin
                if (!(_T_979)) begin
                  if (_T_1117) begin
                    sectored_entries_4_valid_2 <= _GEN_174;
                  end
                end
              end
            end
          end else if (_T_939) begin
            if (!(_T_961)) begin
              if (!(_T_979)) begin
                if (_T_1117) begin
                  sectored_entries_4_valid_2 <= _GEN_174;
                end
              end
            end
          end
        end else if (_T_439) begin
          if (2'h2 == vpn[1:0]) begin
            sectored_entries_4_valid_2 <= 1'h0;
          end else if (_T_939) begin
            if (!(_T_961)) begin
              if (!(_T_979)) begin
                if (_T_1117) begin
                  sectored_entries_4_valid_2 <= _GEN_174;
                end
              end
            end
          end
        end else if (_T_939) begin
          if (!(_T_961)) begin
            if (!(_T_979)) begin
              if (_T_1117) begin
                sectored_entries_4_valid_2 <= _GEN_174;
              end
            end
          end
        end
      end else begin
        sectored_entries_4_valid_2 <= _GEN_766;
      end
    end else begin
      sectored_entries_4_valid_2 <= _GEN_514;
    end
    if (_T_3753) begin
      sectored_entries_4_valid_3 <= 1'h0;
    end else if (io_sfence_valid) begin
      if (io_sfence_bits_rs1) begin
        if (_T_2973) begin
          if (sectored_entries_4_data_3[0]) begin
            sectored_entries_4_valid_3 <= 1'h0;
          end else if (_T_439) begin
            if (2'h3 == vpn[1:0]) begin
              sectored_entries_4_valid_3 <= 1'h0;
            end else if (_T_939) begin
              if (!(_T_961)) begin
                if (!(_T_979)) begin
                  if (_T_1117) begin
                    sectored_entries_4_valid_3 <= _GEN_175;
                  end
                end
              end
            end
          end else if (_T_939) begin
            if (!(_T_961)) begin
              if (!(_T_979)) begin
                if (_T_1117) begin
                  sectored_entries_4_valid_3 <= _GEN_175;
                end
              end
            end
          end
        end else if (_T_439) begin
          if (2'h3 == vpn[1:0]) begin
            sectored_entries_4_valid_3 <= 1'h0;
          end else if (_T_939) begin
            if (!(_T_961)) begin
              if (!(_T_979)) begin
                if (_T_1117) begin
                  sectored_entries_4_valid_3 <= _GEN_175;
                end
              end
            end
          end
        end else if (_T_939) begin
          if (!(_T_961)) begin
            if (!(_T_979)) begin
              if (_T_1117) begin
                sectored_entries_4_valid_3 <= _GEN_175;
              end
            end
          end
        end
      end else begin
        sectored_entries_4_valid_3 <= _GEN_767;
      end
    end else begin
      sectored_entries_4_valid_3 <= _GEN_515;
    end
    if (_T_939) begin
      if (!(_T_961)) begin
        if (!(_T_979)) begin
          if (_T_1135) begin
            sectored_entries_5_tag <= r_refill_tag;
          end
        end
      end
    end
    if (_T_939) begin
      if (!(_T_961)) begin
        if (!(_T_979)) begin
          if (_T_1135) begin
            if (2'h0 == r_refill_tag[1:0]) begin
              sectored_entries_5_data_0 <= _T_978;
            end
          end
        end
      end
    end
    if (_T_939) begin
      if (!(_T_961)) begin
        if (!(_T_979)) begin
          if (_T_1135) begin
            if (2'h1 == r_refill_tag[1:0]) begin
              sectored_entries_5_data_1 <= _T_978;
            end
          end
        end
      end
    end
    if (_T_939) begin
      if (!(_T_961)) begin
        if (!(_T_979)) begin
          if (_T_1135) begin
            if (2'h2 == r_refill_tag[1:0]) begin
              sectored_entries_5_data_2 <= _T_978;
            end
          end
        end
      end
    end
    if (_T_939) begin
      if (!(_T_961)) begin
        if (!(_T_979)) begin
          if (_T_1135) begin
            if (2'h3 == r_refill_tag[1:0]) begin
              sectored_entries_5_data_3 <= _T_978;
            end
          end
        end
      end
    end
    if (_T_3753) begin
      sectored_entries_5_valid_0 <= 1'h0;
    end else if (io_sfence_valid) begin
      if (io_sfence_bits_rs1) begin
        if (_T_3128) begin
          if (sectored_entries_5_data_0[0]) begin
            sectored_entries_5_valid_0 <= 1'h0;
          end else if (_T_445) begin
            if (2'h0 == vpn[1:0]) begin
              sectored_entries_5_valid_0 <= 1'h0;
            end else if (_T_939) begin
              if (!(_T_961)) begin
                if (!(_T_979)) begin
                  if (_T_1135) begin
                    sectored_entries_5_valid_0 <= _GEN_194;
                  end
                end
              end
            end
          end else if (_T_939) begin
            if (!(_T_961)) begin
              if (!(_T_979)) begin
                if (_T_1135) begin
                  sectored_entries_5_valid_0 <= _GEN_194;
                end
              end
            end
          end
        end else if (_T_445) begin
          if (2'h0 == vpn[1:0]) begin
            sectored_entries_5_valid_0 <= 1'h0;
          end else if (_T_939) begin
            if (!(_T_961)) begin
              if (!(_T_979)) begin
                if (_T_1135) begin
                  sectored_entries_5_valid_0 <= _GEN_194;
                end
              end
            end
          end
        end else if (_T_939) begin
          if (!(_T_961)) begin
            if (!(_T_979)) begin
              if (_T_1135) begin
                sectored_entries_5_valid_0 <= _GEN_194;
              end
            end
          end
        end
      end else begin
        sectored_entries_5_valid_0 <= _GEN_792;
      end
    end else begin
      sectored_entries_5_valid_0 <= _GEN_522;
    end
    if (_T_3753) begin
      sectored_entries_5_valid_1 <= 1'h0;
    end else if (io_sfence_valid) begin
      if (io_sfence_bits_rs1) begin
        if (_T_3128) begin
          if (sectored_entries_5_data_1[0]) begin
            sectored_entries_5_valid_1 <= 1'h0;
          end else if (_T_445) begin
            if (2'h1 == vpn[1:0]) begin
              sectored_entries_5_valid_1 <= 1'h0;
            end else if (_T_939) begin
              if (!(_T_961)) begin
                if (!(_T_979)) begin
                  if (_T_1135) begin
                    sectored_entries_5_valid_1 <= _GEN_195;
                  end
                end
              end
            end
          end else if (_T_939) begin
            if (!(_T_961)) begin
              if (!(_T_979)) begin
                if (_T_1135) begin
                  sectored_entries_5_valid_1 <= _GEN_195;
                end
              end
            end
          end
        end else if (_T_445) begin
          if (2'h1 == vpn[1:0]) begin
            sectored_entries_5_valid_1 <= 1'h0;
          end else if (_T_939) begin
            if (!(_T_961)) begin
              if (!(_T_979)) begin
                if (_T_1135) begin
                  sectored_entries_5_valid_1 <= _GEN_195;
                end
              end
            end
          end
        end else if (_T_939) begin
          if (!(_T_961)) begin
            if (!(_T_979)) begin
              if (_T_1135) begin
                sectored_entries_5_valid_1 <= _GEN_195;
              end
            end
          end
        end
      end else begin
        sectored_entries_5_valid_1 <= _GEN_793;
      end
    end else begin
      sectored_entries_5_valid_1 <= _GEN_523;
    end
    if (_T_3753) begin
      sectored_entries_5_valid_2 <= 1'h0;
    end else if (io_sfence_valid) begin
      if (io_sfence_bits_rs1) begin
        if (_T_3128) begin
          if (sectored_entries_5_data_2[0]) begin
            sectored_entries_5_valid_2 <= 1'h0;
          end else if (_T_445) begin
            if (2'h2 == vpn[1:0]) begin
              sectored_entries_5_valid_2 <= 1'h0;
            end else if (_T_939) begin
              if (!(_T_961)) begin
                if (!(_T_979)) begin
                  if (_T_1135) begin
                    sectored_entries_5_valid_2 <= _GEN_196;
                  end
                end
              end
            end
          end else if (_T_939) begin
            if (!(_T_961)) begin
              if (!(_T_979)) begin
                if (_T_1135) begin
                  sectored_entries_5_valid_2 <= _GEN_196;
                end
              end
            end
          end
        end else if (_T_445) begin
          if (2'h2 == vpn[1:0]) begin
            sectored_entries_5_valid_2 <= 1'h0;
          end else if (_T_939) begin
            if (!(_T_961)) begin
              if (!(_T_979)) begin
                if (_T_1135) begin
                  sectored_entries_5_valid_2 <= _GEN_196;
                end
              end
            end
          end
        end else if (_T_939) begin
          if (!(_T_961)) begin
            if (!(_T_979)) begin
              if (_T_1135) begin
                sectored_entries_5_valid_2 <= _GEN_196;
              end
            end
          end
        end
      end else begin
        sectored_entries_5_valid_2 <= _GEN_794;
      end
    end else begin
      sectored_entries_5_valid_2 <= _GEN_524;
    end
    if (_T_3753) begin
      sectored_entries_5_valid_3 <= 1'h0;
    end else if (io_sfence_valid) begin
      if (io_sfence_bits_rs1) begin
        if (_T_3128) begin
          if (sectored_entries_5_data_3[0]) begin
            sectored_entries_5_valid_3 <= 1'h0;
          end else if (_T_445) begin
            if (2'h3 == vpn[1:0]) begin
              sectored_entries_5_valid_3 <= 1'h0;
            end else if (_T_939) begin
              if (!(_T_961)) begin
                if (!(_T_979)) begin
                  if (_T_1135) begin
                    sectored_entries_5_valid_3 <= _GEN_197;
                  end
                end
              end
            end
          end else if (_T_939) begin
            if (!(_T_961)) begin
              if (!(_T_979)) begin
                if (_T_1135) begin
                  sectored_entries_5_valid_3 <= _GEN_197;
                end
              end
            end
          end
        end else if (_T_445) begin
          if (2'h3 == vpn[1:0]) begin
            sectored_entries_5_valid_3 <= 1'h0;
          end else if (_T_939) begin
            if (!(_T_961)) begin
              if (!(_T_979)) begin
                if (_T_1135) begin
                  sectored_entries_5_valid_3 <= _GEN_197;
                end
              end
            end
          end
        end else if (_T_939) begin
          if (!(_T_961)) begin
            if (!(_T_979)) begin
              if (_T_1135) begin
                sectored_entries_5_valid_3 <= _GEN_197;
              end
            end
          end
        end
      end else begin
        sectored_entries_5_valid_3 <= _GEN_795;
      end
    end else begin
      sectored_entries_5_valid_3 <= _GEN_525;
    end
    if (_T_939) begin
      if (!(_T_961)) begin
        if (!(_T_979)) begin
          if (_T_1153) begin
            sectored_entries_6_tag <= r_refill_tag;
          end
        end
      end
    end
    if (_T_939) begin
      if (!(_T_961)) begin
        if (!(_T_979)) begin
          if (_T_1153) begin
            if (2'h0 == r_refill_tag[1:0]) begin
              sectored_entries_6_data_0 <= _T_978;
            end
          end
        end
      end
    end
    if (_T_939) begin
      if (!(_T_961)) begin
        if (!(_T_979)) begin
          if (_T_1153) begin
            if (2'h1 == r_refill_tag[1:0]) begin
              sectored_entries_6_data_1 <= _T_978;
            end
          end
        end
      end
    end
    if (_T_939) begin
      if (!(_T_961)) begin
        if (!(_T_979)) begin
          if (_T_1153) begin
            if (2'h2 == r_refill_tag[1:0]) begin
              sectored_entries_6_data_2 <= _T_978;
            end
          end
        end
      end
    end
    if (_T_939) begin
      if (!(_T_961)) begin
        if (!(_T_979)) begin
          if (_T_1153) begin
            if (2'h3 == r_refill_tag[1:0]) begin
              sectored_entries_6_data_3 <= _T_978;
            end
          end
        end
      end
    end
    if (_T_3753) begin
      sectored_entries_6_valid_0 <= 1'h0;
    end else if (io_sfence_valid) begin
      if (io_sfence_bits_rs1) begin
        if (_T_3283) begin
          if (sectored_entries_6_data_0[0]) begin
            sectored_entries_6_valid_0 <= 1'h0;
          end else if (_T_451) begin
            if (2'h0 == vpn[1:0]) begin
              sectored_entries_6_valid_0 <= 1'h0;
            end else if (_T_939) begin
              if (!(_T_961)) begin
                if (!(_T_979)) begin
                  if (_T_1153) begin
                    sectored_entries_6_valid_0 <= _GEN_216;
                  end
                end
              end
            end
          end else if (_T_939) begin
            if (!(_T_961)) begin
              if (!(_T_979)) begin
                if (_T_1153) begin
                  sectored_entries_6_valid_0 <= _GEN_216;
                end
              end
            end
          end
        end else if (_T_451) begin
          if (2'h0 == vpn[1:0]) begin
            sectored_entries_6_valid_0 <= 1'h0;
          end else if (_T_939) begin
            if (!(_T_961)) begin
              if (!(_T_979)) begin
                if (_T_1153) begin
                  sectored_entries_6_valid_0 <= _GEN_216;
                end
              end
            end
          end
        end else if (_T_939) begin
          if (!(_T_961)) begin
            if (!(_T_979)) begin
              if (_T_1153) begin
                sectored_entries_6_valid_0 <= _GEN_216;
              end
            end
          end
        end
      end else begin
        sectored_entries_6_valid_0 <= _GEN_820;
      end
    end else begin
      sectored_entries_6_valid_0 <= _GEN_532;
    end
    if (_T_3753) begin
      sectored_entries_6_valid_1 <= 1'h0;
    end else if (io_sfence_valid) begin
      if (io_sfence_bits_rs1) begin
        if (_T_3283) begin
          if (sectored_entries_6_data_1[0]) begin
            sectored_entries_6_valid_1 <= 1'h0;
          end else if (_T_451) begin
            if (2'h1 == vpn[1:0]) begin
              sectored_entries_6_valid_1 <= 1'h0;
            end else if (_T_939) begin
              if (!(_T_961)) begin
                if (!(_T_979)) begin
                  if (_T_1153) begin
                    sectored_entries_6_valid_1 <= _GEN_217;
                  end
                end
              end
            end
          end else if (_T_939) begin
            if (!(_T_961)) begin
              if (!(_T_979)) begin
                if (_T_1153) begin
                  sectored_entries_6_valid_1 <= _GEN_217;
                end
              end
            end
          end
        end else if (_T_451) begin
          if (2'h1 == vpn[1:0]) begin
            sectored_entries_6_valid_1 <= 1'h0;
          end else if (_T_939) begin
            if (!(_T_961)) begin
              if (!(_T_979)) begin
                if (_T_1153) begin
                  sectored_entries_6_valid_1 <= _GEN_217;
                end
              end
            end
          end
        end else if (_T_939) begin
          if (!(_T_961)) begin
            if (!(_T_979)) begin
              if (_T_1153) begin
                sectored_entries_6_valid_1 <= _GEN_217;
              end
            end
          end
        end
      end else begin
        sectored_entries_6_valid_1 <= _GEN_821;
      end
    end else begin
      sectored_entries_6_valid_1 <= _GEN_533;
    end
    if (_T_3753) begin
      sectored_entries_6_valid_2 <= 1'h0;
    end else if (io_sfence_valid) begin
      if (io_sfence_bits_rs1) begin
        if (_T_3283) begin
          if (sectored_entries_6_data_2[0]) begin
            sectored_entries_6_valid_2 <= 1'h0;
          end else if (_T_451) begin
            if (2'h2 == vpn[1:0]) begin
              sectored_entries_6_valid_2 <= 1'h0;
            end else if (_T_939) begin
              if (!(_T_961)) begin
                if (!(_T_979)) begin
                  if (_T_1153) begin
                    sectored_entries_6_valid_2 <= _GEN_218;
                  end
                end
              end
            end
          end else if (_T_939) begin
            if (!(_T_961)) begin
              if (!(_T_979)) begin
                if (_T_1153) begin
                  sectored_entries_6_valid_2 <= _GEN_218;
                end
              end
            end
          end
        end else if (_T_451) begin
          if (2'h2 == vpn[1:0]) begin
            sectored_entries_6_valid_2 <= 1'h0;
          end else if (_T_939) begin
            if (!(_T_961)) begin
              if (!(_T_979)) begin
                if (_T_1153) begin
                  sectored_entries_6_valid_2 <= _GEN_218;
                end
              end
            end
          end
        end else if (_T_939) begin
          if (!(_T_961)) begin
            if (!(_T_979)) begin
              if (_T_1153) begin
                sectored_entries_6_valid_2 <= _GEN_218;
              end
            end
          end
        end
      end else begin
        sectored_entries_6_valid_2 <= _GEN_822;
      end
    end else begin
      sectored_entries_6_valid_2 <= _GEN_534;
    end
    if (_T_3753) begin
      sectored_entries_6_valid_3 <= 1'h0;
    end else if (io_sfence_valid) begin
      if (io_sfence_bits_rs1) begin
        if (_T_3283) begin
          if (sectored_entries_6_data_3[0]) begin
            sectored_entries_6_valid_3 <= 1'h0;
          end else if (_T_451) begin
            if (2'h3 == vpn[1:0]) begin
              sectored_entries_6_valid_3 <= 1'h0;
            end else if (_T_939) begin
              if (!(_T_961)) begin
                if (!(_T_979)) begin
                  if (_T_1153) begin
                    sectored_entries_6_valid_3 <= _GEN_219;
                  end
                end
              end
            end
          end else if (_T_939) begin
            if (!(_T_961)) begin
              if (!(_T_979)) begin
                if (_T_1153) begin
                  sectored_entries_6_valid_3 <= _GEN_219;
                end
              end
            end
          end
        end else if (_T_451) begin
          if (2'h3 == vpn[1:0]) begin
            sectored_entries_6_valid_3 <= 1'h0;
          end else if (_T_939) begin
            if (!(_T_961)) begin
              if (!(_T_979)) begin
                if (_T_1153) begin
                  sectored_entries_6_valid_3 <= _GEN_219;
                end
              end
            end
          end
        end else if (_T_939) begin
          if (!(_T_961)) begin
            if (!(_T_979)) begin
              if (_T_1153) begin
                sectored_entries_6_valid_3 <= _GEN_219;
              end
            end
          end
        end
      end else begin
        sectored_entries_6_valid_3 <= _GEN_823;
      end
    end else begin
      sectored_entries_6_valid_3 <= _GEN_535;
    end
    if (_T_939) begin
      if (!(_T_961)) begin
        if (!(_T_979)) begin
          if (_T_1171) begin
            sectored_entries_7_tag <= r_refill_tag;
          end
        end
      end
    end
    if (_T_939) begin
      if (!(_T_961)) begin
        if (!(_T_979)) begin
          if (_T_1171) begin
            if (2'h0 == r_refill_tag[1:0]) begin
              sectored_entries_7_data_0 <= _T_978;
            end
          end
        end
      end
    end
    if (_T_939) begin
      if (!(_T_961)) begin
        if (!(_T_979)) begin
          if (_T_1171) begin
            if (2'h1 == r_refill_tag[1:0]) begin
              sectored_entries_7_data_1 <= _T_978;
            end
          end
        end
      end
    end
    if (_T_939) begin
      if (!(_T_961)) begin
        if (!(_T_979)) begin
          if (_T_1171) begin
            if (2'h2 == r_refill_tag[1:0]) begin
              sectored_entries_7_data_2 <= _T_978;
            end
          end
        end
      end
    end
    if (_T_939) begin
      if (!(_T_961)) begin
        if (!(_T_979)) begin
          if (_T_1171) begin
            if (2'h3 == r_refill_tag[1:0]) begin
              sectored_entries_7_data_3 <= _T_978;
            end
          end
        end
      end
    end
    if (_T_3753) begin
      sectored_entries_7_valid_0 <= 1'h0;
    end else if (io_sfence_valid) begin
      if (io_sfence_bits_rs1) begin
        if (_T_3438) begin
          if (sectored_entries_7_data_0[0]) begin
            sectored_entries_7_valid_0 <= 1'h0;
          end else if (_T_457) begin
            if (2'h0 == vpn[1:0]) begin
              sectored_entries_7_valid_0 <= 1'h0;
            end else if (_T_939) begin
              if (!(_T_961)) begin
                if (!(_T_979)) begin
                  if (_T_1171) begin
                    sectored_entries_7_valid_0 <= _GEN_238;
                  end
                end
              end
            end
          end else if (_T_939) begin
            if (!(_T_961)) begin
              if (!(_T_979)) begin
                if (_T_1171) begin
                  sectored_entries_7_valid_0 <= _GEN_238;
                end
              end
            end
          end
        end else if (_T_457) begin
          if (2'h0 == vpn[1:0]) begin
            sectored_entries_7_valid_0 <= 1'h0;
          end else if (_T_939) begin
            if (!(_T_961)) begin
              if (!(_T_979)) begin
                if (_T_1171) begin
                  sectored_entries_7_valid_0 <= _GEN_238;
                end
              end
            end
          end
        end else if (_T_939) begin
          if (!(_T_961)) begin
            if (!(_T_979)) begin
              if (_T_1171) begin
                sectored_entries_7_valid_0 <= _GEN_238;
              end
            end
          end
        end
      end else begin
        sectored_entries_7_valid_0 <= _GEN_848;
      end
    end else begin
      sectored_entries_7_valid_0 <= _GEN_542;
    end
    if (_T_3753) begin
      sectored_entries_7_valid_1 <= 1'h0;
    end else if (io_sfence_valid) begin
      if (io_sfence_bits_rs1) begin
        if (_T_3438) begin
          if (sectored_entries_7_data_1[0]) begin
            sectored_entries_7_valid_1 <= 1'h0;
          end else if (_T_457) begin
            if (2'h1 == vpn[1:0]) begin
              sectored_entries_7_valid_1 <= 1'h0;
            end else if (_T_939) begin
              if (!(_T_961)) begin
                if (!(_T_979)) begin
                  if (_T_1171) begin
                    sectored_entries_7_valid_1 <= _GEN_239;
                  end
                end
              end
            end
          end else if (_T_939) begin
            if (!(_T_961)) begin
              if (!(_T_979)) begin
                if (_T_1171) begin
                  sectored_entries_7_valid_1 <= _GEN_239;
                end
              end
            end
          end
        end else if (_T_457) begin
          if (2'h1 == vpn[1:0]) begin
            sectored_entries_7_valid_1 <= 1'h0;
          end else if (_T_939) begin
            if (!(_T_961)) begin
              if (!(_T_979)) begin
                if (_T_1171) begin
                  sectored_entries_7_valid_1 <= _GEN_239;
                end
              end
            end
          end
        end else if (_T_939) begin
          if (!(_T_961)) begin
            if (!(_T_979)) begin
              if (_T_1171) begin
                sectored_entries_7_valid_1 <= _GEN_239;
              end
            end
          end
        end
      end else begin
        sectored_entries_7_valid_1 <= _GEN_849;
      end
    end else begin
      sectored_entries_7_valid_1 <= _GEN_543;
    end
    if (_T_3753) begin
      sectored_entries_7_valid_2 <= 1'h0;
    end else if (io_sfence_valid) begin
      if (io_sfence_bits_rs1) begin
        if (_T_3438) begin
          if (sectored_entries_7_data_2[0]) begin
            sectored_entries_7_valid_2 <= 1'h0;
          end else if (_T_457) begin
            if (2'h2 == vpn[1:0]) begin
              sectored_entries_7_valid_2 <= 1'h0;
            end else if (_T_939) begin
              if (!(_T_961)) begin
                if (!(_T_979)) begin
                  if (_T_1171) begin
                    sectored_entries_7_valid_2 <= _GEN_240;
                  end
                end
              end
            end
          end else if (_T_939) begin
            if (!(_T_961)) begin
              if (!(_T_979)) begin
                if (_T_1171) begin
                  sectored_entries_7_valid_2 <= _GEN_240;
                end
              end
            end
          end
        end else if (_T_457) begin
          if (2'h2 == vpn[1:0]) begin
            sectored_entries_7_valid_2 <= 1'h0;
          end else if (_T_939) begin
            if (!(_T_961)) begin
              if (!(_T_979)) begin
                if (_T_1171) begin
                  sectored_entries_7_valid_2 <= _GEN_240;
                end
              end
            end
          end
        end else if (_T_939) begin
          if (!(_T_961)) begin
            if (!(_T_979)) begin
              if (_T_1171) begin
                sectored_entries_7_valid_2 <= _GEN_240;
              end
            end
          end
        end
      end else begin
        sectored_entries_7_valid_2 <= _GEN_850;
      end
    end else begin
      sectored_entries_7_valid_2 <= _GEN_544;
    end
    if (_T_3753) begin
      sectored_entries_7_valid_3 <= 1'h0;
    end else if (io_sfence_valid) begin
      if (io_sfence_bits_rs1) begin
        if (_T_3438) begin
          if (sectored_entries_7_data_3[0]) begin
            sectored_entries_7_valid_3 <= 1'h0;
          end else if (_T_457) begin
            if (2'h3 == vpn[1:0]) begin
              sectored_entries_7_valid_3 <= 1'h0;
            end else if (_T_939) begin
              if (!(_T_961)) begin
                if (!(_T_979)) begin
                  if (_T_1171) begin
                    sectored_entries_7_valid_3 <= _GEN_241;
                  end
                end
              end
            end
          end else if (_T_939) begin
            if (!(_T_961)) begin
              if (!(_T_979)) begin
                if (_T_1171) begin
                  sectored_entries_7_valid_3 <= _GEN_241;
                end
              end
            end
          end
        end else if (_T_457) begin
          if (2'h3 == vpn[1:0]) begin
            sectored_entries_7_valid_3 <= 1'h0;
          end else if (_T_939) begin
            if (!(_T_961)) begin
              if (!(_T_979)) begin
                if (_T_1171) begin
                  sectored_entries_7_valid_3 <= _GEN_241;
                end
              end
            end
          end
        end else if (_T_939) begin
          if (!(_T_961)) begin
            if (!(_T_979)) begin
              if (_T_1171) begin
                sectored_entries_7_valid_3 <= _GEN_241;
              end
            end
          end
        end
      end else begin
        sectored_entries_7_valid_3 <= _GEN_851;
      end
    end else begin
      sectored_entries_7_valid_3 <= _GEN_545;
    end
    if (_T_939) begin
      if (!(_T_961)) begin
        if (_T_979) begin
          if (_T_980) begin
            superpage_entries_0_tag <= r_refill_tag;
          end
        end
      end
    end
    if (_T_939) begin
      if (!(_T_961)) begin
        if (_T_979) begin
          if (_T_980) begin
            superpage_entries_0_data_0 <= _T_978;
          end
        end
      end
    end
    if (_T_3753) begin
      superpage_entries_0_valid_0 <= 1'h0;
    end else if (io_sfence_valid) begin
      if (io_sfence_bits_rs1) begin
        if (superpage_hits_0) begin
          superpage_entries_0_valid_0 <= 1'h0;
        end else if (_T_939) begin
          if (!(_T_961)) begin
            if (_T_979) begin
              superpage_entries_0_valid_0 <= _GEN_66;
            end
          end
        end
      end else begin
        superpage_entries_0_valid_0 <= _GEN_858;
      end
    end else if (_T_939) begin
      if (!(_T_961)) begin
        if (_T_979) begin
          superpage_entries_0_valid_0 <= _GEN_66;
        end
      end
    end
    if (_T_939) begin
      if (!(_T_961)) begin
        if (_T_979) begin
          if (_T_996) begin
            superpage_entries_1_tag <= r_refill_tag;
          end
        end
      end
    end
    if (_T_939) begin
      if (!(_T_961)) begin
        if (_T_979) begin
          if (_T_996) begin
            superpage_entries_1_data_0 <= _T_978;
          end
        end
      end
    end
    if (_T_3753) begin
      superpage_entries_1_valid_0 <= 1'h0;
    end else if (io_sfence_valid) begin
      if (io_sfence_bits_rs1) begin
        if (superpage_hits_1) begin
          superpage_entries_1_valid_0 <= 1'h0;
        end else if (_T_939) begin
          if (!(_T_961)) begin
            if (_T_979) begin
              superpage_entries_1_valid_0 <= _GEN_70;
            end
          end
        end
      end else begin
        superpage_entries_1_valid_0 <= _GEN_862;
      end
    end else if (_T_939) begin
      if (!(_T_961)) begin
        if (_T_979) begin
          superpage_entries_1_valid_0 <= _GEN_70;
        end
      end
    end
    if (_T_939) begin
      if (!(_T_961)) begin
        if (_T_979) begin
          if (_T_1012) begin
            superpage_entries_2_tag <= r_refill_tag;
          end
        end
      end
    end
    if (_T_939) begin
      if (!(_T_961)) begin
        if (_T_979) begin
          if (_T_1012) begin
            superpage_entries_2_data_0 <= _T_978;
          end
        end
      end
    end
    if (_T_3753) begin
      superpage_entries_2_valid_0 <= 1'h0;
    end else if (io_sfence_valid) begin
      if (io_sfence_bits_rs1) begin
        if (superpage_hits_2) begin
          superpage_entries_2_valid_0 <= 1'h0;
        end else if (_T_939) begin
          if (!(_T_961)) begin
            if (_T_979) begin
              superpage_entries_2_valid_0 <= _GEN_74;
            end
          end
        end
      end else begin
        superpage_entries_2_valid_0 <= _GEN_866;
      end
    end else if (_T_939) begin
      if (!(_T_961)) begin
        if (_T_979) begin
          superpage_entries_2_valid_0 <= _GEN_74;
        end
      end
    end
    if (_T_939) begin
      if (!(_T_961)) begin
        if (_T_979) begin
          if (_T_1028) begin
            superpage_entries_3_tag <= r_refill_tag;
          end
        end
      end
    end
    if (_T_939) begin
      if (!(_T_961)) begin
        if (_T_979) begin
          if (_T_1028) begin
            superpage_entries_3_data_0 <= _T_978;
          end
        end
      end
    end
    if (_T_3753) begin
      superpage_entries_3_valid_0 <= 1'h0;
    end else if (io_sfence_valid) begin
      if (io_sfence_bits_rs1) begin
        if (superpage_hits_3) begin
          superpage_entries_3_valid_0 <= 1'h0;
        end else if (_T_939) begin
          if (!(_T_961)) begin
            if (_T_979) begin
              superpage_entries_3_valid_0 <= _GEN_78;
            end
          end
        end
      end else begin
        superpage_entries_3_valid_0 <= _GEN_870;
      end
    end else if (_T_939) begin
      if (!(_T_961)) begin
        if (_T_979) begin
          superpage_entries_3_valid_0 <= _GEN_78;
        end
      end
    end
    if (_T_939) begin
      if (_T_961) begin
        special_entry_level <= io_ptw_resp_bits_level;
      end
    end
    if (_T_939) begin
      if (_T_961) begin
        special_entry_tag <= r_refill_tag;
      end
    end
    if (_T_939) begin
      if (_T_961) begin
        special_entry_data_0 <= _T_978;
      end
    end
    if (_T_3753) begin
      special_entry_valid_0 <= 1'h0;
    end else if (io_sfence_valid) begin
      if (io_sfence_bits_rs1) begin
        if (_T_619) begin
          special_entry_valid_0 <= 1'h0;
        end else if (_T_939) begin
          special_entry_valid_0 <= _GEN_354;
        end
      end else begin
        special_entry_valid_0 <= _GEN_874;
      end
    end else if (_T_939) begin
      special_entry_valid_0 <= _GEN_354;
    end
    if (reset) begin
      state <= 2'h0;
    end else if (io_ptw_resp_valid) begin
      state <= 2'h0;
    end else if (_T_2339) begin
      state <= 2'h3;
    end else if (_T_4) begin
      if (io_kill) begin
        state <= 2'h0;
      end else if (io_ptw_req_ready) begin
        if (io_sfence_valid) begin
          state <= 2'h3;
        end else begin
          state <= 2'h2;
        end
      end else if (io_sfence_valid) begin
        state <= 2'h0;
      end else if (_T_2222) begin
        state <= 2'h1;
      end
    end else if (_T_2222) begin
      state <= 2'h1;
    end
    if (_T_2222) begin
      r_refill_tag <= vpn;
    end
    if (_T_2222) begin
      if (_T_2233) begin
        r_superpage_repl_addr <= _T_2229;
      end else if (_T_2234[0]) begin
        r_superpage_repl_addr <= 2'h0;
      end else if (_T_2234[1]) begin
        r_superpage_repl_addr <= 2'h1;
      end else if (_T_2234[2]) begin
        r_superpage_repl_addr <= 2'h2;
      end else begin
        r_superpage_repl_addr <= 2'h3;
      end
    end
    if (_T_2222) begin
      if (_T_2293) begin
        r_sectored_repl_addr <= _T_2261;
      end else if (_T_2294[0]) begin
        r_sectored_repl_addr <= 3'h0;
      end else if (_T_2294[1]) begin
        r_sectored_repl_addr <= 3'h1;
      end else if (_T_2294[2]) begin
        r_sectored_repl_addr <= 3'h2;
      end else if (_T_2294[3]) begin
        r_sectored_repl_addr <= 3'h3;
      end else if (_T_2294[4]) begin
        r_sectored_repl_addr <= 3'h4;
      end else if (_T_2294[5]) begin
        r_sectored_repl_addr <= 3'h5;
      end else if (_T_2294[6]) begin
        r_sectored_repl_addr <= 3'h6;
      end else begin
        r_sectored_repl_addr <= 3'h7;
      end
    end
    if (_T_2222) begin
      r_sectored_hit_addr <= _T_2034;
    end
    if (_T_2222) begin
      r_sectored_hit <= _T_2016;
    end
    if (_T_2009) begin
      if (_T_2016) begin
        _T_2007 <= _T_2073;
      end
    end
    if (_T_2009) begin
      if (_T_2076) begin
        _T_2008 <= _T_2100;
      end
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_sfence_valid & _T_2346) begin
          $fwrite(32'h80000002,"Assertion failed\n    at TLB.scala:376 assert(!io.sfence.bits.rs1 || (io.sfence.bits.addr >> pgIdxBits) === vpn)\n"); // @[TLB.scala 376:13:freechips.rocketchip.system.DefaultRV32Config.fir@201971.8]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_sfence_valid & _T_2346) begin
          $fatal; // @[TLB.scala 376:13:freechips.rocketchip.system.DefaultRV32Config.fir@201972.8]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
  end
endmodule
