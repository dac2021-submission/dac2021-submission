module CompareRecFN( // @[:freechips.rocketchip.system.DefaultRV32Config.fir@211774.2]
  input  [32:0] io_a, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@211775.4]
  input  [32:0] io_b, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@211775.4]
  input         io_signaling, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@211775.4]
  output        io_lt, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@211775.4]
  output        io_eq, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@211775.4]
  output [4:0]  io_exceptionFlags // @[:freechips.rocketchip.system.DefaultRV32Config.fir@211775.4]
);
  wire  rawA_isZero; // @[rawFloatFromRecFN.scala 51:54:freechips.rocketchip.system.DefaultRV32Config.fir@211780.4]
  wire  _T_4; // @[rawFloatFromRecFN.scala 52:54:freechips.rocketchip.system.DefaultRV32Config.fir@211782.4]
  wire  rawA_isNaN; // @[rawFloatFromRecFN.scala 55:33:freechips.rocketchip.system.DefaultRV32Config.fir@211786.4]
  wire  _T_8; // @[rawFloatFromRecFN.scala 56:36:freechips.rocketchip.system.DefaultRV32Config.fir@211789.4]
  wire  rawA_isInf; // @[rawFloatFromRecFN.scala 56:33:freechips.rocketchip.system.DefaultRV32Config.fir@211790.4]
  wire  rawA_sign; // @[rawFloatFromRecFN.scala 58:25:freechips.rocketchip.system.DefaultRV32Config.fir@211793.4]
  wire [9:0] rawA_sExp; // @[rawFloatFromRecFN.scala 59:27:freechips.rocketchip.system.DefaultRV32Config.fir@211795.4]
  wire  _T_12; // @[rawFloatFromRecFN.scala 60:39:freechips.rocketchip.system.DefaultRV32Config.fir@211797.4]
  wire [24:0] rawA_sig; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@211800.4]
  wire  rawB_isZero; // @[rawFloatFromRecFN.scala 51:54:freechips.rocketchip.system.DefaultRV32Config.fir@211804.4]
  wire  _T_20; // @[rawFloatFromRecFN.scala 52:54:freechips.rocketchip.system.DefaultRV32Config.fir@211806.4]
  wire  rawB_isNaN; // @[rawFloatFromRecFN.scala 55:33:freechips.rocketchip.system.DefaultRV32Config.fir@211810.4]
  wire  _T_24; // @[rawFloatFromRecFN.scala 56:36:freechips.rocketchip.system.DefaultRV32Config.fir@211813.4]
  wire  rawB_isInf; // @[rawFloatFromRecFN.scala 56:33:freechips.rocketchip.system.DefaultRV32Config.fir@211814.4]
  wire  rawB_sign; // @[rawFloatFromRecFN.scala 58:25:freechips.rocketchip.system.DefaultRV32Config.fir@211817.4]
  wire [9:0] rawB_sExp; // @[rawFloatFromRecFN.scala 59:27:freechips.rocketchip.system.DefaultRV32Config.fir@211819.4]
  wire  _T_28; // @[rawFloatFromRecFN.scala 60:39:freechips.rocketchip.system.DefaultRV32Config.fir@211821.4]
  wire [24:0] rawB_sig; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@211824.4]
  wire  _T_32; // @[CompareRecFN.scala 57:19:freechips.rocketchip.system.DefaultRV32Config.fir@211826.4]
  wire  _T_33; // @[CompareRecFN.scala 57:35:freechips.rocketchip.system.DefaultRV32Config.fir@211827.4]
  wire  ordered; // @[CompareRecFN.scala 57:32:freechips.rocketchip.system.DefaultRV32Config.fir@211828.4]
  wire  bothInfs; // @[CompareRecFN.scala 58:33:freechips.rocketchip.system.DefaultRV32Config.fir@211829.4]
  wire  bothZeros; // @[CompareRecFN.scala 59:33:freechips.rocketchip.system.DefaultRV32Config.fir@211830.4]
  wire  eqExps; // @[CompareRecFN.scala 60:29:freechips.rocketchip.system.DefaultRV32Config.fir@211831.4]
  wire  _T_34; // @[CompareRecFN.scala 62:20:freechips.rocketchip.system.DefaultRV32Config.fir@211832.4]
  wire  _T_35; // @[CompareRecFN.scala 62:57:freechips.rocketchip.system.DefaultRV32Config.fir@211833.4]
  wire  _T_36; // @[CompareRecFN.scala 62:44:freechips.rocketchip.system.DefaultRV32Config.fir@211834.4]
  wire  common_ltMags; // @[CompareRecFN.scala 62:33:freechips.rocketchip.system.DefaultRV32Config.fir@211835.4]
  wire  _T_37; // @[CompareRecFN.scala 63:45:freechips.rocketchip.system.DefaultRV32Config.fir@211836.4]
  wire  common_eqMags; // @[CompareRecFN.scala 63:32:freechips.rocketchip.system.DefaultRV32Config.fir@211837.4]
  wire  _T_38; // @[CompareRecFN.scala 66:9:freechips.rocketchip.system.DefaultRV32Config.fir@211838.4]
  wire  _T_39; // @[CompareRecFN.scala 67:28:freechips.rocketchip.system.DefaultRV32Config.fir@211839.4]
  wire  _T_40; // @[CompareRecFN.scala 67:25:freechips.rocketchip.system.DefaultRV32Config.fir@211840.4]
  wire  _T_41; // @[CompareRecFN.scala 68:19:freechips.rocketchip.system.DefaultRV32Config.fir@211841.4]
  wire  _T_42; // @[CompareRecFN.scala 69:38:freechips.rocketchip.system.DefaultRV32Config.fir@211842.4]
  wire  _T_43; // @[CompareRecFN.scala 69:35:freechips.rocketchip.system.DefaultRV32Config.fir@211843.4]
  wire  _T_44; // @[CompareRecFN.scala 69:57:freechips.rocketchip.system.DefaultRV32Config.fir@211844.4]
  wire  _T_45; // @[CompareRecFN.scala 69:54:freechips.rocketchip.system.DefaultRV32Config.fir@211845.4]
  wire  _T_47; // @[CompareRecFN.scala 70:41:freechips.rocketchip.system.DefaultRV32Config.fir@211847.4]
  wire  _T_48; // @[CompareRecFN.scala 69:74:freechips.rocketchip.system.DefaultRV32Config.fir@211848.4]
  wire  _T_49; // @[CompareRecFN.scala 68:30:freechips.rocketchip.system.DefaultRV32Config.fir@211849.4]
  wire  _T_50; // @[CompareRecFN.scala 67:41:freechips.rocketchip.system.DefaultRV32Config.fir@211850.4]
  wire  ordered_lt; // @[CompareRecFN.scala 66:21:freechips.rocketchip.system.DefaultRV32Config.fir@211851.4]
  wire  _T_51; // @[CompareRecFN.scala 72:34:freechips.rocketchip.system.DefaultRV32Config.fir@211852.4]
  wire  _T_52; // @[CompareRecFN.scala 72:62:freechips.rocketchip.system.DefaultRV32Config.fir@211853.4]
  wire  _T_53; // @[CompareRecFN.scala 72:49:freechips.rocketchip.system.DefaultRV32Config.fir@211854.4]
  wire  ordered_eq; // @[CompareRecFN.scala 72:19:freechips.rocketchip.system.DefaultRV32Config.fir@211855.4]
  wire  _T_55; // @[common.scala 81:49:freechips.rocketchip.system.DefaultRV32Config.fir@211857.4]
  wire  _T_56; // @[common.scala 81:46:freechips.rocketchip.system.DefaultRV32Config.fir@211858.4]
  wire  _T_58; // @[common.scala 81:49:freechips.rocketchip.system.DefaultRV32Config.fir@211860.4]
  wire  _T_59; // @[common.scala 81:46:freechips.rocketchip.system.DefaultRV32Config.fir@211861.4]
  wire  _T_60; // @[CompareRecFN.scala 75:32:freechips.rocketchip.system.DefaultRV32Config.fir@211862.4]
  wire  _T_61; // @[CompareRecFN.scala 76:30:freechips.rocketchip.system.DefaultRV32Config.fir@211863.4]
  wire  _T_62; // @[CompareRecFN.scala 76:27:freechips.rocketchip.system.DefaultRV32Config.fir@211864.4]
  wire  invalid; // @[CompareRecFN.scala 75:58:freechips.rocketchip.system.DefaultRV32Config.fir@211865.4]
  assign rawA_isZero = io_a[31:29] == 3'h0; // @[rawFloatFromRecFN.scala 51:54:freechips.rocketchip.system.DefaultRV32Config.fir@211780.4]
  assign _T_4 = io_a[31:30] == 2'h3; // @[rawFloatFromRecFN.scala 52:54:freechips.rocketchip.system.DefaultRV32Config.fir@211782.4]
  assign rawA_isNaN = _T_4 & io_a[29]; // @[rawFloatFromRecFN.scala 55:33:freechips.rocketchip.system.DefaultRV32Config.fir@211786.4]
  assign _T_8 = ~io_a[29]; // @[rawFloatFromRecFN.scala 56:36:freechips.rocketchip.system.DefaultRV32Config.fir@211789.4]
  assign rawA_isInf = _T_4 & _T_8; // @[rawFloatFromRecFN.scala 56:33:freechips.rocketchip.system.DefaultRV32Config.fir@211790.4]
  assign rawA_sign = io_a[32]; // @[rawFloatFromRecFN.scala 58:25:freechips.rocketchip.system.DefaultRV32Config.fir@211793.4]
  assign rawA_sExp = {1'b0,$signed(io_a[31:23])}; // @[rawFloatFromRecFN.scala 59:27:freechips.rocketchip.system.DefaultRV32Config.fir@211795.4]
  assign _T_12 = ~rawA_isZero; // @[rawFloatFromRecFN.scala 60:39:freechips.rocketchip.system.DefaultRV32Config.fir@211797.4]
  assign rawA_sig = {1'h0,_T_12,io_a[22:0]}; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@211800.4]
  assign rawB_isZero = io_b[31:29] == 3'h0; // @[rawFloatFromRecFN.scala 51:54:freechips.rocketchip.system.DefaultRV32Config.fir@211804.4]
  assign _T_20 = io_b[31:30] == 2'h3; // @[rawFloatFromRecFN.scala 52:54:freechips.rocketchip.system.DefaultRV32Config.fir@211806.4]
  assign rawB_isNaN = _T_20 & io_b[29]; // @[rawFloatFromRecFN.scala 55:33:freechips.rocketchip.system.DefaultRV32Config.fir@211810.4]
  assign _T_24 = ~io_b[29]; // @[rawFloatFromRecFN.scala 56:36:freechips.rocketchip.system.DefaultRV32Config.fir@211813.4]
  assign rawB_isInf = _T_20 & _T_24; // @[rawFloatFromRecFN.scala 56:33:freechips.rocketchip.system.DefaultRV32Config.fir@211814.4]
  assign rawB_sign = io_b[32]; // @[rawFloatFromRecFN.scala 58:25:freechips.rocketchip.system.DefaultRV32Config.fir@211817.4]
  assign rawB_sExp = {1'b0,$signed(io_b[31:23])}; // @[rawFloatFromRecFN.scala 59:27:freechips.rocketchip.system.DefaultRV32Config.fir@211819.4]
  assign _T_28 = ~rawB_isZero; // @[rawFloatFromRecFN.scala 60:39:freechips.rocketchip.system.DefaultRV32Config.fir@211821.4]
  assign rawB_sig = {1'h0,_T_28,io_b[22:0]}; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@211824.4]
  assign _T_32 = ~rawA_isNaN; // @[CompareRecFN.scala 57:19:freechips.rocketchip.system.DefaultRV32Config.fir@211826.4]
  assign _T_33 = ~rawB_isNaN; // @[CompareRecFN.scala 57:35:freechips.rocketchip.system.DefaultRV32Config.fir@211827.4]
  assign ordered = _T_32 & _T_33; // @[CompareRecFN.scala 57:32:freechips.rocketchip.system.DefaultRV32Config.fir@211828.4]
  assign bothInfs = rawA_isInf & rawB_isInf; // @[CompareRecFN.scala 58:33:freechips.rocketchip.system.DefaultRV32Config.fir@211829.4]
  assign bothZeros = rawA_isZero & rawB_isZero; // @[CompareRecFN.scala 59:33:freechips.rocketchip.system.DefaultRV32Config.fir@211830.4]
  assign eqExps = $signed(rawA_sExp) == $signed(rawB_sExp); // @[CompareRecFN.scala 60:29:freechips.rocketchip.system.DefaultRV32Config.fir@211831.4]
  assign _T_34 = $signed(rawA_sExp) < $signed(rawB_sExp); // @[CompareRecFN.scala 62:20:freechips.rocketchip.system.DefaultRV32Config.fir@211832.4]
  assign _T_35 = rawA_sig < rawB_sig; // @[CompareRecFN.scala 62:57:freechips.rocketchip.system.DefaultRV32Config.fir@211833.4]
  assign _T_36 = eqExps & _T_35; // @[CompareRecFN.scala 62:44:freechips.rocketchip.system.DefaultRV32Config.fir@211834.4]
  assign common_ltMags = _T_34 | _T_36; // @[CompareRecFN.scala 62:33:freechips.rocketchip.system.DefaultRV32Config.fir@211835.4]
  assign _T_37 = rawA_sig == rawB_sig; // @[CompareRecFN.scala 63:45:freechips.rocketchip.system.DefaultRV32Config.fir@211836.4]
  assign common_eqMags = eqExps & _T_37; // @[CompareRecFN.scala 63:32:freechips.rocketchip.system.DefaultRV32Config.fir@211837.4]
  assign _T_38 = ~bothZeros; // @[CompareRecFN.scala 66:9:freechips.rocketchip.system.DefaultRV32Config.fir@211838.4]
  assign _T_39 = ~rawB_sign; // @[CompareRecFN.scala 67:28:freechips.rocketchip.system.DefaultRV32Config.fir@211839.4]
  assign _T_40 = rawA_sign & _T_39; // @[CompareRecFN.scala 67:25:freechips.rocketchip.system.DefaultRV32Config.fir@211840.4]
  assign _T_41 = ~bothInfs; // @[CompareRecFN.scala 68:19:freechips.rocketchip.system.DefaultRV32Config.fir@211841.4]
  assign _T_42 = ~common_ltMags; // @[CompareRecFN.scala 69:38:freechips.rocketchip.system.DefaultRV32Config.fir@211842.4]
  assign _T_43 = rawA_sign & _T_42; // @[CompareRecFN.scala 69:35:freechips.rocketchip.system.DefaultRV32Config.fir@211843.4]
  assign _T_44 = ~common_eqMags; // @[CompareRecFN.scala 69:57:freechips.rocketchip.system.DefaultRV32Config.fir@211844.4]
  assign _T_45 = _T_43 & _T_44; // @[CompareRecFN.scala 69:54:freechips.rocketchip.system.DefaultRV32Config.fir@211845.4]
  assign _T_47 = _T_39 & common_ltMags; // @[CompareRecFN.scala 70:41:freechips.rocketchip.system.DefaultRV32Config.fir@211847.4]
  assign _T_48 = _T_45 | _T_47; // @[CompareRecFN.scala 69:74:freechips.rocketchip.system.DefaultRV32Config.fir@211848.4]
  assign _T_49 = _T_41 & _T_48; // @[CompareRecFN.scala 68:30:freechips.rocketchip.system.DefaultRV32Config.fir@211849.4]
  assign _T_50 = _T_40 | _T_49; // @[CompareRecFN.scala 67:41:freechips.rocketchip.system.DefaultRV32Config.fir@211850.4]
  assign ordered_lt = _T_38 & _T_50; // @[CompareRecFN.scala 66:21:freechips.rocketchip.system.DefaultRV32Config.fir@211851.4]
  assign _T_51 = rawA_sign == rawB_sign; // @[CompareRecFN.scala 72:34:freechips.rocketchip.system.DefaultRV32Config.fir@211852.4]
  assign _T_52 = bothInfs | common_eqMags; // @[CompareRecFN.scala 72:62:freechips.rocketchip.system.DefaultRV32Config.fir@211853.4]
  assign _T_53 = _T_51 & _T_52; // @[CompareRecFN.scala 72:49:freechips.rocketchip.system.DefaultRV32Config.fir@211854.4]
  assign ordered_eq = bothZeros | _T_53; // @[CompareRecFN.scala 72:19:freechips.rocketchip.system.DefaultRV32Config.fir@211855.4]
  assign _T_55 = ~rawA_sig[22]; // @[common.scala 81:49:freechips.rocketchip.system.DefaultRV32Config.fir@211857.4]
  assign _T_56 = rawA_isNaN & _T_55; // @[common.scala 81:46:freechips.rocketchip.system.DefaultRV32Config.fir@211858.4]
  assign _T_58 = ~rawB_sig[22]; // @[common.scala 81:49:freechips.rocketchip.system.DefaultRV32Config.fir@211860.4]
  assign _T_59 = rawB_isNaN & _T_58; // @[common.scala 81:46:freechips.rocketchip.system.DefaultRV32Config.fir@211861.4]
  assign _T_60 = _T_56 | _T_59; // @[CompareRecFN.scala 75:32:freechips.rocketchip.system.DefaultRV32Config.fir@211862.4]
  assign _T_61 = ~ordered; // @[CompareRecFN.scala 76:30:freechips.rocketchip.system.DefaultRV32Config.fir@211863.4]
  assign _T_62 = io_signaling & _T_61; // @[CompareRecFN.scala 76:27:freechips.rocketchip.system.DefaultRV32Config.fir@211864.4]
  assign invalid = _T_60 | _T_62; // @[CompareRecFN.scala 75:58:freechips.rocketchip.system.DefaultRV32Config.fir@211865.4]
  assign io_lt = ordered & ordered_lt; // @[CompareRecFN.scala 78:11:freechips.rocketchip.system.DefaultRV32Config.fir@211867.4]
  assign io_eq = ordered & ordered_eq; // @[CompareRecFN.scala 79:11:freechips.rocketchip.system.DefaultRV32Config.fir@211869.4]
  assign io_exceptionFlags = {invalid,4'h0}; // @[CompareRecFN.scala 81:23:freechips.rocketchip.system.DefaultRV32Config.fir@211876.4]
endmodule
