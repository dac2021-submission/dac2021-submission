module AXI4Deinterleaver( // @[:freechips.rocketchip.system.DefaultRV32Config.fir@24171.2]
  input         clock, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@24172.4]
  input         reset, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@24173.4]
  output        auto_in_aw_ready, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@24174.4]
  input         auto_in_aw_valid, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@24174.4]
  input  [3:0]  auto_in_aw_bits_id, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@24174.4]
  input  [30:0] auto_in_aw_bits_addr, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@24174.4]
  input  [7:0]  auto_in_aw_bits_len, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@24174.4]
  input  [2:0]  auto_in_aw_bits_size, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@24174.4]
  input  [1:0]  auto_in_aw_bits_burst, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@24174.4]
  input         auto_in_aw_bits_lock, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@24174.4]
  input  [3:0]  auto_in_aw_bits_cache, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@24174.4]
  input  [2:0]  auto_in_aw_bits_prot, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@24174.4]
  input  [3:0]  auto_in_aw_bits_qos, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@24174.4]
  input  [3:0]  auto_in_aw_bits_echo_tl_state_size, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@24174.4]
  input  [4:0]  auto_in_aw_bits_echo_tl_state_source, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@24174.4]
  output        auto_in_w_ready, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@24174.4]
  input         auto_in_w_valid, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@24174.4]
  input  [31:0] auto_in_w_bits_data, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@24174.4]
  input  [3:0]  auto_in_w_bits_strb, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@24174.4]
  input         auto_in_w_bits_last, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@24174.4]
  input         auto_in_b_ready, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@24174.4]
  output        auto_in_b_valid, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@24174.4]
  output [3:0]  auto_in_b_bits_id, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@24174.4]
  output [1:0]  auto_in_b_bits_resp, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@24174.4]
  output [3:0]  auto_in_b_bits_echo_tl_state_size, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@24174.4]
  output [4:0]  auto_in_b_bits_echo_tl_state_source, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@24174.4]
  output        auto_in_ar_ready, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@24174.4]
  input         auto_in_ar_valid, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@24174.4]
  input  [3:0]  auto_in_ar_bits_id, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@24174.4]
  input  [30:0] auto_in_ar_bits_addr, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@24174.4]
  input  [7:0]  auto_in_ar_bits_len, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@24174.4]
  input  [2:0]  auto_in_ar_bits_size, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@24174.4]
  input  [1:0]  auto_in_ar_bits_burst, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@24174.4]
  input         auto_in_ar_bits_lock, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@24174.4]
  input  [3:0]  auto_in_ar_bits_cache, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@24174.4]
  input  [2:0]  auto_in_ar_bits_prot, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@24174.4]
  input  [3:0]  auto_in_ar_bits_qos, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@24174.4]
  input  [3:0]  auto_in_ar_bits_echo_tl_state_size, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@24174.4]
  input  [4:0]  auto_in_ar_bits_echo_tl_state_source, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@24174.4]
  input         auto_in_r_ready, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@24174.4]
  output        auto_in_r_valid, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@24174.4]
  output [3:0]  auto_in_r_bits_id, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@24174.4]
  output [31:0] auto_in_r_bits_data, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@24174.4]
  output [1:0]  auto_in_r_bits_resp, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@24174.4]
  output [3:0]  auto_in_r_bits_echo_tl_state_size, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@24174.4]
  output [4:0]  auto_in_r_bits_echo_tl_state_source, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@24174.4]
  output        auto_in_r_bits_last, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@24174.4]
  input         auto_out_aw_ready, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@24174.4]
  output        auto_out_aw_valid, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@24174.4]
  output [3:0]  auto_out_aw_bits_id, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@24174.4]
  output [30:0] auto_out_aw_bits_addr, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@24174.4]
  output [7:0]  auto_out_aw_bits_len, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@24174.4]
  output [2:0]  auto_out_aw_bits_size, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@24174.4]
  output [1:0]  auto_out_aw_bits_burst, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@24174.4]
  output        auto_out_aw_bits_lock, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@24174.4]
  output [3:0]  auto_out_aw_bits_cache, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@24174.4]
  output [2:0]  auto_out_aw_bits_prot, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@24174.4]
  output [3:0]  auto_out_aw_bits_qos, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@24174.4]
  output [3:0]  auto_out_aw_bits_echo_tl_state_size, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@24174.4]
  output [4:0]  auto_out_aw_bits_echo_tl_state_source, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@24174.4]
  input         auto_out_w_ready, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@24174.4]
  output        auto_out_w_valid, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@24174.4]
  output [31:0] auto_out_w_bits_data, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@24174.4]
  output [3:0]  auto_out_w_bits_strb, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@24174.4]
  output        auto_out_w_bits_last, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@24174.4]
  output        auto_out_b_ready, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@24174.4]
  input         auto_out_b_valid, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@24174.4]
  input  [3:0]  auto_out_b_bits_id, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@24174.4]
  input  [1:0]  auto_out_b_bits_resp, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@24174.4]
  input  [3:0]  auto_out_b_bits_echo_tl_state_size, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@24174.4]
  input  [4:0]  auto_out_b_bits_echo_tl_state_source, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@24174.4]
  input         auto_out_ar_ready, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@24174.4]
  output        auto_out_ar_valid, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@24174.4]
  output [3:0]  auto_out_ar_bits_id, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@24174.4]
  output [30:0] auto_out_ar_bits_addr, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@24174.4]
  output [7:0]  auto_out_ar_bits_len, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@24174.4]
  output [2:0]  auto_out_ar_bits_size, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@24174.4]
  output [1:0]  auto_out_ar_bits_burst, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@24174.4]
  output        auto_out_ar_bits_lock, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@24174.4]
  output [3:0]  auto_out_ar_bits_cache, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@24174.4]
  output [2:0]  auto_out_ar_bits_prot, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@24174.4]
  output [3:0]  auto_out_ar_bits_qos, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@24174.4]
  output [3:0]  auto_out_ar_bits_echo_tl_state_size, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@24174.4]
  output [4:0]  auto_out_ar_bits_echo_tl_state_source, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@24174.4]
  output        auto_out_r_ready, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@24174.4]
  input         auto_out_r_valid, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@24174.4]
  input  [3:0]  auto_out_r_bits_id, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@24174.4]
  input  [31:0] auto_out_r_bits_data, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@24174.4]
  input  [1:0]  auto_out_r_bits_resp, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@24174.4]
  input  [3:0]  auto_out_r_bits_echo_tl_state_size, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@24174.4]
  input  [4:0]  auto_out_r_bits_echo_tl_state_source, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@24174.4]
  input         auto_out_r_bits_last // @[:freechips.rocketchip.system.DefaultRV32Config.fir@24174.4]
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
`endif // RANDOMIZE_REG_INIT
  wire  queue_0_clock; // @[Deinterleaver.scala 44:27:freechips.rocketchip.system.DefaultRV32Config.fir@24222.4]
  wire  queue_0_reset; // @[Deinterleaver.scala 44:27:freechips.rocketchip.system.DefaultRV32Config.fir@24222.4]
  wire  queue_0_io_enq_ready; // @[Deinterleaver.scala 44:27:freechips.rocketchip.system.DefaultRV32Config.fir@24222.4]
  wire  queue_0_io_enq_valid; // @[Deinterleaver.scala 44:27:freechips.rocketchip.system.DefaultRV32Config.fir@24222.4]
  wire [3:0] queue_0_io_enq_bits_id; // @[Deinterleaver.scala 44:27:freechips.rocketchip.system.DefaultRV32Config.fir@24222.4]
  wire [31:0] queue_0_io_enq_bits_data; // @[Deinterleaver.scala 44:27:freechips.rocketchip.system.DefaultRV32Config.fir@24222.4]
  wire [1:0] queue_0_io_enq_bits_resp; // @[Deinterleaver.scala 44:27:freechips.rocketchip.system.DefaultRV32Config.fir@24222.4]
  wire [3:0] queue_0_io_enq_bits_echo_tl_state_size; // @[Deinterleaver.scala 44:27:freechips.rocketchip.system.DefaultRV32Config.fir@24222.4]
  wire [4:0] queue_0_io_enq_bits_echo_tl_state_source; // @[Deinterleaver.scala 44:27:freechips.rocketchip.system.DefaultRV32Config.fir@24222.4]
  wire  queue_0_io_enq_bits_last; // @[Deinterleaver.scala 44:27:freechips.rocketchip.system.DefaultRV32Config.fir@24222.4]
  wire  queue_0_io_deq_ready; // @[Deinterleaver.scala 44:27:freechips.rocketchip.system.DefaultRV32Config.fir@24222.4]
  wire  queue_0_io_deq_valid; // @[Deinterleaver.scala 44:27:freechips.rocketchip.system.DefaultRV32Config.fir@24222.4]
  wire [3:0] queue_0_io_deq_bits_id; // @[Deinterleaver.scala 44:27:freechips.rocketchip.system.DefaultRV32Config.fir@24222.4]
  wire [31:0] queue_0_io_deq_bits_data; // @[Deinterleaver.scala 44:27:freechips.rocketchip.system.DefaultRV32Config.fir@24222.4]
  wire [1:0] queue_0_io_deq_bits_resp; // @[Deinterleaver.scala 44:27:freechips.rocketchip.system.DefaultRV32Config.fir@24222.4]
  wire [3:0] queue_0_io_deq_bits_echo_tl_state_size; // @[Deinterleaver.scala 44:27:freechips.rocketchip.system.DefaultRV32Config.fir@24222.4]
  wire [4:0] queue_0_io_deq_bits_echo_tl_state_source; // @[Deinterleaver.scala 44:27:freechips.rocketchip.system.DefaultRV32Config.fir@24222.4]
  wire  queue_0_io_deq_bits_last; // @[Deinterleaver.scala 44:27:freechips.rocketchip.system.DefaultRV32Config.fir@24222.4]
  wire  queue_1_clock; // @[Deinterleaver.scala 44:27:freechips.rocketchip.system.DefaultRV32Config.fir@24225.4]
  wire  queue_1_reset; // @[Deinterleaver.scala 44:27:freechips.rocketchip.system.DefaultRV32Config.fir@24225.4]
  wire  queue_1_io_enq_ready; // @[Deinterleaver.scala 44:27:freechips.rocketchip.system.DefaultRV32Config.fir@24225.4]
  wire  queue_1_io_enq_valid; // @[Deinterleaver.scala 44:27:freechips.rocketchip.system.DefaultRV32Config.fir@24225.4]
  wire [3:0] queue_1_io_enq_bits_id; // @[Deinterleaver.scala 44:27:freechips.rocketchip.system.DefaultRV32Config.fir@24225.4]
  wire [31:0] queue_1_io_enq_bits_data; // @[Deinterleaver.scala 44:27:freechips.rocketchip.system.DefaultRV32Config.fir@24225.4]
  wire [1:0] queue_1_io_enq_bits_resp; // @[Deinterleaver.scala 44:27:freechips.rocketchip.system.DefaultRV32Config.fir@24225.4]
  wire [3:0] queue_1_io_enq_bits_echo_tl_state_size; // @[Deinterleaver.scala 44:27:freechips.rocketchip.system.DefaultRV32Config.fir@24225.4]
  wire [4:0] queue_1_io_enq_bits_echo_tl_state_source; // @[Deinterleaver.scala 44:27:freechips.rocketchip.system.DefaultRV32Config.fir@24225.4]
  wire  queue_1_io_enq_bits_last; // @[Deinterleaver.scala 44:27:freechips.rocketchip.system.DefaultRV32Config.fir@24225.4]
  wire  queue_1_io_deq_ready; // @[Deinterleaver.scala 44:27:freechips.rocketchip.system.DefaultRV32Config.fir@24225.4]
  wire  queue_1_io_deq_valid; // @[Deinterleaver.scala 44:27:freechips.rocketchip.system.DefaultRV32Config.fir@24225.4]
  wire [3:0] queue_1_io_deq_bits_id; // @[Deinterleaver.scala 44:27:freechips.rocketchip.system.DefaultRV32Config.fir@24225.4]
  wire [31:0] queue_1_io_deq_bits_data; // @[Deinterleaver.scala 44:27:freechips.rocketchip.system.DefaultRV32Config.fir@24225.4]
  wire [1:0] queue_1_io_deq_bits_resp; // @[Deinterleaver.scala 44:27:freechips.rocketchip.system.DefaultRV32Config.fir@24225.4]
  wire [3:0] queue_1_io_deq_bits_echo_tl_state_size; // @[Deinterleaver.scala 44:27:freechips.rocketchip.system.DefaultRV32Config.fir@24225.4]
  wire [4:0] queue_1_io_deq_bits_echo_tl_state_source; // @[Deinterleaver.scala 44:27:freechips.rocketchip.system.DefaultRV32Config.fir@24225.4]
  wire  queue_1_io_deq_bits_last; // @[Deinterleaver.scala 44:27:freechips.rocketchip.system.DefaultRV32Config.fir@24225.4]
  wire  queue_2_clock; // @[Deinterleaver.scala 44:27:freechips.rocketchip.system.DefaultRV32Config.fir@24228.4]
  wire  queue_2_reset; // @[Deinterleaver.scala 44:27:freechips.rocketchip.system.DefaultRV32Config.fir@24228.4]
  wire  queue_2_io_enq_ready; // @[Deinterleaver.scala 44:27:freechips.rocketchip.system.DefaultRV32Config.fir@24228.4]
  wire  queue_2_io_enq_valid; // @[Deinterleaver.scala 44:27:freechips.rocketchip.system.DefaultRV32Config.fir@24228.4]
  wire [3:0] queue_2_io_enq_bits_id; // @[Deinterleaver.scala 44:27:freechips.rocketchip.system.DefaultRV32Config.fir@24228.4]
  wire [31:0] queue_2_io_enq_bits_data; // @[Deinterleaver.scala 44:27:freechips.rocketchip.system.DefaultRV32Config.fir@24228.4]
  wire [1:0] queue_2_io_enq_bits_resp; // @[Deinterleaver.scala 44:27:freechips.rocketchip.system.DefaultRV32Config.fir@24228.4]
  wire [3:0] queue_2_io_enq_bits_echo_tl_state_size; // @[Deinterleaver.scala 44:27:freechips.rocketchip.system.DefaultRV32Config.fir@24228.4]
  wire [4:0] queue_2_io_enq_bits_echo_tl_state_source; // @[Deinterleaver.scala 44:27:freechips.rocketchip.system.DefaultRV32Config.fir@24228.4]
  wire  queue_2_io_enq_bits_last; // @[Deinterleaver.scala 44:27:freechips.rocketchip.system.DefaultRV32Config.fir@24228.4]
  wire  queue_2_io_deq_ready; // @[Deinterleaver.scala 44:27:freechips.rocketchip.system.DefaultRV32Config.fir@24228.4]
  wire  queue_2_io_deq_valid; // @[Deinterleaver.scala 44:27:freechips.rocketchip.system.DefaultRV32Config.fir@24228.4]
  wire [3:0] queue_2_io_deq_bits_id; // @[Deinterleaver.scala 44:27:freechips.rocketchip.system.DefaultRV32Config.fir@24228.4]
  wire [31:0] queue_2_io_deq_bits_data; // @[Deinterleaver.scala 44:27:freechips.rocketchip.system.DefaultRV32Config.fir@24228.4]
  wire [1:0] queue_2_io_deq_bits_resp; // @[Deinterleaver.scala 44:27:freechips.rocketchip.system.DefaultRV32Config.fir@24228.4]
  wire [3:0] queue_2_io_deq_bits_echo_tl_state_size; // @[Deinterleaver.scala 44:27:freechips.rocketchip.system.DefaultRV32Config.fir@24228.4]
  wire [4:0] queue_2_io_deq_bits_echo_tl_state_source; // @[Deinterleaver.scala 44:27:freechips.rocketchip.system.DefaultRV32Config.fir@24228.4]
  wire  queue_2_io_deq_bits_last; // @[Deinterleaver.scala 44:27:freechips.rocketchip.system.DefaultRV32Config.fir@24228.4]
  wire  queue_3_clock; // @[Deinterleaver.scala 44:27:freechips.rocketchip.system.DefaultRV32Config.fir@24231.4]
  wire  queue_3_reset; // @[Deinterleaver.scala 44:27:freechips.rocketchip.system.DefaultRV32Config.fir@24231.4]
  wire  queue_3_io_enq_ready; // @[Deinterleaver.scala 44:27:freechips.rocketchip.system.DefaultRV32Config.fir@24231.4]
  wire  queue_3_io_enq_valid; // @[Deinterleaver.scala 44:27:freechips.rocketchip.system.DefaultRV32Config.fir@24231.4]
  wire [3:0] queue_3_io_enq_bits_id; // @[Deinterleaver.scala 44:27:freechips.rocketchip.system.DefaultRV32Config.fir@24231.4]
  wire [31:0] queue_3_io_enq_bits_data; // @[Deinterleaver.scala 44:27:freechips.rocketchip.system.DefaultRV32Config.fir@24231.4]
  wire [1:0] queue_3_io_enq_bits_resp; // @[Deinterleaver.scala 44:27:freechips.rocketchip.system.DefaultRV32Config.fir@24231.4]
  wire [3:0] queue_3_io_enq_bits_echo_tl_state_size; // @[Deinterleaver.scala 44:27:freechips.rocketchip.system.DefaultRV32Config.fir@24231.4]
  wire [4:0] queue_3_io_enq_bits_echo_tl_state_source; // @[Deinterleaver.scala 44:27:freechips.rocketchip.system.DefaultRV32Config.fir@24231.4]
  wire  queue_3_io_enq_bits_last; // @[Deinterleaver.scala 44:27:freechips.rocketchip.system.DefaultRV32Config.fir@24231.4]
  wire  queue_3_io_deq_ready; // @[Deinterleaver.scala 44:27:freechips.rocketchip.system.DefaultRV32Config.fir@24231.4]
  wire  queue_3_io_deq_valid; // @[Deinterleaver.scala 44:27:freechips.rocketchip.system.DefaultRV32Config.fir@24231.4]
  wire [3:0] queue_3_io_deq_bits_id; // @[Deinterleaver.scala 44:27:freechips.rocketchip.system.DefaultRV32Config.fir@24231.4]
  wire [31:0] queue_3_io_deq_bits_data; // @[Deinterleaver.scala 44:27:freechips.rocketchip.system.DefaultRV32Config.fir@24231.4]
  wire [1:0] queue_3_io_deq_bits_resp; // @[Deinterleaver.scala 44:27:freechips.rocketchip.system.DefaultRV32Config.fir@24231.4]
  wire [3:0] queue_3_io_deq_bits_echo_tl_state_size; // @[Deinterleaver.scala 44:27:freechips.rocketchip.system.DefaultRV32Config.fir@24231.4]
  wire [4:0] queue_3_io_deq_bits_echo_tl_state_source; // @[Deinterleaver.scala 44:27:freechips.rocketchip.system.DefaultRV32Config.fir@24231.4]
  wire  queue_3_io_deq_bits_last; // @[Deinterleaver.scala 44:27:freechips.rocketchip.system.DefaultRV32Config.fir@24231.4]
  wire  queue_4_clock; // @[Deinterleaver.scala 44:27:freechips.rocketchip.system.DefaultRV32Config.fir@24234.4]
  wire  queue_4_reset; // @[Deinterleaver.scala 44:27:freechips.rocketchip.system.DefaultRV32Config.fir@24234.4]
  wire  queue_4_io_enq_ready; // @[Deinterleaver.scala 44:27:freechips.rocketchip.system.DefaultRV32Config.fir@24234.4]
  wire  queue_4_io_enq_valid; // @[Deinterleaver.scala 44:27:freechips.rocketchip.system.DefaultRV32Config.fir@24234.4]
  wire [3:0] queue_4_io_enq_bits_id; // @[Deinterleaver.scala 44:27:freechips.rocketchip.system.DefaultRV32Config.fir@24234.4]
  wire [31:0] queue_4_io_enq_bits_data; // @[Deinterleaver.scala 44:27:freechips.rocketchip.system.DefaultRV32Config.fir@24234.4]
  wire [1:0] queue_4_io_enq_bits_resp; // @[Deinterleaver.scala 44:27:freechips.rocketchip.system.DefaultRV32Config.fir@24234.4]
  wire [3:0] queue_4_io_enq_bits_echo_tl_state_size; // @[Deinterleaver.scala 44:27:freechips.rocketchip.system.DefaultRV32Config.fir@24234.4]
  wire [4:0] queue_4_io_enq_bits_echo_tl_state_source; // @[Deinterleaver.scala 44:27:freechips.rocketchip.system.DefaultRV32Config.fir@24234.4]
  wire  queue_4_io_enq_bits_last; // @[Deinterleaver.scala 44:27:freechips.rocketchip.system.DefaultRV32Config.fir@24234.4]
  wire  queue_4_io_deq_ready; // @[Deinterleaver.scala 44:27:freechips.rocketchip.system.DefaultRV32Config.fir@24234.4]
  wire  queue_4_io_deq_valid; // @[Deinterleaver.scala 44:27:freechips.rocketchip.system.DefaultRV32Config.fir@24234.4]
  wire [3:0] queue_4_io_deq_bits_id; // @[Deinterleaver.scala 44:27:freechips.rocketchip.system.DefaultRV32Config.fir@24234.4]
  wire [31:0] queue_4_io_deq_bits_data; // @[Deinterleaver.scala 44:27:freechips.rocketchip.system.DefaultRV32Config.fir@24234.4]
  wire [1:0] queue_4_io_deq_bits_resp; // @[Deinterleaver.scala 44:27:freechips.rocketchip.system.DefaultRV32Config.fir@24234.4]
  wire [3:0] queue_4_io_deq_bits_echo_tl_state_size; // @[Deinterleaver.scala 44:27:freechips.rocketchip.system.DefaultRV32Config.fir@24234.4]
  wire [4:0] queue_4_io_deq_bits_echo_tl_state_source; // @[Deinterleaver.scala 44:27:freechips.rocketchip.system.DefaultRV32Config.fir@24234.4]
  wire  queue_4_io_deq_bits_last; // @[Deinterleaver.scala 44:27:freechips.rocketchip.system.DefaultRV32Config.fir@24234.4]
  wire [15:0] _T_52; // @[OneHot.scala 65:12:freechips.rocketchip.system.DefaultRV32Config.fir@24529.4]
  wire  queue_wire_5_enq_valid; // @[Deinterleaver.scala 108:28:freechips.rocketchip.system.DefaultRV32Config.fir@25019.4]
  wire  _T_2; // @[Deinterleaver.scala 53:20:freechips.rocketchip.system.DefaultRV32Config.fir@24238.4]
  wire  _T_4; // @[Deinterleaver.scala 53:19:freechips.rocketchip.system.DefaultRV32Config.fir@24240.4]
  wire  _T_5; // @[Deinterleaver.scala 53:19:freechips.rocketchip.system.DefaultRV32Config.fir@24241.4]
  wire  queue_wire_6_enq_valid; // @[Deinterleaver.scala 108:28:freechips.rocketchip.system.DefaultRV32Config.fir@25027.4]
  wire  _T_6; // @[Deinterleaver.scala 53:20:freechips.rocketchip.system.DefaultRV32Config.fir@24264.4]
  wire  _T_8; // @[Deinterleaver.scala 53:19:freechips.rocketchip.system.DefaultRV32Config.fir@24266.4]
  wire  _T_9; // @[Deinterleaver.scala 53:19:freechips.rocketchip.system.DefaultRV32Config.fir@24267.4]
  wire  queue_wire_7_enq_valid; // @[Deinterleaver.scala 108:28:freechips.rocketchip.system.DefaultRV32Config.fir@25035.4]
  wire  _T_10; // @[Deinterleaver.scala 53:20:freechips.rocketchip.system.DefaultRV32Config.fir@24290.4]
  wire  _T_12; // @[Deinterleaver.scala 53:19:freechips.rocketchip.system.DefaultRV32Config.fir@24292.4]
  wire  _T_13; // @[Deinterleaver.scala 53:19:freechips.rocketchip.system.DefaultRV32Config.fir@24293.4]
  wire  queue_wire_8_enq_valid; // @[Deinterleaver.scala 108:28:freechips.rocketchip.system.DefaultRV32Config.fir@25043.4]
  wire  _T_14; // @[Deinterleaver.scala 53:20:freechips.rocketchip.system.DefaultRV32Config.fir@24316.4]
  wire  _T_16; // @[Deinterleaver.scala 53:19:freechips.rocketchip.system.DefaultRV32Config.fir@24318.4]
  wire  _T_17; // @[Deinterleaver.scala 53:19:freechips.rocketchip.system.DefaultRV32Config.fir@24319.4]
  wire  queue_wire_9_enq_valid; // @[Deinterleaver.scala 108:28:freechips.rocketchip.system.DefaultRV32Config.fir@25051.4]
  wire  _T_18; // @[Deinterleaver.scala 53:20:freechips.rocketchip.system.DefaultRV32Config.fir@24342.4]
  wire  _T_20; // @[Deinterleaver.scala 53:19:freechips.rocketchip.system.DefaultRV32Config.fir@24344.4]
  wire  _T_21; // @[Deinterleaver.scala 53:19:freechips.rocketchip.system.DefaultRV32Config.fir@24345.4]
  wire  queue_wire_10_enq_valid; // @[Deinterleaver.scala 108:28:freechips.rocketchip.system.DefaultRV32Config.fir@25059.4]
  wire  _T_22; // @[Deinterleaver.scala 53:20:freechips.rocketchip.system.DefaultRV32Config.fir@24368.4]
  wire  _T_24; // @[Deinterleaver.scala 53:19:freechips.rocketchip.system.DefaultRV32Config.fir@24370.4]
  wire  _T_25; // @[Deinterleaver.scala 53:19:freechips.rocketchip.system.DefaultRV32Config.fir@24371.4]
  wire  queue_wire_11_enq_valid; // @[Deinterleaver.scala 108:28:freechips.rocketchip.system.DefaultRV32Config.fir@25067.4]
  wire  _T_26; // @[Deinterleaver.scala 53:20:freechips.rocketchip.system.DefaultRV32Config.fir@24394.4]
  wire  _T_28; // @[Deinterleaver.scala 53:19:freechips.rocketchip.system.DefaultRV32Config.fir@24396.4]
  wire  _T_29; // @[Deinterleaver.scala 53:19:freechips.rocketchip.system.DefaultRV32Config.fir@24397.4]
  wire  queue_wire_12_enq_valid; // @[Deinterleaver.scala 108:28:freechips.rocketchip.system.DefaultRV32Config.fir@25075.4]
  wire  _T_30; // @[Deinterleaver.scala 53:20:freechips.rocketchip.system.DefaultRV32Config.fir@24420.4]
  wire  _T_32; // @[Deinterleaver.scala 53:19:freechips.rocketchip.system.DefaultRV32Config.fir@24422.4]
  wire  _T_33; // @[Deinterleaver.scala 53:19:freechips.rocketchip.system.DefaultRV32Config.fir@24423.4]
  wire  queue_wire_13_enq_valid; // @[Deinterleaver.scala 108:28:freechips.rocketchip.system.DefaultRV32Config.fir@25083.4]
  wire  _T_34; // @[Deinterleaver.scala 53:20:freechips.rocketchip.system.DefaultRV32Config.fir@24446.4]
  wire  _T_36; // @[Deinterleaver.scala 53:19:freechips.rocketchip.system.DefaultRV32Config.fir@24448.4]
  wire  _T_37; // @[Deinterleaver.scala 53:19:freechips.rocketchip.system.DefaultRV32Config.fir@24449.4]
  wire  queue_wire_14_enq_valid; // @[Deinterleaver.scala 108:28:freechips.rocketchip.system.DefaultRV32Config.fir@25091.4]
  wire  _T_38; // @[Deinterleaver.scala 53:20:freechips.rocketchip.system.DefaultRV32Config.fir@24472.4]
  wire  _T_40; // @[Deinterleaver.scala 53:19:freechips.rocketchip.system.DefaultRV32Config.fir@24474.4]
  wire  _T_41; // @[Deinterleaver.scala 53:19:freechips.rocketchip.system.DefaultRV32Config.fir@24475.4]
  wire  queue_wire_15_enq_valid; // @[Deinterleaver.scala 108:28:freechips.rocketchip.system.DefaultRV32Config.fir@25099.4]
  wire  _T_42; // @[Deinterleaver.scala 53:20:freechips.rocketchip.system.DefaultRV32Config.fir@24498.4]
  wire  _T_44; // @[Deinterleaver.scala 53:19:freechips.rocketchip.system.DefaultRV32Config.fir@24500.4]
  wire  _T_45; // @[Deinterleaver.scala 53:19:freechips.rocketchip.system.DefaultRV32Config.fir@24501.4]
  reg  _T_46; // @[Deinterleaver.scala 60:29:freechips.rocketchip.system.DefaultRV32Config.fir@24523.4]
  reg [3:0] _T_47; // @[Deinterleaver.scala 61:25:freechips.rocketchip.system.DefaultRV32Config.fir@24524.4]
  wire [15:0] _T_49; // @[OneHot.scala 65:12:freechips.rocketchip.system.DefaultRV32Config.fir@24526.4]
  reg [4:0] _T_54; // @[Deinterleaver.scala 72:32:freechips.rocketchip.system.DefaultRV32Config.fir@24531.4]
  wire  _T_311_4; // @[Deinterleaver.scala 105:33:freechips.rocketchip.system.DefaultRV32Config.fir@24961.4 Deinterleaver.scala 105:33:freechips.rocketchip.system.DefaultRV32Config.fir@24966.4]
  wire  _T_311_3; // @[Deinterleaver.scala 105:33:freechips.rocketchip.system.DefaultRV32Config.fir@24961.4 Deinterleaver.scala 105:33:freechips.rocketchip.system.DefaultRV32Config.fir@24965.4]
  wire  _T_311_2; // @[Deinterleaver.scala 105:33:freechips.rocketchip.system.DefaultRV32Config.fir@24961.4 Deinterleaver.scala 105:33:freechips.rocketchip.system.DefaultRV32Config.fir@24964.4]
  wire  _T_311_1; // @[Deinterleaver.scala 105:33:freechips.rocketchip.system.DefaultRV32Config.fir@24961.4 Deinterleaver.scala 105:33:freechips.rocketchip.system.DefaultRV32Config.fir@24963.4]
  wire  _T_311_0; // @[Deinterleaver.scala 105:33:freechips.rocketchip.system.DefaultRV32Config.fir@24961.4 Deinterleaver.scala 105:33:freechips.rocketchip.system.DefaultRV32Config.fir@24962.4]
  wire  _GEN_99; // @[Deinterleaver.scala 106:21:freechips.rocketchip.system.DefaultRV32Config.fir@24978.4]
  wire  _GEN_100; // @[Deinterleaver.scala 106:21:freechips.rocketchip.system.DefaultRV32Config.fir@24978.4]
  wire  _GEN_101; // @[Deinterleaver.scala 106:21:freechips.rocketchip.system.DefaultRV32Config.fir@24978.4]
  wire  _GEN_102; // @[Deinterleaver.scala 106:21:freechips.rocketchip.system.DefaultRV32Config.fir@24978.4]
  wire  _GEN_103; // @[Deinterleaver.scala 106:21:freechips.rocketchip.system.DefaultRV32Config.fir@24978.4]
  wire  _GEN_104; // @[Deinterleaver.scala 106:21:freechips.rocketchip.system.DefaultRV32Config.fir@24978.4]
  wire  _GEN_105; // @[Deinterleaver.scala 106:21:freechips.rocketchip.system.DefaultRV32Config.fir@24978.4]
  wire  _GEN_106; // @[Deinterleaver.scala 106:21:freechips.rocketchip.system.DefaultRV32Config.fir@24978.4]
  wire  _GEN_107; // @[Deinterleaver.scala 106:21:freechips.rocketchip.system.DefaultRV32Config.fir@24978.4]
  wire  _GEN_108; // @[Deinterleaver.scala 106:21:freechips.rocketchip.system.DefaultRV32Config.fir@24978.4]
  wire  _GEN_109; // @[Deinterleaver.scala 106:21:freechips.rocketchip.system.DefaultRV32Config.fir@24978.4]
  wire  _GEN_110; // @[Deinterleaver.scala 106:21:freechips.rocketchip.system.DefaultRV32Config.fir@24978.4]
  wire  _GEN_111; // @[Deinterleaver.scala 106:21:freechips.rocketchip.system.DefaultRV32Config.fir@24978.4]
  wire  _GEN_112; // @[Deinterleaver.scala 106:21:freechips.rocketchip.system.DefaultRV32Config.fir@24978.4]
  wire  _GEN_113; // @[Deinterleaver.scala 106:21:freechips.rocketchip.system.DefaultRV32Config.fir@24978.4]
  wire  _T_57; // @[Decoupled.scala 40:37:freechips.rocketchip.system.DefaultRV32Config.fir@24534.4]
  wire  _T_58; // @[Deinterleaver.scala 74:33:freechips.rocketchip.system.DefaultRV32Config.fir@24535.4]
  wire  _T_59; // @[Deinterleaver.scala 74:49:freechips.rocketchip.system.DefaultRV32Config.fir@24536.4]
  wire  _T_61; // @[Decoupled.scala 40:37:freechips.rocketchip.system.DefaultRV32Config.fir@24538.4]
  wire  _T_62; // @[Deinterleaver.scala 75:33:freechips.rocketchip.system.DefaultRV32Config.fir@24539.4]
  wire  _T_246_4_last; // @[Deinterleaver.scala 94:31:freechips.rocketchip.system.DefaultRV32Config.fir@24778.4 Deinterleaver.scala 94:31:freechips.rocketchip.system.DefaultRV32Config.fir@24803.4]
  wire  _T_246_3_last; // @[Deinterleaver.scala 94:31:freechips.rocketchip.system.DefaultRV32Config.fir@24778.4 Deinterleaver.scala 94:31:freechips.rocketchip.system.DefaultRV32Config.fir@24797.4]
  wire  _T_246_2_last; // @[Deinterleaver.scala 94:31:freechips.rocketchip.system.DefaultRV32Config.fir@24778.4 Deinterleaver.scala 94:31:freechips.rocketchip.system.DefaultRV32Config.fir@24791.4]
  wire  _T_246_1_last; // @[Deinterleaver.scala 94:31:freechips.rocketchip.system.DefaultRV32Config.fir@24778.4 Deinterleaver.scala 94:31:freechips.rocketchip.system.DefaultRV32Config.fir@24785.4]
  wire  _T_246_0_last; // @[Deinterleaver.scala 94:31:freechips.rocketchip.system.DefaultRV32Config.fir@24778.4 Deinterleaver.scala 94:31:freechips.rocketchip.system.DefaultRV32Config.fir@24779.4]
  wire  _GEN_13; // @[Deinterleaver.scala 95:20:freechips.rocketchip.system.DefaultRV32Config.fir@24875.4]
  wire  _GEN_19; // @[Deinterleaver.scala 95:20:freechips.rocketchip.system.DefaultRV32Config.fir@24875.4]
  wire  _GEN_25; // @[Deinterleaver.scala 95:20:freechips.rocketchip.system.DefaultRV32Config.fir@24875.4]
  wire  _GEN_31; // @[Deinterleaver.scala 95:20:freechips.rocketchip.system.DefaultRV32Config.fir@24875.4]
  wire  _GEN_37; // @[Deinterleaver.scala 95:20:freechips.rocketchip.system.DefaultRV32Config.fir@24875.4]
  wire  _GEN_43; // @[Deinterleaver.scala 95:20:freechips.rocketchip.system.DefaultRV32Config.fir@24875.4]
  wire  _GEN_49; // @[Deinterleaver.scala 95:20:freechips.rocketchip.system.DefaultRV32Config.fir@24875.4]
  wire  _GEN_55; // @[Deinterleaver.scala 95:20:freechips.rocketchip.system.DefaultRV32Config.fir@24875.4]
  wire  _GEN_61; // @[Deinterleaver.scala 95:20:freechips.rocketchip.system.DefaultRV32Config.fir@24875.4]
  wire  _GEN_67; // @[Deinterleaver.scala 95:20:freechips.rocketchip.system.DefaultRV32Config.fir@24875.4]
  wire  _GEN_73; // @[Deinterleaver.scala 95:20:freechips.rocketchip.system.DefaultRV32Config.fir@24875.4]
  wire  _GEN_79; // @[Deinterleaver.scala 95:20:freechips.rocketchip.system.DefaultRV32Config.fir@24875.4]
  wire  _GEN_85; // @[Deinterleaver.scala 95:20:freechips.rocketchip.system.DefaultRV32Config.fir@24875.4]
  wire  _GEN_91; // @[Deinterleaver.scala 95:20:freechips.rocketchip.system.DefaultRV32Config.fir@24875.4]
  wire  _GEN_97; // @[Deinterleaver.scala 95:20:freechips.rocketchip.system.DefaultRV32Config.fir@24875.4]
  wire  _T_63; // @[Deinterleaver.scala 75:48:freechips.rocketchip.system.DefaultRV32Config.fir@24540.4]
  wire [4:0] _GEN_114; // @[Deinterleaver.scala 76:27:freechips.rocketchip.system.DefaultRV32Config.fir@24541.4]
  wire [4:0] _T_65; // @[Deinterleaver.scala 76:27:freechips.rocketchip.system.DefaultRV32Config.fir@24542.4]
  wire [4:0] _GEN_115; // @[Deinterleaver.scala 76:40:freechips.rocketchip.system.DefaultRV32Config.fir@24543.4]
  wire [4:0] _T_67; // @[Deinterleaver.scala 76:40:freechips.rocketchip.system.DefaultRV32Config.fir@24544.4]
  wire  _T_68; // @[Deinterleaver.scala 79:21:freechips.rocketchip.system.DefaultRV32Config.fir@24547.4]
  wire  _T_69; // @[Deinterleaver.scala 79:35:freechips.rocketchip.system.DefaultRV32Config.fir@24548.4]
  wire  _T_70; // @[Deinterleaver.scala 79:26:freechips.rocketchip.system.DefaultRV32Config.fir@24549.4]
  wire  _T_72; // @[Deinterleaver.scala 79:20:freechips.rocketchip.system.DefaultRV32Config.fir@24551.4]
  wire  _T_73; // @[Deinterleaver.scala 79:20:freechips.rocketchip.system.DefaultRV32Config.fir@24552.4]
  wire  _T_74; // @[Deinterleaver.scala 80:21:freechips.rocketchip.system.DefaultRV32Config.fir@24557.4]
  wire  _T_75; // @[Deinterleaver.scala 80:35:freechips.rocketchip.system.DefaultRV32Config.fir@24558.4]
  wire  _T_76; // @[Deinterleaver.scala 80:26:freechips.rocketchip.system.DefaultRV32Config.fir@24559.4]
  wire  _T_78; // @[Deinterleaver.scala 80:20:freechips.rocketchip.system.DefaultRV32Config.fir@24561.4]
  wire  _T_79; // @[Deinterleaver.scala 80:20:freechips.rocketchip.system.DefaultRV32Config.fir@24562.4]
  wire  _T_80; // @[Deinterleaver.scala 81:18:freechips.rocketchip.system.DefaultRV32Config.fir@24567.4]
  reg [4:0] _T_81; // @[Deinterleaver.scala 72:32:freechips.rocketchip.system.DefaultRV32Config.fir@24568.4]
  wire  _T_85; // @[Deinterleaver.scala 74:33:freechips.rocketchip.system.DefaultRV32Config.fir@24572.4]
  wire  _T_86; // @[Deinterleaver.scala 74:49:freechips.rocketchip.system.DefaultRV32Config.fir@24573.4]
  wire  _T_89; // @[Deinterleaver.scala 75:33:freechips.rocketchip.system.DefaultRV32Config.fir@24576.4]
  wire  _T_90; // @[Deinterleaver.scala 75:48:freechips.rocketchip.system.DefaultRV32Config.fir@24577.4]
  wire [4:0] _GEN_116; // @[Deinterleaver.scala 76:27:freechips.rocketchip.system.DefaultRV32Config.fir@24578.4]
  wire [4:0] _T_92; // @[Deinterleaver.scala 76:27:freechips.rocketchip.system.DefaultRV32Config.fir@24579.4]
  wire [4:0] _GEN_117; // @[Deinterleaver.scala 76:40:freechips.rocketchip.system.DefaultRV32Config.fir@24580.4]
  wire [4:0] _T_94; // @[Deinterleaver.scala 76:40:freechips.rocketchip.system.DefaultRV32Config.fir@24581.4]
  wire  _T_95; // @[Deinterleaver.scala 79:21:freechips.rocketchip.system.DefaultRV32Config.fir@24584.4]
  wire  _T_96; // @[Deinterleaver.scala 79:35:freechips.rocketchip.system.DefaultRV32Config.fir@24585.4]
  wire  _T_97; // @[Deinterleaver.scala 79:26:freechips.rocketchip.system.DefaultRV32Config.fir@24586.4]
  wire  _T_99; // @[Deinterleaver.scala 79:20:freechips.rocketchip.system.DefaultRV32Config.fir@24588.4]
  wire  _T_100; // @[Deinterleaver.scala 79:20:freechips.rocketchip.system.DefaultRV32Config.fir@24589.4]
  wire  _T_101; // @[Deinterleaver.scala 80:21:freechips.rocketchip.system.DefaultRV32Config.fir@24594.4]
  wire  _T_102; // @[Deinterleaver.scala 80:35:freechips.rocketchip.system.DefaultRV32Config.fir@24595.4]
  wire  _T_103; // @[Deinterleaver.scala 80:26:freechips.rocketchip.system.DefaultRV32Config.fir@24596.4]
  wire  _T_105; // @[Deinterleaver.scala 80:20:freechips.rocketchip.system.DefaultRV32Config.fir@24598.4]
  wire  _T_106; // @[Deinterleaver.scala 80:20:freechips.rocketchip.system.DefaultRV32Config.fir@24599.4]
  wire  _T_107; // @[Deinterleaver.scala 81:18:freechips.rocketchip.system.DefaultRV32Config.fir@24604.4]
  reg [4:0] _T_108; // @[Deinterleaver.scala 72:32:freechips.rocketchip.system.DefaultRV32Config.fir@24605.4]
  wire  _T_112; // @[Deinterleaver.scala 74:33:freechips.rocketchip.system.DefaultRV32Config.fir@24609.4]
  wire  _T_113; // @[Deinterleaver.scala 74:49:freechips.rocketchip.system.DefaultRV32Config.fir@24610.4]
  wire  _T_116; // @[Deinterleaver.scala 75:33:freechips.rocketchip.system.DefaultRV32Config.fir@24613.4]
  wire  _T_117; // @[Deinterleaver.scala 75:48:freechips.rocketchip.system.DefaultRV32Config.fir@24614.4]
  wire [4:0] _GEN_118; // @[Deinterleaver.scala 76:27:freechips.rocketchip.system.DefaultRV32Config.fir@24615.4]
  wire [4:0] _T_119; // @[Deinterleaver.scala 76:27:freechips.rocketchip.system.DefaultRV32Config.fir@24616.4]
  wire [4:0] _GEN_119; // @[Deinterleaver.scala 76:40:freechips.rocketchip.system.DefaultRV32Config.fir@24617.4]
  wire [4:0] _T_121; // @[Deinterleaver.scala 76:40:freechips.rocketchip.system.DefaultRV32Config.fir@24618.4]
  wire  _T_122; // @[Deinterleaver.scala 79:21:freechips.rocketchip.system.DefaultRV32Config.fir@24621.4]
  wire  _T_123; // @[Deinterleaver.scala 79:35:freechips.rocketchip.system.DefaultRV32Config.fir@24622.4]
  wire  _T_124; // @[Deinterleaver.scala 79:26:freechips.rocketchip.system.DefaultRV32Config.fir@24623.4]
  wire  _T_126; // @[Deinterleaver.scala 79:20:freechips.rocketchip.system.DefaultRV32Config.fir@24625.4]
  wire  _T_127; // @[Deinterleaver.scala 79:20:freechips.rocketchip.system.DefaultRV32Config.fir@24626.4]
  wire  _T_128; // @[Deinterleaver.scala 80:21:freechips.rocketchip.system.DefaultRV32Config.fir@24631.4]
  wire  _T_129; // @[Deinterleaver.scala 80:35:freechips.rocketchip.system.DefaultRV32Config.fir@24632.4]
  wire  _T_130; // @[Deinterleaver.scala 80:26:freechips.rocketchip.system.DefaultRV32Config.fir@24633.4]
  wire  _T_132; // @[Deinterleaver.scala 80:20:freechips.rocketchip.system.DefaultRV32Config.fir@24635.4]
  wire  _T_133; // @[Deinterleaver.scala 80:20:freechips.rocketchip.system.DefaultRV32Config.fir@24636.4]
  wire  _T_134; // @[Deinterleaver.scala 81:18:freechips.rocketchip.system.DefaultRV32Config.fir@24641.4]
  reg [4:0] _T_135; // @[Deinterleaver.scala 72:32:freechips.rocketchip.system.DefaultRV32Config.fir@24642.4]
  wire  _T_139; // @[Deinterleaver.scala 74:33:freechips.rocketchip.system.DefaultRV32Config.fir@24646.4]
  wire  _T_140; // @[Deinterleaver.scala 74:49:freechips.rocketchip.system.DefaultRV32Config.fir@24647.4]
  wire  _T_143; // @[Deinterleaver.scala 75:33:freechips.rocketchip.system.DefaultRV32Config.fir@24650.4]
  wire  _T_144; // @[Deinterleaver.scala 75:48:freechips.rocketchip.system.DefaultRV32Config.fir@24651.4]
  wire [4:0] _GEN_120; // @[Deinterleaver.scala 76:27:freechips.rocketchip.system.DefaultRV32Config.fir@24652.4]
  wire [4:0] _T_146; // @[Deinterleaver.scala 76:27:freechips.rocketchip.system.DefaultRV32Config.fir@24653.4]
  wire [4:0] _GEN_121; // @[Deinterleaver.scala 76:40:freechips.rocketchip.system.DefaultRV32Config.fir@24654.4]
  wire [4:0] _T_148; // @[Deinterleaver.scala 76:40:freechips.rocketchip.system.DefaultRV32Config.fir@24655.4]
  wire  _T_149; // @[Deinterleaver.scala 79:21:freechips.rocketchip.system.DefaultRV32Config.fir@24658.4]
  wire  _T_150; // @[Deinterleaver.scala 79:35:freechips.rocketchip.system.DefaultRV32Config.fir@24659.4]
  wire  _T_151; // @[Deinterleaver.scala 79:26:freechips.rocketchip.system.DefaultRV32Config.fir@24660.4]
  wire  _T_153; // @[Deinterleaver.scala 79:20:freechips.rocketchip.system.DefaultRV32Config.fir@24662.4]
  wire  _T_154; // @[Deinterleaver.scala 79:20:freechips.rocketchip.system.DefaultRV32Config.fir@24663.4]
  wire  _T_155; // @[Deinterleaver.scala 80:21:freechips.rocketchip.system.DefaultRV32Config.fir@24668.4]
  wire  _T_156; // @[Deinterleaver.scala 80:35:freechips.rocketchip.system.DefaultRV32Config.fir@24669.4]
  wire  _T_157; // @[Deinterleaver.scala 80:26:freechips.rocketchip.system.DefaultRV32Config.fir@24670.4]
  wire  _T_159; // @[Deinterleaver.scala 80:20:freechips.rocketchip.system.DefaultRV32Config.fir@24672.4]
  wire  _T_160; // @[Deinterleaver.scala 80:20:freechips.rocketchip.system.DefaultRV32Config.fir@24673.4]
  wire  _T_161; // @[Deinterleaver.scala 81:18:freechips.rocketchip.system.DefaultRV32Config.fir@24678.4]
  reg [4:0] _T_162; // @[Deinterleaver.scala 72:32:freechips.rocketchip.system.DefaultRV32Config.fir@24679.4]
  wire  _T_166; // @[Deinterleaver.scala 74:33:freechips.rocketchip.system.DefaultRV32Config.fir@24683.4]
  wire  _T_167; // @[Deinterleaver.scala 74:49:freechips.rocketchip.system.DefaultRV32Config.fir@24684.4]
  wire  _T_170; // @[Deinterleaver.scala 75:33:freechips.rocketchip.system.DefaultRV32Config.fir@24687.4]
  wire  _T_171; // @[Deinterleaver.scala 75:48:freechips.rocketchip.system.DefaultRV32Config.fir@24688.4]
  wire [4:0] _GEN_122; // @[Deinterleaver.scala 76:27:freechips.rocketchip.system.DefaultRV32Config.fir@24689.4]
  wire [4:0] _T_173; // @[Deinterleaver.scala 76:27:freechips.rocketchip.system.DefaultRV32Config.fir@24690.4]
  wire [4:0] _GEN_123; // @[Deinterleaver.scala 76:40:freechips.rocketchip.system.DefaultRV32Config.fir@24691.4]
  wire [4:0] _T_175; // @[Deinterleaver.scala 76:40:freechips.rocketchip.system.DefaultRV32Config.fir@24692.4]
  wire  _T_176; // @[Deinterleaver.scala 79:21:freechips.rocketchip.system.DefaultRV32Config.fir@24695.4]
  wire  _T_177; // @[Deinterleaver.scala 79:35:freechips.rocketchip.system.DefaultRV32Config.fir@24696.4]
  wire  _T_178; // @[Deinterleaver.scala 79:26:freechips.rocketchip.system.DefaultRV32Config.fir@24697.4]
  wire  _T_180; // @[Deinterleaver.scala 79:20:freechips.rocketchip.system.DefaultRV32Config.fir@24699.4]
  wire  _T_181; // @[Deinterleaver.scala 79:20:freechips.rocketchip.system.DefaultRV32Config.fir@24700.4]
  wire  _T_182; // @[Deinterleaver.scala 80:21:freechips.rocketchip.system.DefaultRV32Config.fir@24705.4]
  wire  _T_183; // @[Deinterleaver.scala 80:35:freechips.rocketchip.system.DefaultRV32Config.fir@24706.4]
  wire  _T_184; // @[Deinterleaver.scala 80:26:freechips.rocketchip.system.DefaultRV32Config.fir@24707.4]
  wire  _T_186; // @[Deinterleaver.scala 80:20:freechips.rocketchip.system.DefaultRV32Config.fir@24709.4]
  wire  _T_187; // @[Deinterleaver.scala 80:20:freechips.rocketchip.system.DefaultRV32Config.fir@24710.4]
  wire  _T_188; // @[Deinterleaver.scala 81:18:freechips.rocketchip.system.DefaultRV32Config.fir@24715.4]
  wire [15:0] _T_203; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@24730.4]
  wire [16:0] _T_204; // @[package.scala 217:48:freechips.rocketchip.system.DefaultRV32Config.fir@24731.4]
  wire [15:0] _T_206; // @[package.scala 217:43:freechips.rocketchip.system.DefaultRV32Config.fir@24733.4]
  wire [17:0] _T_207; // @[package.scala 217:48:freechips.rocketchip.system.DefaultRV32Config.fir@24734.4]
  wire [15:0] _T_209; // @[package.scala 217:43:freechips.rocketchip.system.DefaultRV32Config.fir@24736.4]
  wire [19:0] _T_210; // @[package.scala 217:48:freechips.rocketchip.system.DefaultRV32Config.fir@24737.4]
  wire [15:0] _T_212; // @[package.scala 217:43:freechips.rocketchip.system.DefaultRV32Config.fir@24739.4]
  wire [23:0] _T_213; // @[package.scala 217:48:freechips.rocketchip.system.DefaultRV32Config.fir@24740.4]
  wire [15:0] _T_215; // @[package.scala 217:43:freechips.rocketchip.system.DefaultRV32Config.fir@24742.4]
  wire [16:0] _T_217; // @[Deinterleaver.scala 86:51:freechips.rocketchip.system.DefaultRV32Config.fir@24744.4]
  wire [16:0] _T_218; // @[Deinterleaver.scala 86:33:freechips.rocketchip.system.DefaultRV32Config.fir@24745.4]
  wire [16:0] _GEN_124; // @[Deinterleaver.scala 86:31:freechips.rocketchip.system.DefaultRV32Config.fir@24746.4]
  wire [16:0] _T_219; // @[Deinterleaver.scala 86:31:freechips.rocketchip.system.DefaultRV32Config.fir@24746.4]
  wire  _T_220; // @[Deinterleaver.scala 87:15:freechips.rocketchip.system.DefaultRV32Config.fir@24747.4]
  wire  _T_222; // @[Deinterleaver.scala 87:39:freechips.rocketchip.system.DefaultRV32Config.fir@24749.4]
  wire  _T_223; // @[Deinterleaver.scala 87:23:freechips.rocketchip.system.DefaultRV32Config.fir@24750.4]
  wire  _T_224; // @[Deinterleaver.scala 88:29:freechips.rocketchip.system.DefaultRV32Config.fir@24752.6]
  wire  _T_227; // @[OneHot.scala 32:14:freechips.rocketchip.system.DefaultRV32Config.fir@24756.6]
  wire [15:0] _GEN_125; // @[OneHot.scala 32:28:freechips.rocketchip.system.DefaultRV32Config.fir@24757.6]
  wire [15:0] _T_228; // @[OneHot.scala 32:28:freechips.rocketchip.system.DefaultRV32Config.fir@24757.6]
  wire  _T_231; // @[OneHot.scala 32:14:freechips.rocketchip.system.DefaultRV32Config.fir@24760.6]
  wire [7:0] _T_232; // @[OneHot.scala 32:28:freechips.rocketchip.system.DefaultRV32Config.fir@24761.6]
  wire  _T_235; // @[OneHot.scala 32:14:freechips.rocketchip.system.DefaultRV32Config.fir@24764.6]
  wire [3:0] _T_236; // @[OneHot.scala 32:28:freechips.rocketchip.system.DefaultRV32Config.fir@24765.6]
  wire  _T_239; // @[OneHot.scala 32:14:freechips.rocketchip.system.DefaultRV32Config.fir@24768.6]
  wire [1:0] _T_240; // @[OneHot.scala 32:28:freechips.rocketchip.system.DefaultRV32Config.fir@24769.6]
  wire [4:0] _T_245; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@24774.6]
  wire [4:0] _GEN_1; // @[Deinterleaver.scala 87:59:freechips.rocketchip.system.DefaultRV32Config.fir@24751.4]
  wire [3:0] _T_246_0_id; // @[Deinterleaver.scala 94:31:freechips.rocketchip.system.DefaultRV32Config.fir@24778.4 Deinterleaver.scala 94:31:freechips.rocketchip.system.DefaultRV32Config.fir@24784.4]
  wire [31:0] _T_246_0_data; // @[Deinterleaver.scala 94:31:freechips.rocketchip.system.DefaultRV32Config.fir@24778.4 Deinterleaver.scala 94:31:freechips.rocketchip.system.DefaultRV32Config.fir@24783.4]
  wire [1:0] _T_246_0_resp; // @[Deinterleaver.scala 94:31:freechips.rocketchip.system.DefaultRV32Config.fir@24778.4 Deinterleaver.scala 94:31:freechips.rocketchip.system.DefaultRV32Config.fir@24782.4]
  wire [3:0] _T_246_0_echo_tl_state_size; // @[Deinterleaver.scala 94:31:freechips.rocketchip.system.DefaultRV32Config.fir@24778.4 Deinterleaver.scala 94:31:freechips.rocketchip.system.DefaultRV32Config.fir@24781.4]
  wire [4:0] _T_246_0_echo_tl_state_source; // @[Deinterleaver.scala 94:31:freechips.rocketchip.system.DefaultRV32Config.fir@24778.4 Deinterleaver.scala 94:31:freechips.rocketchip.system.DefaultRV32Config.fir@24780.4]
  wire [3:0] _T_246_1_id; // @[Deinterleaver.scala 94:31:freechips.rocketchip.system.DefaultRV32Config.fir@24778.4 Deinterleaver.scala 94:31:freechips.rocketchip.system.DefaultRV32Config.fir@24790.4]
  wire [3:0] _GEN_8; // @[Deinterleaver.scala 95:20:freechips.rocketchip.system.DefaultRV32Config.fir@24875.4]
  wire [31:0] _T_246_1_data; // @[Deinterleaver.scala 94:31:freechips.rocketchip.system.DefaultRV32Config.fir@24778.4 Deinterleaver.scala 94:31:freechips.rocketchip.system.DefaultRV32Config.fir@24789.4]
  wire [31:0] _GEN_9; // @[Deinterleaver.scala 95:20:freechips.rocketchip.system.DefaultRV32Config.fir@24875.4]
  wire [1:0] _T_246_1_resp; // @[Deinterleaver.scala 94:31:freechips.rocketchip.system.DefaultRV32Config.fir@24778.4 Deinterleaver.scala 94:31:freechips.rocketchip.system.DefaultRV32Config.fir@24788.4]
  wire [1:0] _GEN_10; // @[Deinterleaver.scala 95:20:freechips.rocketchip.system.DefaultRV32Config.fir@24875.4]
  wire [3:0] _T_246_1_echo_tl_state_size; // @[Deinterleaver.scala 94:31:freechips.rocketchip.system.DefaultRV32Config.fir@24778.4 Deinterleaver.scala 94:31:freechips.rocketchip.system.DefaultRV32Config.fir@24787.4]
  wire [3:0] _GEN_11; // @[Deinterleaver.scala 95:20:freechips.rocketchip.system.DefaultRV32Config.fir@24875.4]
  wire [4:0] _T_246_1_echo_tl_state_source; // @[Deinterleaver.scala 94:31:freechips.rocketchip.system.DefaultRV32Config.fir@24778.4 Deinterleaver.scala 94:31:freechips.rocketchip.system.DefaultRV32Config.fir@24786.4]
  wire [4:0] _GEN_12; // @[Deinterleaver.scala 95:20:freechips.rocketchip.system.DefaultRV32Config.fir@24875.4]
  wire [3:0] _T_246_2_id; // @[Deinterleaver.scala 94:31:freechips.rocketchip.system.DefaultRV32Config.fir@24778.4 Deinterleaver.scala 94:31:freechips.rocketchip.system.DefaultRV32Config.fir@24796.4]
  wire [3:0] _GEN_14; // @[Deinterleaver.scala 95:20:freechips.rocketchip.system.DefaultRV32Config.fir@24875.4]
  wire [31:0] _T_246_2_data; // @[Deinterleaver.scala 94:31:freechips.rocketchip.system.DefaultRV32Config.fir@24778.4 Deinterleaver.scala 94:31:freechips.rocketchip.system.DefaultRV32Config.fir@24795.4]
  wire [31:0] _GEN_15; // @[Deinterleaver.scala 95:20:freechips.rocketchip.system.DefaultRV32Config.fir@24875.4]
  wire [1:0] _T_246_2_resp; // @[Deinterleaver.scala 94:31:freechips.rocketchip.system.DefaultRV32Config.fir@24778.4 Deinterleaver.scala 94:31:freechips.rocketchip.system.DefaultRV32Config.fir@24794.4]
  wire [1:0] _GEN_16; // @[Deinterleaver.scala 95:20:freechips.rocketchip.system.DefaultRV32Config.fir@24875.4]
  wire [3:0] _T_246_2_echo_tl_state_size; // @[Deinterleaver.scala 94:31:freechips.rocketchip.system.DefaultRV32Config.fir@24778.4 Deinterleaver.scala 94:31:freechips.rocketchip.system.DefaultRV32Config.fir@24793.4]
  wire [3:0] _GEN_17; // @[Deinterleaver.scala 95:20:freechips.rocketchip.system.DefaultRV32Config.fir@24875.4]
  wire [4:0] _T_246_2_echo_tl_state_source; // @[Deinterleaver.scala 94:31:freechips.rocketchip.system.DefaultRV32Config.fir@24778.4 Deinterleaver.scala 94:31:freechips.rocketchip.system.DefaultRV32Config.fir@24792.4]
  wire [4:0] _GEN_18; // @[Deinterleaver.scala 95:20:freechips.rocketchip.system.DefaultRV32Config.fir@24875.4]
  wire [3:0] _T_246_3_id; // @[Deinterleaver.scala 94:31:freechips.rocketchip.system.DefaultRV32Config.fir@24778.4 Deinterleaver.scala 94:31:freechips.rocketchip.system.DefaultRV32Config.fir@24802.4]
  wire [3:0] _GEN_20; // @[Deinterleaver.scala 95:20:freechips.rocketchip.system.DefaultRV32Config.fir@24875.4]
  wire [31:0] _T_246_3_data; // @[Deinterleaver.scala 94:31:freechips.rocketchip.system.DefaultRV32Config.fir@24778.4 Deinterleaver.scala 94:31:freechips.rocketchip.system.DefaultRV32Config.fir@24801.4]
  wire [31:0] _GEN_21; // @[Deinterleaver.scala 95:20:freechips.rocketchip.system.DefaultRV32Config.fir@24875.4]
  wire [1:0] _T_246_3_resp; // @[Deinterleaver.scala 94:31:freechips.rocketchip.system.DefaultRV32Config.fir@24778.4 Deinterleaver.scala 94:31:freechips.rocketchip.system.DefaultRV32Config.fir@24800.4]
  wire [1:0] _GEN_22; // @[Deinterleaver.scala 95:20:freechips.rocketchip.system.DefaultRV32Config.fir@24875.4]
  wire [3:0] _T_246_3_echo_tl_state_size; // @[Deinterleaver.scala 94:31:freechips.rocketchip.system.DefaultRV32Config.fir@24778.4 Deinterleaver.scala 94:31:freechips.rocketchip.system.DefaultRV32Config.fir@24799.4]
  wire [3:0] _GEN_23; // @[Deinterleaver.scala 95:20:freechips.rocketchip.system.DefaultRV32Config.fir@24875.4]
  wire [4:0] _T_246_3_echo_tl_state_source; // @[Deinterleaver.scala 94:31:freechips.rocketchip.system.DefaultRV32Config.fir@24778.4 Deinterleaver.scala 94:31:freechips.rocketchip.system.DefaultRV32Config.fir@24798.4]
  wire [4:0] _GEN_24; // @[Deinterleaver.scala 95:20:freechips.rocketchip.system.DefaultRV32Config.fir@24875.4]
  wire [3:0] _T_246_4_id; // @[Deinterleaver.scala 94:31:freechips.rocketchip.system.DefaultRV32Config.fir@24778.4 Deinterleaver.scala 94:31:freechips.rocketchip.system.DefaultRV32Config.fir@24808.4]
  wire [3:0] _GEN_26; // @[Deinterleaver.scala 95:20:freechips.rocketchip.system.DefaultRV32Config.fir@24875.4]
  wire [31:0] _T_246_4_data; // @[Deinterleaver.scala 94:31:freechips.rocketchip.system.DefaultRV32Config.fir@24778.4 Deinterleaver.scala 94:31:freechips.rocketchip.system.DefaultRV32Config.fir@24807.4]
  wire [31:0] _GEN_27; // @[Deinterleaver.scala 95:20:freechips.rocketchip.system.DefaultRV32Config.fir@24875.4]
  wire [1:0] _T_246_4_resp; // @[Deinterleaver.scala 94:31:freechips.rocketchip.system.DefaultRV32Config.fir@24778.4 Deinterleaver.scala 94:31:freechips.rocketchip.system.DefaultRV32Config.fir@24806.4]
  wire [1:0] _GEN_28; // @[Deinterleaver.scala 95:20:freechips.rocketchip.system.DefaultRV32Config.fir@24875.4]
  wire [3:0] _T_246_4_echo_tl_state_size; // @[Deinterleaver.scala 94:31:freechips.rocketchip.system.DefaultRV32Config.fir@24778.4 Deinterleaver.scala 94:31:freechips.rocketchip.system.DefaultRV32Config.fir@24805.4]
  wire [3:0] _GEN_29; // @[Deinterleaver.scala 95:20:freechips.rocketchip.system.DefaultRV32Config.fir@24875.4]
  wire [4:0] _T_246_4_echo_tl_state_source; // @[Deinterleaver.scala 94:31:freechips.rocketchip.system.DefaultRV32Config.fir@24778.4 Deinterleaver.scala 94:31:freechips.rocketchip.system.DefaultRV32Config.fir@24804.4]
  wire [4:0] _GEN_30; // @[Deinterleaver.scala 95:20:freechips.rocketchip.system.DefaultRV32Config.fir@24875.4]
  wire [3:0] _GEN_32; // @[Deinterleaver.scala 95:20:freechips.rocketchip.system.DefaultRV32Config.fir@24875.4]
  wire [31:0] _GEN_33; // @[Deinterleaver.scala 95:20:freechips.rocketchip.system.DefaultRV32Config.fir@24875.4]
  wire [1:0] _GEN_34; // @[Deinterleaver.scala 95:20:freechips.rocketchip.system.DefaultRV32Config.fir@24875.4]
  wire [3:0] _GEN_35; // @[Deinterleaver.scala 95:20:freechips.rocketchip.system.DefaultRV32Config.fir@24875.4]
  wire [4:0] _GEN_36; // @[Deinterleaver.scala 95:20:freechips.rocketchip.system.DefaultRV32Config.fir@24875.4]
  wire [3:0] _GEN_38; // @[Deinterleaver.scala 95:20:freechips.rocketchip.system.DefaultRV32Config.fir@24875.4]
  wire [31:0] _GEN_39; // @[Deinterleaver.scala 95:20:freechips.rocketchip.system.DefaultRV32Config.fir@24875.4]
  wire [1:0] _GEN_40; // @[Deinterleaver.scala 95:20:freechips.rocketchip.system.DefaultRV32Config.fir@24875.4]
  wire [3:0] _GEN_41; // @[Deinterleaver.scala 95:20:freechips.rocketchip.system.DefaultRV32Config.fir@24875.4]
  wire [4:0] _GEN_42; // @[Deinterleaver.scala 95:20:freechips.rocketchip.system.DefaultRV32Config.fir@24875.4]
  wire [3:0] _GEN_44; // @[Deinterleaver.scala 95:20:freechips.rocketchip.system.DefaultRV32Config.fir@24875.4]
  wire [31:0] _GEN_45; // @[Deinterleaver.scala 95:20:freechips.rocketchip.system.DefaultRV32Config.fir@24875.4]
  wire [1:0] _GEN_46; // @[Deinterleaver.scala 95:20:freechips.rocketchip.system.DefaultRV32Config.fir@24875.4]
  wire [3:0] _GEN_47; // @[Deinterleaver.scala 95:20:freechips.rocketchip.system.DefaultRV32Config.fir@24875.4]
  wire [4:0] _GEN_48; // @[Deinterleaver.scala 95:20:freechips.rocketchip.system.DefaultRV32Config.fir@24875.4]
  wire [3:0] _GEN_50; // @[Deinterleaver.scala 95:20:freechips.rocketchip.system.DefaultRV32Config.fir@24875.4]
  wire [31:0] _GEN_51; // @[Deinterleaver.scala 95:20:freechips.rocketchip.system.DefaultRV32Config.fir@24875.4]
  wire [1:0] _GEN_52; // @[Deinterleaver.scala 95:20:freechips.rocketchip.system.DefaultRV32Config.fir@24875.4]
  wire [3:0] _GEN_53; // @[Deinterleaver.scala 95:20:freechips.rocketchip.system.DefaultRV32Config.fir@24875.4]
  wire [4:0] _GEN_54; // @[Deinterleaver.scala 95:20:freechips.rocketchip.system.DefaultRV32Config.fir@24875.4]
  wire [3:0] _GEN_56; // @[Deinterleaver.scala 95:20:freechips.rocketchip.system.DefaultRV32Config.fir@24875.4]
  wire [31:0] _GEN_57; // @[Deinterleaver.scala 95:20:freechips.rocketchip.system.DefaultRV32Config.fir@24875.4]
  wire [1:0] _GEN_58; // @[Deinterleaver.scala 95:20:freechips.rocketchip.system.DefaultRV32Config.fir@24875.4]
  wire [3:0] _GEN_59; // @[Deinterleaver.scala 95:20:freechips.rocketchip.system.DefaultRV32Config.fir@24875.4]
  wire [4:0] _GEN_60; // @[Deinterleaver.scala 95:20:freechips.rocketchip.system.DefaultRV32Config.fir@24875.4]
  wire [3:0] _GEN_62; // @[Deinterleaver.scala 95:20:freechips.rocketchip.system.DefaultRV32Config.fir@24875.4]
  wire [31:0] _GEN_63; // @[Deinterleaver.scala 95:20:freechips.rocketchip.system.DefaultRV32Config.fir@24875.4]
  wire [1:0] _GEN_64; // @[Deinterleaver.scala 95:20:freechips.rocketchip.system.DefaultRV32Config.fir@24875.4]
  wire [3:0] _GEN_65; // @[Deinterleaver.scala 95:20:freechips.rocketchip.system.DefaultRV32Config.fir@24875.4]
  wire [4:0] _GEN_66; // @[Deinterleaver.scala 95:20:freechips.rocketchip.system.DefaultRV32Config.fir@24875.4]
  wire [3:0] _GEN_68; // @[Deinterleaver.scala 95:20:freechips.rocketchip.system.DefaultRV32Config.fir@24875.4]
  wire [31:0] _GEN_69; // @[Deinterleaver.scala 95:20:freechips.rocketchip.system.DefaultRV32Config.fir@24875.4]
  wire [1:0] _GEN_70; // @[Deinterleaver.scala 95:20:freechips.rocketchip.system.DefaultRV32Config.fir@24875.4]
  wire [3:0] _GEN_71; // @[Deinterleaver.scala 95:20:freechips.rocketchip.system.DefaultRV32Config.fir@24875.4]
  wire [4:0] _GEN_72; // @[Deinterleaver.scala 95:20:freechips.rocketchip.system.DefaultRV32Config.fir@24875.4]
  wire [3:0] _GEN_74; // @[Deinterleaver.scala 95:20:freechips.rocketchip.system.DefaultRV32Config.fir@24875.4]
  wire [31:0] _GEN_75; // @[Deinterleaver.scala 95:20:freechips.rocketchip.system.DefaultRV32Config.fir@24875.4]
  wire [1:0] _GEN_76; // @[Deinterleaver.scala 95:20:freechips.rocketchip.system.DefaultRV32Config.fir@24875.4]
  wire [3:0] _GEN_77; // @[Deinterleaver.scala 95:20:freechips.rocketchip.system.DefaultRV32Config.fir@24875.4]
  wire [4:0] _GEN_78; // @[Deinterleaver.scala 95:20:freechips.rocketchip.system.DefaultRV32Config.fir@24875.4]
  wire [3:0] _GEN_80; // @[Deinterleaver.scala 95:20:freechips.rocketchip.system.DefaultRV32Config.fir@24875.4]
  wire [31:0] _GEN_81; // @[Deinterleaver.scala 95:20:freechips.rocketchip.system.DefaultRV32Config.fir@24875.4]
  wire [1:0] _GEN_82; // @[Deinterleaver.scala 95:20:freechips.rocketchip.system.DefaultRV32Config.fir@24875.4]
  wire [3:0] _GEN_83; // @[Deinterleaver.scala 95:20:freechips.rocketchip.system.DefaultRV32Config.fir@24875.4]
  wire [4:0] _GEN_84; // @[Deinterleaver.scala 95:20:freechips.rocketchip.system.DefaultRV32Config.fir@24875.4]
  wire [3:0] _GEN_86; // @[Deinterleaver.scala 95:20:freechips.rocketchip.system.DefaultRV32Config.fir@24875.4]
  wire [31:0] _GEN_87; // @[Deinterleaver.scala 95:20:freechips.rocketchip.system.DefaultRV32Config.fir@24875.4]
  wire [1:0] _GEN_88; // @[Deinterleaver.scala 95:20:freechips.rocketchip.system.DefaultRV32Config.fir@24875.4]
  wire [3:0] _GEN_89; // @[Deinterleaver.scala 95:20:freechips.rocketchip.system.DefaultRV32Config.fir@24875.4]
  wire [4:0] _GEN_90; // @[Deinterleaver.scala 95:20:freechips.rocketchip.system.DefaultRV32Config.fir@24875.4]
  Queue_5 queue_0 ( // @[Deinterleaver.scala 44:27:freechips.rocketchip.system.DefaultRV32Config.fir@24222.4]
    .clock(queue_0_clock),
    .reset(queue_0_reset),
    .io_enq_ready(queue_0_io_enq_ready),
    .io_enq_valid(queue_0_io_enq_valid),
    .io_enq_bits_id(queue_0_io_enq_bits_id),
    .io_enq_bits_data(queue_0_io_enq_bits_data),
    .io_enq_bits_resp(queue_0_io_enq_bits_resp),
    .io_enq_bits_echo_tl_state_size(queue_0_io_enq_bits_echo_tl_state_size),
    .io_enq_bits_echo_tl_state_source(queue_0_io_enq_bits_echo_tl_state_source),
    .io_enq_bits_last(queue_0_io_enq_bits_last),
    .io_deq_ready(queue_0_io_deq_ready),
    .io_deq_valid(queue_0_io_deq_valid),
    .io_deq_bits_id(queue_0_io_deq_bits_id),
    .io_deq_bits_data(queue_0_io_deq_bits_data),
    .io_deq_bits_resp(queue_0_io_deq_bits_resp),
    .io_deq_bits_echo_tl_state_size(queue_0_io_deq_bits_echo_tl_state_size),
    .io_deq_bits_echo_tl_state_source(queue_0_io_deq_bits_echo_tl_state_source),
    .io_deq_bits_last(queue_0_io_deq_bits_last)
  );
  Queue_5 queue_1 ( // @[Deinterleaver.scala 44:27:freechips.rocketchip.system.DefaultRV32Config.fir@24225.4]
    .clock(queue_1_clock),
    .reset(queue_1_reset),
    .io_enq_ready(queue_1_io_enq_ready),
    .io_enq_valid(queue_1_io_enq_valid),
    .io_enq_bits_id(queue_1_io_enq_bits_id),
    .io_enq_bits_data(queue_1_io_enq_bits_data),
    .io_enq_bits_resp(queue_1_io_enq_bits_resp),
    .io_enq_bits_echo_tl_state_size(queue_1_io_enq_bits_echo_tl_state_size),
    .io_enq_bits_echo_tl_state_source(queue_1_io_enq_bits_echo_tl_state_source),
    .io_enq_bits_last(queue_1_io_enq_bits_last),
    .io_deq_ready(queue_1_io_deq_ready),
    .io_deq_valid(queue_1_io_deq_valid),
    .io_deq_bits_id(queue_1_io_deq_bits_id),
    .io_deq_bits_data(queue_1_io_deq_bits_data),
    .io_deq_bits_resp(queue_1_io_deq_bits_resp),
    .io_deq_bits_echo_tl_state_size(queue_1_io_deq_bits_echo_tl_state_size),
    .io_deq_bits_echo_tl_state_source(queue_1_io_deq_bits_echo_tl_state_source),
    .io_deq_bits_last(queue_1_io_deq_bits_last)
  );
  Queue_5 queue_2 ( // @[Deinterleaver.scala 44:27:freechips.rocketchip.system.DefaultRV32Config.fir@24228.4]
    .clock(queue_2_clock),
    .reset(queue_2_reset),
    .io_enq_ready(queue_2_io_enq_ready),
    .io_enq_valid(queue_2_io_enq_valid),
    .io_enq_bits_id(queue_2_io_enq_bits_id),
    .io_enq_bits_data(queue_2_io_enq_bits_data),
    .io_enq_bits_resp(queue_2_io_enq_bits_resp),
    .io_enq_bits_echo_tl_state_size(queue_2_io_enq_bits_echo_tl_state_size),
    .io_enq_bits_echo_tl_state_source(queue_2_io_enq_bits_echo_tl_state_source),
    .io_enq_bits_last(queue_2_io_enq_bits_last),
    .io_deq_ready(queue_2_io_deq_ready),
    .io_deq_valid(queue_2_io_deq_valid),
    .io_deq_bits_id(queue_2_io_deq_bits_id),
    .io_deq_bits_data(queue_2_io_deq_bits_data),
    .io_deq_bits_resp(queue_2_io_deq_bits_resp),
    .io_deq_bits_echo_tl_state_size(queue_2_io_deq_bits_echo_tl_state_size),
    .io_deq_bits_echo_tl_state_source(queue_2_io_deq_bits_echo_tl_state_source),
    .io_deq_bits_last(queue_2_io_deq_bits_last)
  );
  Queue_5 queue_3 ( // @[Deinterleaver.scala 44:27:freechips.rocketchip.system.DefaultRV32Config.fir@24231.4]
    .clock(queue_3_clock),
    .reset(queue_3_reset),
    .io_enq_ready(queue_3_io_enq_ready),
    .io_enq_valid(queue_3_io_enq_valid),
    .io_enq_bits_id(queue_3_io_enq_bits_id),
    .io_enq_bits_data(queue_3_io_enq_bits_data),
    .io_enq_bits_resp(queue_3_io_enq_bits_resp),
    .io_enq_bits_echo_tl_state_size(queue_3_io_enq_bits_echo_tl_state_size),
    .io_enq_bits_echo_tl_state_source(queue_3_io_enq_bits_echo_tl_state_source),
    .io_enq_bits_last(queue_3_io_enq_bits_last),
    .io_deq_ready(queue_3_io_deq_ready),
    .io_deq_valid(queue_3_io_deq_valid),
    .io_deq_bits_id(queue_3_io_deq_bits_id),
    .io_deq_bits_data(queue_3_io_deq_bits_data),
    .io_deq_bits_resp(queue_3_io_deq_bits_resp),
    .io_deq_bits_echo_tl_state_size(queue_3_io_deq_bits_echo_tl_state_size),
    .io_deq_bits_echo_tl_state_source(queue_3_io_deq_bits_echo_tl_state_source),
    .io_deq_bits_last(queue_3_io_deq_bits_last)
  );
  Queue_5 queue_4 ( // @[Deinterleaver.scala 44:27:freechips.rocketchip.system.DefaultRV32Config.fir@24234.4]
    .clock(queue_4_clock),
    .reset(queue_4_reset),
    .io_enq_ready(queue_4_io_enq_ready),
    .io_enq_valid(queue_4_io_enq_valid),
    .io_enq_bits_id(queue_4_io_enq_bits_id),
    .io_enq_bits_data(queue_4_io_enq_bits_data),
    .io_enq_bits_resp(queue_4_io_enq_bits_resp),
    .io_enq_bits_echo_tl_state_size(queue_4_io_enq_bits_echo_tl_state_size),
    .io_enq_bits_echo_tl_state_source(queue_4_io_enq_bits_echo_tl_state_source),
    .io_enq_bits_last(queue_4_io_enq_bits_last),
    .io_deq_ready(queue_4_io_deq_ready),
    .io_deq_valid(queue_4_io_deq_valid),
    .io_deq_bits_id(queue_4_io_deq_bits_id),
    .io_deq_bits_data(queue_4_io_deq_bits_data),
    .io_deq_bits_resp(queue_4_io_deq_bits_resp),
    .io_deq_bits_echo_tl_state_size(queue_4_io_deq_bits_echo_tl_state_size),
    .io_deq_bits_echo_tl_state_source(queue_4_io_deq_bits_echo_tl_state_source),
    .io_deq_bits_last(queue_4_io_deq_bits_last)
  );
  assign _T_52 = 16'h1 << auto_out_r_bits_id; // @[OneHot.scala 65:12:freechips.rocketchip.system.DefaultRV32Config.fir@24529.4]
  assign queue_wire_5_enq_valid = _T_52[5] & auto_out_r_valid; // @[Deinterleaver.scala 108:28:freechips.rocketchip.system.DefaultRV32Config.fir@25019.4]
  assign _T_2 = ~queue_wire_5_enq_valid; // @[Deinterleaver.scala 53:20:freechips.rocketchip.system.DefaultRV32Config.fir@24238.4]
  assign _T_4 = _T_2 | reset; // @[Deinterleaver.scala 53:19:freechips.rocketchip.system.DefaultRV32Config.fir@24240.4]
  assign _T_5 = ~_T_4; // @[Deinterleaver.scala 53:19:freechips.rocketchip.system.DefaultRV32Config.fir@24241.4]
  assign queue_wire_6_enq_valid = _T_52[6] & auto_out_r_valid; // @[Deinterleaver.scala 108:28:freechips.rocketchip.system.DefaultRV32Config.fir@25027.4]
  assign _T_6 = ~queue_wire_6_enq_valid; // @[Deinterleaver.scala 53:20:freechips.rocketchip.system.DefaultRV32Config.fir@24264.4]
  assign _T_8 = _T_6 | reset; // @[Deinterleaver.scala 53:19:freechips.rocketchip.system.DefaultRV32Config.fir@24266.4]
  assign _T_9 = ~_T_8; // @[Deinterleaver.scala 53:19:freechips.rocketchip.system.DefaultRV32Config.fir@24267.4]
  assign queue_wire_7_enq_valid = _T_52[7] & auto_out_r_valid; // @[Deinterleaver.scala 108:28:freechips.rocketchip.system.DefaultRV32Config.fir@25035.4]
  assign _T_10 = ~queue_wire_7_enq_valid; // @[Deinterleaver.scala 53:20:freechips.rocketchip.system.DefaultRV32Config.fir@24290.4]
  assign _T_12 = _T_10 | reset; // @[Deinterleaver.scala 53:19:freechips.rocketchip.system.DefaultRV32Config.fir@24292.4]
  assign _T_13 = ~_T_12; // @[Deinterleaver.scala 53:19:freechips.rocketchip.system.DefaultRV32Config.fir@24293.4]
  assign queue_wire_8_enq_valid = _T_52[8] & auto_out_r_valid; // @[Deinterleaver.scala 108:28:freechips.rocketchip.system.DefaultRV32Config.fir@25043.4]
  assign _T_14 = ~queue_wire_8_enq_valid; // @[Deinterleaver.scala 53:20:freechips.rocketchip.system.DefaultRV32Config.fir@24316.4]
  assign _T_16 = _T_14 | reset; // @[Deinterleaver.scala 53:19:freechips.rocketchip.system.DefaultRV32Config.fir@24318.4]
  assign _T_17 = ~_T_16; // @[Deinterleaver.scala 53:19:freechips.rocketchip.system.DefaultRV32Config.fir@24319.4]
  assign queue_wire_9_enq_valid = _T_52[9] & auto_out_r_valid; // @[Deinterleaver.scala 108:28:freechips.rocketchip.system.DefaultRV32Config.fir@25051.4]
  assign _T_18 = ~queue_wire_9_enq_valid; // @[Deinterleaver.scala 53:20:freechips.rocketchip.system.DefaultRV32Config.fir@24342.4]
  assign _T_20 = _T_18 | reset; // @[Deinterleaver.scala 53:19:freechips.rocketchip.system.DefaultRV32Config.fir@24344.4]
  assign _T_21 = ~_T_20; // @[Deinterleaver.scala 53:19:freechips.rocketchip.system.DefaultRV32Config.fir@24345.4]
  assign queue_wire_10_enq_valid = _T_52[10] & auto_out_r_valid; // @[Deinterleaver.scala 108:28:freechips.rocketchip.system.DefaultRV32Config.fir@25059.4]
  assign _T_22 = ~queue_wire_10_enq_valid; // @[Deinterleaver.scala 53:20:freechips.rocketchip.system.DefaultRV32Config.fir@24368.4]
  assign _T_24 = _T_22 | reset; // @[Deinterleaver.scala 53:19:freechips.rocketchip.system.DefaultRV32Config.fir@24370.4]
  assign _T_25 = ~_T_24; // @[Deinterleaver.scala 53:19:freechips.rocketchip.system.DefaultRV32Config.fir@24371.4]
  assign queue_wire_11_enq_valid = _T_52[11] & auto_out_r_valid; // @[Deinterleaver.scala 108:28:freechips.rocketchip.system.DefaultRV32Config.fir@25067.4]
  assign _T_26 = ~queue_wire_11_enq_valid; // @[Deinterleaver.scala 53:20:freechips.rocketchip.system.DefaultRV32Config.fir@24394.4]
  assign _T_28 = _T_26 | reset; // @[Deinterleaver.scala 53:19:freechips.rocketchip.system.DefaultRV32Config.fir@24396.4]
  assign _T_29 = ~_T_28; // @[Deinterleaver.scala 53:19:freechips.rocketchip.system.DefaultRV32Config.fir@24397.4]
  assign queue_wire_12_enq_valid = _T_52[12] & auto_out_r_valid; // @[Deinterleaver.scala 108:28:freechips.rocketchip.system.DefaultRV32Config.fir@25075.4]
  assign _T_30 = ~queue_wire_12_enq_valid; // @[Deinterleaver.scala 53:20:freechips.rocketchip.system.DefaultRV32Config.fir@24420.4]
  assign _T_32 = _T_30 | reset; // @[Deinterleaver.scala 53:19:freechips.rocketchip.system.DefaultRV32Config.fir@24422.4]
  assign _T_33 = ~_T_32; // @[Deinterleaver.scala 53:19:freechips.rocketchip.system.DefaultRV32Config.fir@24423.4]
  assign queue_wire_13_enq_valid = _T_52[13] & auto_out_r_valid; // @[Deinterleaver.scala 108:28:freechips.rocketchip.system.DefaultRV32Config.fir@25083.4]
  assign _T_34 = ~queue_wire_13_enq_valid; // @[Deinterleaver.scala 53:20:freechips.rocketchip.system.DefaultRV32Config.fir@24446.4]
  assign _T_36 = _T_34 | reset; // @[Deinterleaver.scala 53:19:freechips.rocketchip.system.DefaultRV32Config.fir@24448.4]
  assign _T_37 = ~_T_36; // @[Deinterleaver.scala 53:19:freechips.rocketchip.system.DefaultRV32Config.fir@24449.4]
  assign queue_wire_14_enq_valid = _T_52[14] & auto_out_r_valid; // @[Deinterleaver.scala 108:28:freechips.rocketchip.system.DefaultRV32Config.fir@25091.4]
  assign _T_38 = ~queue_wire_14_enq_valid; // @[Deinterleaver.scala 53:20:freechips.rocketchip.system.DefaultRV32Config.fir@24472.4]
  assign _T_40 = _T_38 | reset; // @[Deinterleaver.scala 53:19:freechips.rocketchip.system.DefaultRV32Config.fir@24474.4]
  assign _T_41 = ~_T_40; // @[Deinterleaver.scala 53:19:freechips.rocketchip.system.DefaultRV32Config.fir@24475.4]
  assign queue_wire_15_enq_valid = _T_52[15] & auto_out_r_valid; // @[Deinterleaver.scala 108:28:freechips.rocketchip.system.DefaultRV32Config.fir@25099.4]
  assign _T_42 = ~queue_wire_15_enq_valid; // @[Deinterleaver.scala 53:20:freechips.rocketchip.system.DefaultRV32Config.fir@24498.4]
  assign _T_44 = _T_42 | reset; // @[Deinterleaver.scala 53:19:freechips.rocketchip.system.DefaultRV32Config.fir@24500.4]
  assign _T_45 = ~_T_44; // @[Deinterleaver.scala 53:19:freechips.rocketchip.system.DefaultRV32Config.fir@24501.4]
  assign _T_49 = 16'h1 << _T_47; // @[OneHot.scala 65:12:freechips.rocketchip.system.DefaultRV32Config.fir@24526.4]
  assign _T_311_4 = queue_4_io_enq_ready; // @[Deinterleaver.scala 105:33:freechips.rocketchip.system.DefaultRV32Config.fir@24961.4 Deinterleaver.scala 105:33:freechips.rocketchip.system.DefaultRV32Config.fir@24966.4]
  assign _T_311_3 = queue_3_io_enq_ready; // @[Deinterleaver.scala 105:33:freechips.rocketchip.system.DefaultRV32Config.fir@24961.4 Deinterleaver.scala 105:33:freechips.rocketchip.system.DefaultRV32Config.fir@24965.4]
  assign _T_311_2 = queue_2_io_enq_ready; // @[Deinterleaver.scala 105:33:freechips.rocketchip.system.DefaultRV32Config.fir@24961.4 Deinterleaver.scala 105:33:freechips.rocketchip.system.DefaultRV32Config.fir@24964.4]
  assign _T_311_1 = queue_1_io_enq_ready; // @[Deinterleaver.scala 105:33:freechips.rocketchip.system.DefaultRV32Config.fir@24961.4 Deinterleaver.scala 105:33:freechips.rocketchip.system.DefaultRV32Config.fir@24963.4]
  assign _T_311_0 = queue_0_io_enq_ready; // @[Deinterleaver.scala 105:33:freechips.rocketchip.system.DefaultRV32Config.fir@24961.4 Deinterleaver.scala 105:33:freechips.rocketchip.system.DefaultRV32Config.fir@24962.4]
  assign _GEN_99 = 4'h1 == auto_out_r_bits_id ? _T_311_1 : _T_311_0; // @[Deinterleaver.scala 106:21:freechips.rocketchip.system.DefaultRV32Config.fir@24978.4]
  assign _GEN_100 = 4'h2 == auto_out_r_bits_id ? _T_311_2 : _GEN_99; // @[Deinterleaver.scala 106:21:freechips.rocketchip.system.DefaultRV32Config.fir@24978.4]
  assign _GEN_101 = 4'h3 == auto_out_r_bits_id ? _T_311_3 : _GEN_100; // @[Deinterleaver.scala 106:21:freechips.rocketchip.system.DefaultRV32Config.fir@24978.4]
  assign _GEN_102 = 4'h4 == auto_out_r_bits_id ? _T_311_4 : _GEN_101; // @[Deinterleaver.scala 106:21:freechips.rocketchip.system.DefaultRV32Config.fir@24978.4]
  assign _GEN_103 = 4'h5 == auto_out_r_bits_id ? 1'h0 : _GEN_102; // @[Deinterleaver.scala 106:21:freechips.rocketchip.system.DefaultRV32Config.fir@24978.4]
  assign _GEN_104 = 4'h6 == auto_out_r_bits_id ? 1'h0 : _GEN_103; // @[Deinterleaver.scala 106:21:freechips.rocketchip.system.DefaultRV32Config.fir@24978.4]
  assign _GEN_105 = 4'h7 == auto_out_r_bits_id ? 1'h0 : _GEN_104; // @[Deinterleaver.scala 106:21:freechips.rocketchip.system.DefaultRV32Config.fir@24978.4]
  assign _GEN_106 = 4'h8 == auto_out_r_bits_id ? 1'h0 : _GEN_105; // @[Deinterleaver.scala 106:21:freechips.rocketchip.system.DefaultRV32Config.fir@24978.4]
  assign _GEN_107 = 4'h9 == auto_out_r_bits_id ? 1'h0 : _GEN_106; // @[Deinterleaver.scala 106:21:freechips.rocketchip.system.DefaultRV32Config.fir@24978.4]
  assign _GEN_108 = 4'ha == auto_out_r_bits_id ? 1'h0 : _GEN_107; // @[Deinterleaver.scala 106:21:freechips.rocketchip.system.DefaultRV32Config.fir@24978.4]
  assign _GEN_109 = 4'hb == auto_out_r_bits_id ? 1'h0 : _GEN_108; // @[Deinterleaver.scala 106:21:freechips.rocketchip.system.DefaultRV32Config.fir@24978.4]
  assign _GEN_110 = 4'hc == auto_out_r_bits_id ? 1'h0 : _GEN_109; // @[Deinterleaver.scala 106:21:freechips.rocketchip.system.DefaultRV32Config.fir@24978.4]
  assign _GEN_111 = 4'hd == auto_out_r_bits_id ? 1'h0 : _GEN_110; // @[Deinterleaver.scala 106:21:freechips.rocketchip.system.DefaultRV32Config.fir@24978.4]
  assign _GEN_112 = 4'he == auto_out_r_bits_id ? 1'h0 : _GEN_111; // @[Deinterleaver.scala 106:21:freechips.rocketchip.system.DefaultRV32Config.fir@24978.4]
  assign _GEN_113 = 4'hf == auto_out_r_bits_id ? 1'h0 : _GEN_112; // @[Deinterleaver.scala 106:21:freechips.rocketchip.system.DefaultRV32Config.fir@24978.4]
  assign _T_57 = _GEN_113 & auto_out_r_valid; // @[Decoupled.scala 40:37:freechips.rocketchip.system.DefaultRV32Config.fir@24534.4]
  assign _T_58 = _T_52[0] & _T_57; // @[Deinterleaver.scala 74:33:freechips.rocketchip.system.DefaultRV32Config.fir@24535.4]
  assign _T_59 = _T_58 & auto_out_r_bits_last; // @[Deinterleaver.scala 74:49:freechips.rocketchip.system.DefaultRV32Config.fir@24536.4]
  assign _T_61 = auto_in_r_ready & _T_46; // @[Decoupled.scala 40:37:freechips.rocketchip.system.DefaultRV32Config.fir@24538.4]
  assign _T_62 = _T_49[0] & _T_61; // @[Deinterleaver.scala 75:33:freechips.rocketchip.system.DefaultRV32Config.fir@24539.4]
  assign _T_246_4_last = queue_4_io_deq_bits_last; // @[Deinterleaver.scala 94:31:freechips.rocketchip.system.DefaultRV32Config.fir@24778.4 Deinterleaver.scala 94:31:freechips.rocketchip.system.DefaultRV32Config.fir@24803.4]
  assign _T_246_3_last = queue_3_io_deq_bits_last; // @[Deinterleaver.scala 94:31:freechips.rocketchip.system.DefaultRV32Config.fir@24778.4 Deinterleaver.scala 94:31:freechips.rocketchip.system.DefaultRV32Config.fir@24797.4]
  assign _T_246_2_last = queue_2_io_deq_bits_last; // @[Deinterleaver.scala 94:31:freechips.rocketchip.system.DefaultRV32Config.fir@24778.4 Deinterleaver.scala 94:31:freechips.rocketchip.system.DefaultRV32Config.fir@24791.4]
  assign _T_246_1_last = queue_1_io_deq_bits_last; // @[Deinterleaver.scala 94:31:freechips.rocketchip.system.DefaultRV32Config.fir@24778.4 Deinterleaver.scala 94:31:freechips.rocketchip.system.DefaultRV32Config.fir@24785.4]
  assign _T_246_0_last = queue_0_io_deq_bits_last; // @[Deinterleaver.scala 94:31:freechips.rocketchip.system.DefaultRV32Config.fir@24778.4 Deinterleaver.scala 94:31:freechips.rocketchip.system.DefaultRV32Config.fir@24779.4]
  assign _GEN_13 = 4'h1 == _T_47 ? _T_246_1_last : _T_246_0_last; // @[Deinterleaver.scala 95:20:freechips.rocketchip.system.DefaultRV32Config.fir@24875.4]
  assign _GEN_19 = 4'h2 == _T_47 ? _T_246_2_last : _GEN_13; // @[Deinterleaver.scala 95:20:freechips.rocketchip.system.DefaultRV32Config.fir@24875.4]
  assign _GEN_25 = 4'h3 == _T_47 ? _T_246_3_last : _GEN_19; // @[Deinterleaver.scala 95:20:freechips.rocketchip.system.DefaultRV32Config.fir@24875.4]
  assign _GEN_31 = 4'h4 == _T_47 ? _T_246_4_last : _GEN_25; // @[Deinterleaver.scala 95:20:freechips.rocketchip.system.DefaultRV32Config.fir@24875.4]
  assign _GEN_37 = 4'h5 == _T_47 ? 1'h0 : _GEN_31; // @[Deinterleaver.scala 95:20:freechips.rocketchip.system.DefaultRV32Config.fir@24875.4]
  assign _GEN_43 = 4'h6 == _T_47 ? 1'h0 : _GEN_37; // @[Deinterleaver.scala 95:20:freechips.rocketchip.system.DefaultRV32Config.fir@24875.4]
  assign _GEN_49 = 4'h7 == _T_47 ? 1'h0 : _GEN_43; // @[Deinterleaver.scala 95:20:freechips.rocketchip.system.DefaultRV32Config.fir@24875.4]
  assign _GEN_55 = 4'h8 == _T_47 ? 1'h0 : _GEN_49; // @[Deinterleaver.scala 95:20:freechips.rocketchip.system.DefaultRV32Config.fir@24875.4]
  assign _GEN_61 = 4'h9 == _T_47 ? 1'h0 : _GEN_55; // @[Deinterleaver.scala 95:20:freechips.rocketchip.system.DefaultRV32Config.fir@24875.4]
  assign _GEN_67 = 4'ha == _T_47 ? 1'h0 : _GEN_61; // @[Deinterleaver.scala 95:20:freechips.rocketchip.system.DefaultRV32Config.fir@24875.4]
  assign _GEN_73 = 4'hb == _T_47 ? 1'h0 : _GEN_67; // @[Deinterleaver.scala 95:20:freechips.rocketchip.system.DefaultRV32Config.fir@24875.4]
  assign _GEN_79 = 4'hc == _T_47 ? 1'h0 : _GEN_73; // @[Deinterleaver.scala 95:20:freechips.rocketchip.system.DefaultRV32Config.fir@24875.4]
  assign _GEN_85 = 4'hd == _T_47 ? 1'h0 : _GEN_79; // @[Deinterleaver.scala 95:20:freechips.rocketchip.system.DefaultRV32Config.fir@24875.4]
  assign _GEN_91 = 4'he == _T_47 ? 1'h0 : _GEN_85; // @[Deinterleaver.scala 95:20:freechips.rocketchip.system.DefaultRV32Config.fir@24875.4]
  assign _GEN_97 = 4'hf == _T_47 ? 1'h0 : _GEN_91; // @[Deinterleaver.scala 95:20:freechips.rocketchip.system.DefaultRV32Config.fir@24875.4]
  assign _T_63 = _T_62 & _GEN_97; // @[Deinterleaver.scala 75:48:freechips.rocketchip.system.DefaultRV32Config.fir@24540.4]
  assign _GEN_114 = {{4'd0}, _T_59}; // @[Deinterleaver.scala 76:27:freechips.rocketchip.system.DefaultRV32Config.fir@24541.4]
  assign _T_65 = _T_54 + _GEN_114; // @[Deinterleaver.scala 76:27:freechips.rocketchip.system.DefaultRV32Config.fir@24542.4]
  assign _GEN_115 = {{4'd0}, _T_63}; // @[Deinterleaver.scala 76:40:freechips.rocketchip.system.DefaultRV32Config.fir@24543.4]
  assign _T_67 = _T_65 - _GEN_115; // @[Deinterleaver.scala 76:40:freechips.rocketchip.system.DefaultRV32Config.fir@24544.4]
  assign _T_68 = ~_T_63; // @[Deinterleaver.scala 79:21:freechips.rocketchip.system.DefaultRV32Config.fir@24547.4]
  assign _T_69 = _T_54 != 5'h0; // @[Deinterleaver.scala 79:35:freechips.rocketchip.system.DefaultRV32Config.fir@24548.4]
  assign _T_70 = _T_68 | _T_69; // @[Deinterleaver.scala 79:26:freechips.rocketchip.system.DefaultRV32Config.fir@24549.4]
  assign _T_72 = _T_70 | reset; // @[Deinterleaver.scala 79:20:freechips.rocketchip.system.DefaultRV32Config.fir@24551.4]
  assign _T_73 = ~_T_72; // @[Deinterleaver.scala 79:20:freechips.rocketchip.system.DefaultRV32Config.fir@24552.4]
  assign _T_74 = ~_T_59; // @[Deinterleaver.scala 80:21:freechips.rocketchip.system.DefaultRV32Config.fir@24557.4]
  assign _T_75 = _T_54 != 5'h10; // @[Deinterleaver.scala 80:35:freechips.rocketchip.system.DefaultRV32Config.fir@24558.4]
  assign _T_76 = _T_74 | _T_75; // @[Deinterleaver.scala 80:26:freechips.rocketchip.system.DefaultRV32Config.fir@24559.4]
  assign _T_78 = _T_76 | reset; // @[Deinterleaver.scala 80:20:freechips.rocketchip.system.DefaultRV32Config.fir@24561.4]
  assign _T_79 = ~_T_78; // @[Deinterleaver.scala 80:20:freechips.rocketchip.system.DefaultRV32Config.fir@24562.4]
  assign _T_80 = _T_67 != 5'h0; // @[Deinterleaver.scala 81:18:freechips.rocketchip.system.DefaultRV32Config.fir@24567.4]
  assign _T_85 = _T_52[1] & _T_57; // @[Deinterleaver.scala 74:33:freechips.rocketchip.system.DefaultRV32Config.fir@24572.4]
  assign _T_86 = _T_85 & auto_out_r_bits_last; // @[Deinterleaver.scala 74:49:freechips.rocketchip.system.DefaultRV32Config.fir@24573.4]
  assign _T_89 = _T_49[1] & _T_61; // @[Deinterleaver.scala 75:33:freechips.rocketchip.system.DefaultRV32Config.fir@24576.4]
  assign _T_90 = _T_89 & _GEN_97; // @[Deinterleaver.scala 75:48:freechips.rocketchip.system.DefaultRV32Config.fir@24577.4]
  assign _GEN_116 = {{4'd0}, _T_86}; // @[Deinterleaver.scala 76:27:freechips.rocketchip.system.DefaultRV32Config.fir@24578.4]
  assign _T_92 = _T_81 + _GEN_116; // @[Deinterleaver.scala 76:27:freechips.rocketchip.system.DefaultRV32Config.fir@24579.4]
  assign _GEN_117 = {{4'd0}, _T_90}; // @[Deinterleaver.scala 76:40:freechips.rocketchip.system.DefaultRV32Config.fir@24580.4]
  assign _T_94 = _T_92 - _GEN_117; // @[Deinterleaver.scala 76:40:freechips.rocketchip.system.DefaultRV32Config.fir@24581.4]
  assign _T_95 = ~_T_90; // @[Deinterleaver.scala 79:21:freechips.rocketchip.system.DefaultRV32Config.fir@24584.4]
  assign _T_96 = _T_81 != 5'h0; // @[Deinterleaver.scala 79:35:freechips.rocketchip.system.DefaultRV32Config.fir@24585.4]
  assign _T_97 = _T_95 | _T_96; // @[Deinterleaver.scala 79:26:freechips.rocketchip.system.DefaultRV32Config.fir@24586.4]
  assign _T_99 = _T_97 | reset; // @[Deinterleaver.scala 79:20:freechips.rocketchip.system.DefaultRV32Config.fir@24588.4]
  assign _T_100 = ~_T_99; // @[Deinterleaver.scala 79:20:freechips.rocketchip.system.DefaultRV32Config.fir@24589.4]
  assign _T_101 = ~_T_86; // @[Deinterleaver.scala 80:21:freechips.rocketchip.system.DefaultRV32Config.fir@24594.4]
  assign _T_102 = _T_81 != 5'h10; // @[Deinterleaver.scala 80:35:freechips.rocketchip.system.DefaultRV32Config.fir@24595.4]
  assign _T_103 = _T_101 | _T_102; // @[Deinterleaver.scala 80:26:freechips.rocketchip.system.DefaultRV32Config.fir@24596.4]
  assign _T_105 = _T_103 | reset; // @[Deinterleaver.scala 80:20:freechips.rocketchip.system.DefaultRV32Config.fir@24598.4]
  assign _T_106 = ~_T_105; // @[Deinterleaver.scala 80:20:freechips.rocketchip.system.DefaultRV32Config.fir@24599.4]
  assign _T_107 = _T_94 != 5'h0; // @[Deinterleaver.scala 81:18:freechips.rocketchip.system.DefaultRV32Config.fir@24604.4]
  assign _T_112 = _T_52[2] & _T_57; // @[Deinterleaver.scala 74:33:freechips.rocketchip.system.DefaultRV32Config.fir@24609.4]
  assign _T_113 = _T_112 & auto_out_r_bits_last; // @[Deinterleaver.scala 74:49:freechips.rocketchip.system.DefaultRV32Config.fir@24610.4]
  assign _T_116 = _T_49[2] & _T_61; // @[Deinterleaver.scala 75:33:freechips.rocketchip.system.DefaultRV32Config.fir@24613.4]
  assign _T_117 = _T_116 & _GEN_97; // @[Deinterleaver.scala 75:48:freechips.rocketchip.system.DefaultRV32Config.fir@24614.4]
  assign _GEN_118 = {{4'd0}, _T_113}; // @[Deinterleaver.scala 76:27:freechips.rocketchip.system.DefaultRV32Config.fir@24615.4]
  assign _T_119 = _T_108 + _GEN_118; // @[Deinterleaver.scala 76:27:freechips.rocketchip.system.DefaultRV32Config.fir@24616.4]
  assign _GEN_119 = {{4'd0}, _T_117}; // @[Deinterleaver.scala 76:40:freechips.rocketchip.system.DefaultRV32Config.fir@24617.4]
  assign _T_121 = _T_119 - _GEN_119; // @[Deinterleaver.scala 76:40:freechips.rocketchip.system.DefaultRV32Config.fir@24618.4]
  assign _T_122 = ~_T_117; // @[Deinterleaver.scala 79:21:freechips.rocketchip.system.DefaultRV32Config.fir@24621.4]
  assign _T_123 = _T_108 != 5'h0; // @[Deinterleaver.scala 79:35:freechips.rocketchip.system.DefaultRV32Config.fir@24622.4]
  assign _T_124 = _T_122 | _T_123; // @[Deinterleaver.scala 79:26:freechips.rocketchip.system.DefaultRV32Config.fir@24623.4]
  assign _T_126 = _T_124 | reset; // @[Deinterleaver.scala 79:20:freechips.rocketchip.system.DefaultRV32Config.fir@24625.4]
  assign _T_127 = ~_T_126; // @[Deinterleaver.scala 79:20:freechips.rocketchip.system.DefaultRV32Config.fir@24626.4]
  assign _T_128 = ~_T_113; // @[Deinterleaver.scala 80:21:freechips.rocketchip.system.DefaultRV32Config.fir@24631.4]
  assign _T_129 = _T_108 != 5'h10; // @[Deinterleaver.scala 80:35:freechips.rocketchip.system.DefaultRV32Config.fir@24632.4]
  assign _T_130 = _T_128 | _T_129; // @[Deinterleaver.scala 80:26:freechips.rocketchip.system.DefaultRV32Config.fir@24633.4]
  assign _T_132 = _T_130 | reset; // @[Deinterleaver.scala 80:20:freechips.rocketchip.system.DefaultRV32Config.fir@24635.4]
  assign _T_133 = ~_T_132; // @[Deinterleaver.scala 80:20:freechips.rocketchip.system.DefaultRV32Config.fir@24636.4]
  assign _T_134 = _T_121 != 5'h0; // @[Deinterleaver.scala 81:18:freechips.rocketchip.system.DefaultRV32Config.fir@24641.4]
  assign _T_139 = _T_52[3] & _T_57; // @[Deinterleaver.scala 74:33:freechips.rocketchip.system.DefaultRV32Config.fir@24646.4]
  assign _T_140 = _T_139 & auto_out_r_bits_last; // @[Deinterleaver.scala 74:49:freechips.rocketchip.system.DefaultRV32Config.fir@24647.4]
  assign _T_143 = _T_49[3] & _T_61; // @[Deinterleaver.scala 75:33:freechips.rocketchip.system.DefaultRV32Config.fir@24650.4]
  assign _T_144 = _T_143 & _GEN_97; // @[Deinterleaver.scala 75:48:freechips.rocketchip.system.DefaultRV32Config.fir@24651.4]
  assign _GEN_120 = {{4'd0}, _T_140}; // @[Deinterleaver.scala 76:27:freechips.rocketchip.system.DefaultRV32Config.fir@24652.4]
  assign _T_146 = _T_135 + _GEN_120; // @[Deinterleaver.scala 76:27:freechips.rocketchip.system.DefaultRV32Config.fir@24653.4]
  assign _GEN_121 = {{4'd0}, _T_144}; // @[Deinterleaver.scala 76:40:freechips.rocketchip.system.DefaultRV32Config.fir@24654.4]
  assign _T_148 = _T_146 - _GEN_121; // @[Deinterleaver.scala 76:40:freechips.rocketchip.system.DefaultRV32Config.fir@24655.4]
  assign _T_149 = ~_T_144; // @[Deinterleaver.scala 79:21:freechips.rocketchip.system.DefaultRV32Config.fir@24658.4]
  assign _T_150 = _T_135 != 5'h0; // @[Deinterleaver.scala 79:35:freechips.rocketchip.system.DefaultRV32Config.fir@24659.4]
  assign _T_151 = _T_149 | _T_150; // @[Deinterleaver.scala 79:26:freechips.rocketchip.system.DefaultRV32Config.fir@24660.4]
  assign _T_153 = _T_151 | reset; // @[Deinterleaver.scala 79:20:freechips.rocketchip.system.DefaultRV32Config.fir@24662.4]
  assign _T_154 = ~_T_153; // @[Deinterleaver.scala 79:20:freechips.rocketchip.system.DefaultRV32Config.fir@24663.4]
  assign _T_155 = ~_T_140; // @[Deinterleaver.scala 80:21:freechips.rocketchip.system.DefaultRV32Config.fir@24668.4]
  assign _T_156 = _T_135 != 5'h10; // @[Deinterleaver.scala 80:35:freechips.rocketchip.system.DefaultRV32Config.fir@24669.4]
  assign _T_157 = _T_155 | _T_156; // @[Deinterleaver.scala 80:26:freechips.rocketchip.system.DefaultRV32Config.fir@24670.4]
  assign _T_159 = _T_157 | reset; // @[Deinterleaver.scala 80:20:freechips.rocketchip.system.DefaultRV32Config.fir@24672.4]
  assign _T_160 = ~_T_159; // @[Deinterleaver.scala 80:20:freechips.rocketchip.system.DefaultRV32Config.fir@24673.4]
  assign _T_161 = _T_148 != 5'h0; // @[Deinterleaver.scala 81:18:freechips.rocketchip.system.DefaultRV32Config.fir@24678.4]
  assign _T_166 = _T_52[4] & _T_57; // @[Deinterleaver.scala 74:33:freechips.rocketchip.system.DefaultRV32Config.fir@24683.4]
  assign _T_167 = _T_166 & auto_out_r_bits_last; // @[Deinterleaver.scala 74:49:freechips.rocketchip.system.DefaultRV32Config.fir@24684.4]
  assign _T_170 = _T_49[4] & _T_61; // @[Deinterleaver.scala 75:33:freechips.rocketchip.system.DefaultRV32Config.fir@24687.4]
  assign _T_171 = _T_170 & _GEN_97; // @[Deinterleaver.scala 75:48:freechips.rocketchip.system.DefaultRV32Config.fir@24688.4]
  assign _GEN_122 = {{4'd0}, _T_167}; // @[Deinterleaver.scala 76:27:freechips.rocketchip.system.DefaultRV32Config.fir@24689.4]
  assign _T_173 = _T_162 + _GEN_122; // @[Deinterleaver.scala 76:27:freechips.rocketchip.system.DefaultRV32Config.fir@24690.4]
  assign _GEN_123 = {{4'd0}, _T_171}; // @[Deinterleaver.scala 76:40:freechips.rocketchip.system.DefaultRV32Config.fir@24691.4]
  assign _T_175 = _T_173 - _GEN_123; // @[Deinterleaver.scala 76:40:freechips.rocketchip.system.DefaultRV32Config.fir@24692.4]
  assign _T_176 = ~_T_171; // @[Deinterleaver.scala 79:21:freechips.rocketchip.system.DefaultRV32Config.fir@24695.4]
  assign _T_177 = _T_162 != 5'h0; // @[Deinterleaver.scala 79:35:freechips.rocketchip.system.DefaultRV32Config.fir@24696.4]
  assign _T_178 = _T_176 | _T_177; // @[Deinterleaver.scala 79:26:freechips.rocketchip.system.DefaultRV32Config.fir@24697.4]
  assign _T_180 = _T_178 | reset; // @[Deinterleaver.scala 79:20:freechips.rocketchip.system.DefaultRV32Config.fir@24699.4]
  assign _T_181 = ~_T_180; // @[Deinterleaver.scala 79:20:freechips.rocketchip.system.DefaultRV32Config.fir@24700.4]
  assign _T_182 = ~_T_167; // @[Deinterleaver.scala 80:21:freechips.rocketchip.system.DefaultRV32Config.fir@24705.4]
  assign _T_183 = _T_162 != 5'h10; // @[Deinterleaver.scala 80:35:freechips.rocketchip.system.DefaultRV32Config.fir@24706.4]
  assign _T_184 = _T_182 | _T_183; // @[Deinterleaver.scala 80:26:freechips.rocketchip.system.DefaultRV32Config.fir@24707.4]
  assign _T_186 = _T_184 | reset; // @[Deinterleaver.scala 80:20:freechips.rocketchip.system.DefaultRV32Config.fir@24709.4]
  assign _T_187 = ~_T_186; // @[Deinterleaver.scala 80:20:freechips.rocketchip.system.DefaultRV32Config.fir@24710.4]
  assign _T_188 = _T_175 != 5'h0; // @[Deinterleaver.scala 81:18:freechips.rocketchip.system.DefaultRV32Config.fir@24715.4]
  assign _T_203 = {8'h0,2'h0,1'h0,_T_188,_T_161,_T_134,_T_107,_T_80}; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@24730.4]
  assign _T_204 = {_T_203, 1'h0}; // @[package.scala 217:48:freechips.rocketchip.system.DefaultRV32Config.fir@24731.4]
  assign _T_206 = _T_203 | _T_204[15:0]; // @[package.scala 217:43:freechips.rocketchip.system.DefaultRV32Config.fir@24733.4]
  assign _T_207 = {_T_206, 2'h0}; // @[package.scala 217:48:freechips.rocketchip.system.DefaultRV32Config.fir@24734.4]
  assign _T_209 = _T_206 | _T_207[15:0]; // @[package.scala 217:43:freechips.rocketchip.system.DefaultRV32Config.fir@24736.4]
  assign _T_210 = {_T_209, 4'h0}; // @[package.scala 217:48:freechips.rocketchip.system.DefaultRV32Config.fir@24737.4]
  assign _T_212 = _T_209 | _T_210[15:0]; // @[package.scala 217:43:freechips.rocketchip.system.DefaultRV32Config.fir@24739.4]
  assign _T_213 = {_T_212, 8'h0}; // @[package.scala 217:48:freechips.rocketchip.system.DefaultRV32Config.fir@24740.4]
  assign _T_215 = _T_212 | _T_213[15:0]; // @[package.scala 217:43:freechips.rocketchip.system.DefaultRV32Config.fir@24742.4]
  assign _T_217 = {_T_215, 1'h0}; // @[Deinterleaver.scala 86:51:freechips.rocketchip.system.DefaultRV32Config.fir@24744.4]
  assign _T_218 = ~_T_217; // @[Deinterleaver.scala 86:33:freechips.rocketchip.system.DefaultRV32Config.fir@24745.4]
  assign _GEN_124 = {{1'd0}, _T_203}; // @[Deinterleaver.scala 86:31:freechips.rocketchip.system.DefaultRV32Config.fir@24746.4]
  assign _T_219 = _GEN_124 & _T_218; // @[Deinterleaver.scala 86:31:freechips.rocketchip.system.DefaultRV32Config.fir@24746.4]
  assign _T_220 = ~_T_46; // @[Deinterleaver.scala 87:15:freechips.rocketchip.system.DefaultRV32Config.fir@24747.4]
  assign _T_222 = _T_61 & _GEN_97; // @[Deinterleaver.scala 87:39:freechips.rocketchip.system.DefaultRV32Config.fir@24749.4]
  assign _T_223 = _T_220 | _T_222; // @[Deinterleaver.scala 87:23:freechips.rocketchip.system.DefaultRV32Config.fir@24750.4]
  assign _T_224 = |_T_203; // @[Deinterleaver.scala 88:29:freechips.rocketchip.system.DefaultRV32Config.fir@24752.6]
  assign _T_227 = |_T_219[16]; // @[OneHot.scala 32:14:freechips.rocketchip.system.DefaultRV32Config.fir@24756.6]
  assign _GEN_125 = {{15'd0}, _T_219[16]}; // @[OneHot.scala 32:28:freechips.rocketchip.system.DefaultRV32Config.fir@24757.6]
  assign _T_228 = _GEN_125 | _T_219[15:0]; // @[OneHot.scala 32:28:freechips.rocketchip.system.DefaultRV32Config.fir@24757.6]
  assign _T_231 = |_T_228[15:8]; // @[OneHot.scala 32:14:freechips.rocketchip.system.DefaultRV32Config.fir@24760.6]
  assign _T_232 = _T_228[15:8] | _T_228[7:0]; // @[OneHot.scala 32:28:freechips.rocketchip.system.DefaultRV32Config.fir@24761.6]
  assign _T_235 = |_T_232[7:4]; // @[OneHot.scala 32:14:freechips.rocketchip.system.DefaultRV32Config.fir@24764.6]
  assign _T_236 = _T_232[7:4] | _T_232[3:0]; // @[OneHot.scala 32:28:freechips.rocketchip.system.DefaultRV32Config.fir@24765.6]
  assign _T_239 = |_T_236[3:2]; // @[OneHot.scala 32:14:freechips.rocketchip.system.DefaultRV32Config.fir@24768.6]
  assign _T_240 = _T_236[3:2] | _T_236[1:0]; // @[OneHot.scala 32:28:freechips.rocketchip.system.DefaultRV32Config.fir@24769.6]
  assign _T_245 = {_T_227,_T_231,_T_235,_T_239,_T_240[1]}; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@24774.6]
  assign _GEN_1 = _T_223 ? _T_245 : {{1'd0}, _T_47}; // @[Deinterleaver.scala 87:59:freechips.rocketchip.system.DefaultRV32Config.fir@24751.4]
  assign _T_246_0_id = queue_0_io_deq_bits_id; // @[Deinterleaver.scala 94:31:freechips.rocketchip.system.DefaultRV32Config.fir@24778.4 Deinterleaver.scala 94:31:freechips.rocketchip.system.DefaultRV32Config.fir@24784.4]
  assign _T_246_0_data = queue_0_io_deq_bits_data; // @[Deinterleaver.scala 94:31:freechips.rocketchip.system.DefaultRV32Config.fir@24778.4 Deinterleaver.scala 94:31:freechips.rocketchip.system.DefaultRV32Config.fir@24783.4]
  assign _T_246_0_resp = queue_0_io_deq_bits_resp; // @[Deinterleaver.scala 94:31:freechips.rocketchip.system.DefaultRV32Config.fir@24778.4 Deinterleaver.scala 94:31:freechips.rocketchip.system.DefaultRV32Config.fir@24782.4]
  assign _T_246_0_echo_tl_state_size = queue_0_io_deq_bits_echo_tl_state_size; // @[Deinterleaver.scala 94:31:freechips.rocketchip.system.DefaultRV32Config.fir@24778.4 Deinterleaver.scala 94:31:freechips.rocketchip.system.DefaultRV32Config.fir@24781.4]
  assign _T_246_0_echo_tl_state_source = queue_0_io_deq_bits_echo_tl_state_source; // @[Deinterleaver.scala 94:31:freechips.rocketchip.system.DefaultRV32Config.fir@24778.4 Deinterleaver.scala 94:31:freechips.rocketchip.system.DefaultRV32Config.fir@24780.4]
  assign _T_246_1_id = queue_1_io_deq_bits_id; // @[Deinterleaver.scala 94:31:freechips.rocketchip.system.DefaultRV32Config.fir@24778.4 Deinterleaver.scala 94:31:freechips.rocketchip.system.DefaultRV32Config.fir@24790.4]
  assign _GEN_8 = 4'h1 == _T_47 ? _T_246_1_id : _T_246_0_id; // @[Deinterleaver.scala 95:20:freechips.rocketchip.system.DefaultRV32Config.fir@24875.4]
  assign _T_246_1_data = queue_1_io_deq_bits_data; // @[Deinterleaver.scala 94:31:freechips.rocketchip.system.DefaultRV32Config.fir@24778.4 Deinterleaver.scala 94:31:freechips.rocketchip.system.DefaultRV32Config.fir@24789.4]
  assign _GEN_9 = 4'h1 == _T_47 ? _T_246_1_data : _T_246_0_data; // @[Deinterleaver.scala 95:20:freechips.rocketchip.system.DefaultRV32Config.fir@24875.4]
  assign _T_246_1_resp = queue_1_io_deq_bits_resp; // @[Deinterleaver.scala 94:31:freechips.rocketchip.system.DefaultRV32Config.fir@24778.4 Deinterleaver.scala 94:31:freechips.rocketchip.system.DefaultRV32Config.fir@24788.4]
  assign _GEN_10 = 4'h1 == _T_47 ? _T_246_1_resp : _T_246_0_resp; // @[Deinterleaver.scala 95:20:freechips.rocketchip.system.DefaultRV32Config.fir@24875.4]
  assign _T_246_1_echo_tl_state_size = queue_1_io_deq_bits_echo_tl_state_size; // @[Deinterleaver.scala 94:31:freechips.rocketchip.system.DefaultRV32Config.fir@24778.4 Deinterleaver.scala 94:31:freechips.rocketchip.system.DefaultRV32Config.fir@24787.4]
  assign _GEN_11 = 4'h1 == _T_47 ? _T_246_1_echo_tl_state_size : _T_246_0_echo_tl_state_size; // @[Deinterleaver.scala 95:20:freechips.rocketchip.system.DefaultRV32Config.fir@24875.4]
  assign _T_246_1_echo_tl_state_source = queue_1_io_deq_bits_echo_tl_state_source; // @[Deinterleaver.scala 94:31:freechips.rocketchip.system.DefaultRV32Config.fir@24778.4 Deinterleaver.scala 94:31:freechips.rocketchip.system.DefaultRV32Config.fir@24786.4]
  assign _GEN_12 = 4'h1 == _T_47 ? _T_246_1_echo_tl_state_source : _T_246_0_echo_tl_state_source; // @[Deinterleaver.scala 95:20:freechips.rocketchip.system.DefaultRV32Config.fir@24875.4]
  assign _T_246_2_id = queue_2_io_deq_bits_id; // @[Deinterleaver.scala 94:31:freechips.rocketchip.system.DefaultRV32Config.fir@24778.4 Deinterleaver.scala 94:31:freechips.rocketchip.system.DefaultRV32Config.fir@24796.4]
  assign _GEN_14 = 4'h2 == _T_47 ? _T_246_2_id : _GEN_8; // @[Deinterleaver.scala 95:20:freechips.rocketchip.system.DefaultRV32Config.fir@24875.4]
  assign _T_246_2_data = queue_2_io_deq_bits_data; // @[Deinterleaver.scala 94:31:freechips.rocketchip.system.DefaultRV32Config.fir@24778.4 Deinterleaver.scala 94:31:freechips.rocketchip.system.DefaultRV32Config.fir@24795.4]
  assign _GEN_15 = 4'h2 == _T_47 ? _T_246_2_data : _GEN_9; // @[Deinterleaver.scala 95:20:freechips.rocketchip.system.DefaultRV32Config.fir@24875.4]
  assign _T_246_2_resp = queue_2_io_deq_bits_resp; // @[Deinterleaver.scala 94:31:freechips.rocketchip.system.DefaultRV32Config.fir@24778.4 Deinterleaver.scala 94:31:freechips.rocketchip.system.DefaultRV32Config.fir@24794.4]
  assign _GEN_16 = 4'h2 == _T_47 ? _T_246_2_resp : _GEN_10; // @[Deinterleaver.scala 95:20:freechips.rocketchip.system.DefaultRV32Config.fir@24875.4]
  assign _T_246_2_echo_tl_state_size = queue_2_io_deq_bits_echo_tl_state_size; // @[Deinterleaver.scala 94:31:freechips.rocketchip.system.DefaultRV32Config.fir@24778.4 Deinterleaver.scala 94:31:freechips.rocketchip.system.DefaultRV32Config.fir@24793.4]
  assign _GEN_17 = 4'h2 == _T_47 ? _T_246_2_echo_tl_state_size : _GEN_11; // @[Deinterleaver.scala 95:20:freechips.rocketchip.system.DefaultRV32Config.fir@24875.4]
  assign _T_246_2_echo_tl_state_source = queue_2_io_deq_bits_echo_tl_state_source; // @[Deinterleaver.scala 94:31:freechips.rocketchip.system.DefaultRV32Config.fir@24778.4 Deinterleaver.scala 94:31:freechips.rocketchip.system.DefaultRV32Config.fir@24792.4]
  assign _GEN_18 = 4'h2 == _T_47 ? _T_246_2_echo_tl_state_source : _GEN_12; // @[Deinterleaver.scala 95:20:freechips.rocketchip.system.DefaultRV32Config.fir@24875.4]
  assign _T_246_3_id = queue_3_io_deq_bits_id; // @[Deinterleaver.scala 94:31:freechips.rocketchip.system.DefaultRV32Config.fir@24778.4 Deinterleaver.scala 94:31:freechips.rocketchip.system.DefaultRV32Config.fir@24802.4]
  assign _GEN_20 = 4'h3 == _T_47 ? _T_246_3_id : _GEN_14; // @[Deinterleaver.scala 95:20:freechips.rocketchip.system.DefaultRV32Config.fir@24875.4]
  assign _T_246_3_data = queue_3_io_deq_bits_data; // @[Deinterleaver.scala 94:31:freechips.rocketchip.system.DefaultRV32Config.fir@24778.4 Deinterleaver.scala 94:31:freechips.rocketchip.system.DefaultRV32Config.fir@24801.4]
  assign _GEN_21 = 4'h3 == _T_47 ? _T_246_3_data : _GEN_15; // @[Deinterleaver.scala 95:20:freechips.rocketchip.system.DefaultRV32Config.fir@24875.4]
  assign _T_246_3_resp = queue_3_io_deq_bits_resp; // @[Deinterleaver.scala 94:31:freechips.rocketchip.system.DefaultRV32Config.fir@24778.4 Deinterleaver.scala 94:31:freechips.rocketchip.system.DefaultRV32Config.fir@24800.4]
  assign _GEN_22 = 4'h3 == _T_47 ? _T_246_3_resp : _GEN_16; // @[Deinterleaver.scala 95:20:freechips.rocketchip.system.DefaultRV32Config.fir@24875.4]
  assign _T_246_3_echo_tl_state_size = queue_3_io_deq_bits_echo_tl_state_size; // @[Deinterleaver.scala 94:31:freechips.rocketchip.system.DefaultRV32Config.fir@24778.4 Deinterleaver.scala 94:31:freechips.rocketchip.system.DefaultRV32Config.fir@24799.4]
  assign _GEN_23 = 4'h3 == _T_47 ? _T_246_3_echo_tl_state_size : _GEN_17; // @[Deinterleaver.scala 95:20:freechips.rocketchip.system.DefaultRV32Config.fir@24875.4]
  assign _T_246_3_echo_tl_state_source = queue_3_io_deq_bits_echo_tl_state_source; // @[Deinterleaver.scala 94:31:freechips.rocketchip.system.DefaultRV32Config.fir@24778.4 Deinterleaver.scala 94:31:freechips.rocketchip.system.DefaultRV32Config.fir@24798.4]
  assign _GEN_24 = 4'h3 == _T_47 ? _T_246_3_echo_tl_state_source : _GEN_18; // @[Deinterleaver.scala 95:20:freechips.rocketchip.system.DefaultRV32Config.fir@24875.4]
  assign _T_246_4_id = queue_4_io_deq_bits_id; // @[Deinterleaver.scala 94:31:freechips.rocketchip.system.DefaultRV32Config.fir@24778.4 Deinterleaver.scala 94:31:freechips.rocketchip.system.DefaultRV32Config.fir@24808.4]
  assign _GEN_26 = 4'h4 == _T_47 ? _T_246_4_id : _GEN_20; // @[Deinterleaver.scala 95:20:freechips.rocketchip.system.DefaultRV32Config.fir@24875.4]
  assign _T_246_4_data = queue_4_io_deq_bits_data; // @[Deinterleaver.scala 94:31:freechips.rocketchip.system.DefaultRV32Config.fir@24778.4 Deinterleaver.scala 94:31:freechips.rocketchip.system.DefaultRV32Config.fir@24807.4]
  assign _GEN_27 = 4'h4 == _T_47 ? _T_246_4_data : _GEN_21; // @[Deinterleaver.scala 95:20:freechips.rocketchip.system.DefaultRV32Config.fir@24875.4]
  assign _T_246_4_resp = queue_4_io_deq_bits_resp; // @[Deinterleaver.scala 94:31:freechips.rocketchip.system.DefaultRV32Config.fir@24778.4 Deinterleaver.scala 94:31:freechips.rocketchip.system.DefaultRV32Config.fir@24806.4]
  assign _GEN_28 = 4'h4 == _T_47 ? _T_246_4_resp : _GEN_22; // @[Deinterleaver.scala 95:20:freechips.rocketchip.system.DefaultRV32Config.fir@24875.4]
  assign _T_246_4_echo_tl_state_size = queue_4_io_deq_bits_echo_tl_state_size; // @[Deinterleaver.scala 94:31:freechips.rocketchip.system.DefaultRV32Config.fir@24778.4 Deinterleaver.scala 94:31:freechips.rocketchip.system.DefaultRV32Config.fir@24805.4]
  assign _GEN_29 = 4'h4 == _T_47 ? _T_246_4_echo_tl_state_size : _GEN_23; // @[Deinterleaver.scala 95:20:freechips.rocketchip.system.DefaultRV32Config.fir@24875.4]
  assign _T_246_4_echo_tl_state_source = queue_4_io_deq_bits_echo_tl_state_source; // @[Deinterleaver.scala 94:31:freechips.rocketchip.system.DefaultRV32Config.fir@24778.4 Deinterleaver.scala 94:31:freechips.rocketchip.system.DefaultRV32Config.fir@24804.4]
  assign _GEN_30 = 4'h4 == _T_47 ? _T_246_4_echo_tl_state_source : _GEN_24; // @[Deinterleaver.scala 95:20:freechips.rocketchip.system.DefaultRV32Config.fir@24875.4]
  assign _GEN_32 = 4'h5 == _T_47 ? 4'h0 : _GEN_26; // @[Deinterleaver.scala 95:20:freechips.rocketchip.system.DefaultRV32Config.fir@24875.4]
  assign _GEN_33 = 4'h5 == _T_47 ? 32'h0 : _GEN_27; // @[Deinterleaver.scala 95:20:freechips.rocketchip.system.DefaultRV32Config.fir@24875.4]
  assign _GEN_34 = 4'h5 == _T_47 ? 2'h0 : _GEN_28; // @[Deinterleaver.scala 95:20:freechips.rocketchip.system.DefaultRV32Config.fir@24875.4]
  assign _GEN_35 = 4'h5 == _T_47 ? 4'h0 : _GEN_29; // @[Deinterleaver.scala 95:20:freechips.rocketchip.system.DefaultRV32Config.fir@24875.4]
  assign _GEN_36 = 4'h5 == _T_47 ? 5'h0 : _GEN_30; // @[Deinterleaver.scala 95:20:freechips.rocketchip.system.DefaultRV32Config.fir@24875.4]
  assign _GEN_38 = 4'h6 == _T_47 ? 4'h0 : _GEN_32; // @[Deinterleaver.scala 95:20:freechips.rocketchip.system.DefaultRV32Config.fir@24875.4]
  assign _GEN_39 = 4'h6 == _T_47 ? 32'h0 : _GEN_33; // @[Deinterleaver.scala 95:20:freechips.rocketchip.system.DefaultRV32Config.fir@24875.4]
  assign _GEN_40 = 4'h6 == _T_47 ? 2'h0 : _GEN_34; // @[Deinterleaver.scala 95:20:freechips.rocketchip.system.DefaultRV32Config.fir@24875.4]
  assign _GEN_41 = 4'h6 == _T_47 ? 4'h0 : _GEN_35; // @[Deinterleaver.scala 95:20:freechips.rocketchip.system.DefaultRV32Config.fir@24875.4]
  assign _GEN_42 = 4'h6 == _T_47 ? 5'h0 : _GEN_36; // @[Deinterleaver.scala 95:20:freechips.rocketchip.system.DefaultRV32Config.fir@24875.4]
  assign _GEN_44 = 4'h7 == _T_47 ? 4'h0 : _GEN_38; // @[Deinterleaver.scala 95:20:freechips.rocketchip.system.DefaultRV32Config.fir@24875.4]
  assign _GEN_45 = 4'h7 == _T_47 ? 32'h0 : _GEN_39; // @[Deinterleaver.scala 95:20:freechips.rocketchip.system.DefaultRV32Config.fir@24875.4]
  assign _GEN_46 = 4'h7 == _T_47 ? 2'h0 : _GEN_40; // @[Deinterleaver.scala 95:20:freechips.rocketchip.system.DefaultRV32Config.fir@24875.4]
  assign _GEN_47 = 4'h7 == _T_47 ? 4'h0 : _GEN_41; // @[Deinterleaver.scala 95:20:freechips.rocketchip.system.DefaultRV32Config.fir@24875.4]
  assign _GEN_48 = 4'h7 == _T_47 ? 5'h0 : _GEN_42; // @[Deinterleaver.scala 95:20:freechips.rocketchip.system.DefaultRV32Config.fir@24875.4]
  assign _GEN_50 = 4'h8 == _T_47 ? 4'h0 : _GEN_44; // @[Deinterleaver.scala 95:20:freechips.rocketchip.system.DefaultRV32Config.fir@24875.4]
  assign _GEN_51 = 4'h8 == _T_47 ? 32'h0 : _GEN_45; // @[Deinterleaver.scala 95:20:freechips.rocketchip.system.DefaultRV32Config.fir@24875.4]
  assign _GEN_52 = 4'h8 == _T_47 ? 2'h0 : _GEN_46; // @[Deinterleaver.scala 95:20:freechips.rocketchip.system.DefaultRV32Config.fir@24875.4]
  assign _GEN_53 = 4'h8 == _T_47 ? 4'h0 : _GEN_47; // @[Deinterleaver.scala 95:20:freechips.rocketchip.system.DefaultRV32Config.fir@24875.4]
  assign _GEN_54 = 4'h8 == _T_47 ? 5'h0 : _GEN_48; // @[Deinterleaver.scala 95:20:freechips.rocketchip.system.DefaultRV32Config.fir@24875.4]
  assign _GEN_56 = 4'h9 == _T_47 ? 4'h0 : _GEN_50; // @[Deinterleaver.scala 95:20:freechips.rocketchip.system.DefaultRV32Config.fir@24875.4]
  assign _GEN_57 = 4'h9 == _T_47 ? 32'h0 : _GEN_51; // @[Deinterleaver.scala 95:20:freechips.rocketchip.system.DefaultRV32Config.fir@24875.4]
  assign _GEN_58 = 4'h9 == _T_47 ? 2'h0 : _GEN_52; // @[Deinterleaver.scala 95:20:freechips.rocketchip.system.DefaultRV32Config.fir@24875.4]
  assign _GEN_59 = 4'h9 == _T_47 ? 4'h0 : _GEN_53; // @[Deinterleaver.scala 95:20:freechips.rocketchip.system.DefaultRV32Config.fir@24875.4]
  assign _GEN_60 = 4'h9 == _T_47 ? 5'h0 : _GEN_54; // @[Deinterleaver.scala 95:20:freechips.rocketchip.system.DefaultRV32Config.fir@24875.4]
  assign _GEN_62 = 4'ha == _T_47 ? 4'h0 : _GEN_56; // @[Deinterleaver.scala 95:20:freechips.rocketchip.system.DefaultRV32Config.fir@24875.4]
  assign _GEN_63 = 4'ha == _T_47 ? 32'h0 : _GEN_57; // @[Deinterleaver.scala 95:20:freechips.rocketchip.system.DefaultRV32Config.fir@24875.4]
  assign _GEN_64 = 4'ha == _T_47 ? 2'h0 : _GEN_58; // @[Deinterleaver.scala 95:20:freechips.rocketchip.system.DefaultRV32Config.fir@24875.4]
  assign _GEN_65 = 4'ha == _T_47 ? 4'h0 : _GEN_59; // @[Deinterleaver.scala 95:20:freechips.rocketchip.system.DefaultRV32Config.fir@24875.4]
  assign _GEN_66 = 4'ha == _T_47 ? 5'h0 : _GEN_60; // @[Deinterleaver.scala 95:20:freechips.rocketchip.system.DefaultRV32Config.fir@24875.4]
  assign _GEN_68 = 4'hb == _T_47 ? 4'h0 : _GEN_62; // @[Deinterleaver.scala 95:20:freechips.rocketchip.system.DefaultRV32Config.fir@24875.4]
  assign _GEN_69 = 4'hb == _T_47 ? 32'h0 : _GEN_63; // @[Deinterleaver.scala 95:20:freechips.rocketchip.system.DefaultRV32Config.fir@24875.4]
  assign _GEN_70 = 4'hb == _T_47 ? 2'h0 : _GEN_64; // @[Deinterleaver.scala 95:20:freechips.rocketchip.system.DefaultRV32Config.fir@24875.4]
  assign _GEN_71 = 4'hb == _T_47 ? 4'h0 : _GEN_65; // @[Deinterleaver.scala 95:20:freechips.rocketchip.system.DefaultRV32Config.fir@24875.4]
  assign _GEN_72 = 4'hb == _T_47 ? 5'h0 : _GEN_66; // @[Deinterleaver.scala 95:20:freechips.rocketchip.system.DefaultRV32Config.fir@24875.4]
  assign _GEN_74 = 4'hc == _T_47 ? 4'h0 : _GEN_68; // @[Deinterleaver.scala 95:20:freechips.rocketchip.system.DefaultRV32Config.fir@24875.4]
  assign _GEN_75 = 4'hc == _T_47 ? 32'h0 : _GEN_69; // @[Deinterleaver.scala 95:20:freechips.rocketchip.system.DefaultRV32Config.fir@24875.4]
  assign _GEN_76 = 4'hc == _T_47 ? 2'h0 : _GEN_70; // @[Deinterleaver.scala 95:20:freechips.rocketchip.system.DefaultRV32Config.fir@24875.4]
  assign _GEN_77 = 4'hc == _T_47 ? 4'h0 : _GEN_71; // @[Deinterleaver.scala 95:20:freechips.rocketchip.system.DefaultRV32Config.fir@24875.4]
  assign _GEN_78 = 4'hc == _T_47 ? 5'h0 : _GEN_72; // @[Deinterleaver.scala 95:20:freechips.rocketchip.system.DefaultRV32Config.fir@24875.4]
  assign _GEN_80 = 4'hd == _T_47 ? 4'h0 : _GEN_74; // @[Deinterleaver.scala 95:20:freechips.rocketchip.system.DefaultRV32Config.fir@24875.4]
  assign _GEN_81 = 4'hd == _T_47 ? 32'h0 : _GEN_75; // @[Deinterleaver.scala 95:20:freechips.rocketchip.system.DefaultRV32Config.fir@24875.4]
  assign _GEN_82 = 4'hd == _T_47 ? 2'h0 : _GEN_76; // @[Deinterleaver.scala 95:20:freechips.rocketchip.system.DefaultRV32Config.fir@24875.4]
  assign _GEN_83 = 4'hd == _T_47 ? 4'h0 : _GEN_77; // @[Deinterleaver.scala 95:20:freechips.rocketchip.system.DefaultRV32Config.fir@24875.4]
  assign _GEN_84 = 4'hd == _T_47 ? 5'h0 : _GEN_78; // @[Deinterleaver.scala 95:20:freechips.rocketchip.system.DefaultRV32Config.fir@24875.4]
  assign _GEN_86 = 4'he == _T_47 ? 4'h0 : _GEN_80; // @[Deinterleaver.scala 95:20:freechips.rocketchip.system.DefaultRV32Config.fir@24875.4]
  assign _GEN_87 = 4'he == _T_47 ? 32'h0 : _GEN_81; // @[Deinterleaver.scala 95:20:freechips.rocketchip.system.DefaultRV32Config.fir@24875.4]
  assign _GEN_88 = 4'he == _T_47 ? 2'h0 : _GEN_82; // @[Deinterleaver.scala 95:20:freechips.rocketchip.system.DefaultRV32Config.fir@24875.4]
  assign _GEN_89 = 4'he == _T_47 ? 4'h0 : _GEN_83; // @[Deinterleaver.scala 95:20:freechips.rocketchip.system.DefaultRV32Config.fir@24875.4]
  assign _GEN_90 = 4'he == _T_47 ? 5'h0 : _GEN_84; // @[Deinterleaver.scala 95:20:freechips.rocketchip.system.DefaultRV32Config.fir@24875.4]
  assign auto_in_aw_ready = auto_out_aw_ready; // @[LazyModule.scala 303:16:freechips.rocketchip.system.DefaultRV32Config.fir@24184.4]
  assign auto_in_w_ready = auto_out_w_ready; // @[LazyModule.scala 303:16:freechips.rocketchip.system.DefaultRV32Config.fir@24184.4]
  assign auto_in_b_valid = auto_out_b_valid; // @[LazyModule.scala 303:16:freechips.rocketchip.system.DefaultRV32Config.fir@24184.4]
  assign auto_in_b_bits_id = auto_out_b_bits_id; // @[LazyModule.scala 303:16:freechips.rocketchip.system.DefaultRV32Config.fir@24184.4]
  assign auto_in_b_bits_resp = auto_out_b_bits_resp; // @[LazyModule.scala 303:16:freechips.rocketchip.system.DefaultRV32Config.fir@24184.4]
  assign auto_in_b_bits_echo_tl_state_size = auto_out_b_bits_echo_tl_state_size; // @[LazyModule.scala 303:16:freechips.rocketchip.system.DefaultRV32Config.fir@24184.4]
  assign auto_in_b_bits_echo_tl_state_source = auto_out_b_bits_echo_tl_state_source; // @[LazyModule.scala 303:16:freechips.rocketchip.system.DefaultRV32Config.fir@24184.4]
  assign auto_in_ar_ready = auto_out_ar_ready; // @[LazyModule.scala 303:16:freechips.rocketchip.system.DefaultRV32Config.fir@24184.4]
  assign auto_in_r_valid = _T_46; // @[LazyModule.scala 303:16:freechips.rocketchip.system.DefaultRV32Config.fir@24184.4]
  assign auto_in_r_bits_id = 4'hf == _T_47 ? 4'h0 : _GEN_86; // @[LazyModule.scala 303:16:freechips.rocketchip.system.DefaultRV32Config.fir@24184.4]
  assign auto_in_r_bits_data = 4'hf == _T_47 ? 32'h0 : _GEN_87; // @[LazyModule.scala 303:16:freechips.rocketchip.system.DefaultRV32Config.fir@24184.4]
  assign auto_in_r_bits_resp = 4'hf == _T_47 ? 2'h0 : _GEN_88; // @[LazyModule.scala 303:16:freechips.rocketchip.system.DefaultRV32Config.fir@24184.4]
  assign auto_in_r_bits_echo_tl_state_size = 4'hf == _T_47 ? 4'h0 : _GEN_89; // @[LazyModule.scala 303:16:freechips.rocketchip.system.DefaultRV32Config.fir@24184.4]
  assign auto_in_r_bits_echo_tl_state_source = 4'hf == _T_47 ? 5'h0 : _GEN_90; // @[LazyModule.scala 303:16:freechips.rocketchip.system.DefaultRV32Config.fir@24184.4]
  assign auto_in_r_bits_last = 4'hf == _T_47 ? 1'h0 : _GEN_91; // @[LazyModule.scala 303:16:freechips.rocketchip.system.DefaultRV32Config.fir@24184.4]
  assign auto_out_aw_valid = auto_in_aw_valid; // @[LazyModule.scala 305:12:freechips.rocketchip.system.DefaultRV32Config.fir@24183.4]
  assign auto_out_aw_bits_id = auto_in_aw_bits_id; // @[LazyModule.scala 305:12:freechips.rocketchip.system.DefaultRV32Config.fir@24183.4]
  assign auto_out_aw_bits_addr = auto_in_aw_bits_addr; // @[LazyModule.scala 305:12:freechips.rocketchip.system.DefaultRV32Config.fir@24183.4]
  assign auto_out_aw_bits_len = auto_in_aw_bits_len; // @[LazyModule.scala 305:12:freechips.rocketchip.system.DefaultRV32Config.fir@24183.4]
  assign auto_out_aw_bits_size = auto_in_aw_bits_size; // @[LazyModule.scala 305:12:freechips.rocketchip.system.DefaultRV32Config.fir@24183.4]
  assign auto_out_aw_bits_burst = auto_in_aw_bits_burst; // @[LazyModule.scala 305:12:freechips.rocketchip.system.DefaultRV32Config.fir@24183.4]
  assign auto_out_aw_bits_lock = auto_in_aw_bits_lock; // @[LazyModule.scala 305:12:freechips.rocketchip.system.DefaultRV32Config.fir@24183.4]
  assign auto_out_aw_bits_cache = auto_in_aw_bits_cache; // @[LazyModule.scala 305:12:freechips.rocketchip.system.DefaultRV32Config.fir@24183.4]
  assign auto_out_aw_bits_prot = auto_in_aw_bits_prot; // @[LazyModule.scala 305:12:freechips.rocketchip.system.DefaultRV32Config.fir@24183.4]
  assign auto_out_aw_bits_qos = auto_in_aw_bits_qos; // @[LazyModule.scala 305:12:freechips.rocketchip.system.DefaultRV32Config.fir@24183.4]
  assign auto_out_aw_bits_echo_tl_state_size = auto_in_aw_bits_echo_tl_state_size; // @[LazyModule.scala 305:12:freechips.rocketchip.system.DefaultRV32Config.fir@24183.4]
  assign auto_out_aw_bits_echo_tl_state_source = auto_in_aw_bits_echo_tl_state_source; // @[LazyModule.scala 305:12:freechips.rocketchip.system.DefaultRV32Config.fir@24183.4]
  assign auto_out_w_valid = auto_in_w_valid; // @[LazyModule.scala 305:12:freechips.rocketchip.system.DefaultRV32Config.fir@24183.4]
  assign auto_out_w_bits_data = auto_in_w_bits_data; // @[LazyModule.scala 305:12:freechips.rocketchip.system.DefaultRV32Config.fir@24183.4]
  assign auto_out_w_bits_strb = auto_in_w_bits_strb; // @[LazyModule.scala 305:12:freechips.rocketchip.system.DefaultRV32Config.fir@24183.4]
  assign auto_out_w_bits_last = auto_in_w_bits_last; // @[LazyModule.scala 305:12:freechips.rocketchip.system.DefaultRV32Config.fir@24183.4]
  assign auto_out_b_ready = auto_in_b_ready; // @[LazyModule.scala 305:12:freechips.rocketchip.system.DefaultRV32Config.fir@24183.4]
  assign auto_out_ar_valid = auto_in_ar_valid; // @[LazyModule.scala 305:12:freechips.rocketchip.system.DefaultRV32Config.fir@24183.4]
  assign auto_out_ar_bits_id = auto_in_ar_bits_id; // @[LazyModule.scala 305:12:freechips.rocketchip.system.DefaultRV32Config.fir@24183.4]
  assign auto_out_ar_bits_addr = auto_in_ar_bits_addr; // @[LazyModule.scala 305:12:freechips.rocketchip.system.DefaultRV32Config.fir@24183.4]
  assign auto_out_ar_bits_len = auto_in_ar_bits_len; // @[LazyModule.scala 305:12:freechips.rocketchip.system.DefaultRV32Config.fir@24183.4]
  assign auto_out_ar_bits_size = auto_in_ar_bits_size; // @[LazyModule.scala 305:12:freechips.rocketchip.system.DefaultRV32Config.fir@24183.4]
  assign auto_out_ar_bits_burst = auto_in_ar_bits_burst; // @[LazyModule.scala 305:12:freechips.rocketchip.system.DefaultRV32Config.fir@24183.4]
  assign auto_out_ar_bits_lock = auto_in_ar_bits_lock; // @[LazyModule.scala 305:12:freechips.rocketchip.system.DefaultRV32Config.fir@24183.4]
  assign auto_out_ar_bits_cache = auto_in_ar_bits_cache; // @[LazyModule.scala 305:12:freechips.rocketchip.system.DefaultRV32Config.fir@24183.4]
  assign auto_out_ar_bits_prot = auto_in_ar_bits_prot; // @[LazyModule.scala 305:12:freechips.rocketchip.system.DefaultRV32Config.fir@24183.4]
  assign auto_out_ar_bits_qos = auto_in_ar_bits_qos; // @[LazyModule.scala 305:12:freechips.rocketchip.system.DefaultRV32Config.fir@24183.4]
  assign auto_out_ar_bits_echo_tl_state_size = auto_in_ar_bits_echo_tl_state_size; // @[LazyModule.scala 305:12:freechips.rocketchip.system.DefaultRV32Config.fir@24183.4]
  assign auto_out_ar_bits_echo_tl_state_source = auto_in_ar_bits_echo_tl_state_source; // @[LazyModule.scala 305:12:freechips.rocketchip.system.DefaultRV32Config.fir@24183.4]
  assign auto_out_r_ready = 4'hf == auto_out_r_bits_id ? 1'h0 : _GEN_112; // @[LazyModule.scala 305:12:freechips.rocketchip.system.DefaultRV32Config.fir@24183.4]
  assign queue_0_clock = clock; // @[:freechips.rocketchip.system.DefaultRV32Config.fir@24223.4]
  assign queue_0_reset = reset; // @[:freechips.rocketchip.system.DefaultRV32Config.fir@24224.4]
  assign queue_0_io_enq_valid = _T_52[0] & auto_out_r_valid; // @[Deinterleaver.scala 108:23:freechips.rocketchip.system.DefaultRV32Config.fir@24980.4]
  assign queue_0_io_enq_bits_id = auto_out_r_bits_id; // @[Deinterleaver.scala 109:22:freechips.rocketchip.system.DefaultRV32Config.fir@24986.4]
  assign queue_0_io_enq_bits_data = auto_out_r_bits_data; // @[Deinterleaver.scala 109:22:freechips.rocketchip.system.DefaultRV32Config.fir@24985.4]
  assign queue_0_io_enq_bits_resp = auto_out_r_bits_resp; // @[Deinterleaver.scala 109:22:freechips.rocketchip.system.DefaultRV32Config.fir@24984.4]
  assign queue_0_io_enq_bits_echo_tl_state_size = auto_out_r_bits_echo_tl_state_size; // @[Deinterleaver.scala 109:22:freechips.rocketchip.system.DefaultRV32Config.fir@24983.4]
  assign queue_0_io_enq_bits_echo_tl_state_source = auto_out_r_bits_echo_tl_state_source; // @[Deinterleaver.scala 109:22:freechips.rocketchip.system.DefaultRV32Config.fir@24982.4]
  assign queue_0_io_enq_bits_last = auto_out_r_bits_last; // @[Deinterleaver.scala 109:22:freechips.rocketchip.system.DefaultRV32Config.fir@24981.4]
  assign queue_0_io_deq_ready = _T_49[0] & _T_61; // @[Deinterleaver.scala 99:23:freechips.rocketchip.system.DefaultRV32Config.fir@24899.4]
  assign queue_1_clock = clock; // @[:freechips.rocketchip.system.DefaultRV32Config.fir@24226.4]
  assign queue_1_reset = reset; // @[:freechips.rocketchip.system.DefaultRV32Config.fir@24227.4]
  assign queue_1_io_enq_valid = _T_52[1] & auto_out_r_valid; // @[Deinterleaver.scala 108:23:freechips.rocketchip.system.DefaultRV32Config.fir@24988.4]
  assign queue_1_io_enq_bits_id = auto_out_r_bits_id; // @[Deinterleaver.scala 109:22:freechips.rocketchip.system.DefaultRV32Config.fir@24994.4]
  assign queue_1_io_enq_bits_data = auto_out_r_bits_data; // @[Deinterleaver.scala 109:22:freechips.rocketchip.system.DefaultRV32Config.fir@24993.4]
  assign queue_1_io_enq_bits_resp = auto_out_r_bits_resp; // @[Deinterleaver.scala 109:22:freechips.rocketchip.system.DefaultRV32Config.fir@24992.4]
  assign queue_1_io_enq_bits_echo_tl_state_size = auto_out_r_bits_echo_tl_state_size; // @[Deinterleaver.scala 109:22:freechips.rocketchip.system.DefaultRV32Config.fir@24991.4]
  assign queue_1_io_enq_bits_echo_tl_state_source = auto_out_r_bits_echo_tl_state_source; // @[Deinterleaver.scala 109:22:freechips.rocketchip.system.DefaultRV32Config.fir@24990.4]
  assign queue_1_io_enq_bits_last = auto_out_r_bits_last; // @[Deinterleaver.scala 109:22:freechips.rocketchip.system.DefaultRV32Config.fir@24989.4]
  assign queue_1_io_deq_ready = _T_49[1] & _T_61; // @[Deinterleaver.scala 99:23:freechips.rocketchip.system.DefaultRV32Config.fir@24902.4]
  assign queue_2_clock = clock; // @[:freechips.rocketchip.system.DefaultRV32Config.fir@24229.4]
  assign queue_2_reset = reset; // @[:freechips.rocketchip.system.DefaultRV32Config.fir@24230.4]
  assign queue_2_io_enq_valid = _T_52[2] & auto_out_r_valid; // @[Deinterleaver.scala 108:23:freechips.rocketchip.system.DefaultRV32Config.fir@24996.4]
  assign queue_2_io_enq_bits_id = auto_out_r_bits_id; // @[Deinterleaver.scala 109:22:freechips.rocketchip.system.DefaultRV32Config.fir@25002.4]
  assign queue_2_io_enq_bits_data = auto_out_r_bits_data; // @[Deinterleaver.scala 109:22:freechips.rocketchip.system.DefaultRV32Config.fir@25001.4]
  assign queue_2_io_enq_bits_resp = auto_out_r_bits_resp; // @[Deinterleaver.scala 109:22:freechips.rocketchip.system.DefaultRV32Config.fir@25000.4]
  assign queue_2_io_enq_bits_echo_tl_state_size = auto_out_r_bits_echo_tl_state_size; // @[Deinterleaver.scala 109:22:freechips.rocketchip.system.DefaultRV32Config.fir@24999.4]
  assign queue_2_io_enq_bits_echo_tl_state_source = auto_out_r_bits_echo_tl_state_source; // @[Deinterleaver.scala 109:22:freechips.rocketchip.system.DefaultRV32Config.fir@24998.4]
  assign queue_2_io_enq_bits_last = auto_out_r_bits_last; // @[Deinterleaver.scala 109:22:freechips.rocketchip.system.DefaultRV32Config.fir@24997.4]
  assign queue_2_io_deq_ready = _T_49[2] & _T_61; // @[Deinterleaver.scala 99:23:freechips.rocketchip.system.DefaultRV32Config.fir@24905.4]
  assign queue_3_clock = clock; // @[:freechips.rocketchip.system.DefaultRV32Config.fir@24232.4]
  assign queue_3_reset = reset; // @[:freechips.rocketchip.system.DefaultRV32Config.fir@24233.4]
  assign queue_3_io_enq_valid = _T_52[3] & auto_out_r_valid; // @[Deinterleaver.scala 108:23:freechips.rocketchip.system.DefaultRV32Config.fir@25004.4]
  assign queue_3_io_enq_bits_id = auto_out_r_bits_id; // @[Deinterleaver.scala 109:22:freechips.rocketchip.system.DefaultRV32Config.fir@25010.4]
  assign queue_3_io_enq_bits_data = auto_out_r_bits_data; // @[Deinterleaver.scala 109:22:freechips.rocketchip.system.DefaultRV32Config.fir@25009.4]
  assign queue_3_io_enq_bits_resp = auto_out_r_bits_resp; // @[Deinterleaver.scala 109:22:freechips.rocketchip.system.DefaultRV32Config.fir@25008.4]
  assign queue_3_io_enq_bits_echo_tl_state_size = auto_out_r_bits_echo_tl_state_size; // @[Deinterleaver.scala 109:22:freechips.rocketchip.system.DefaultRV32Config.fir@25007.4]
  assign queue_3_io_enq_bits_echo_tl_state_source = auto_out_r_bits_echo_tl_state_source; // @[Deinterleaver.scala 109:22:freechips.rocketchip.system.DefaultRV32Config.fir@25006.4]
  assign queue_3_io_enq_bits_last = auto_out_r_bits_last; // @[Deinterleaver.scala 109:22:freechips.rocketchip.system.DefaultRV32Config.fir@25005.4]
  assign queue_3_io_deq_ready = _T_49[3] & _T_61; // @[Deinterleaver.scala 99:23:freechips.rocketchip.system.DefaultRV32Config.fir@24908.4]
  assign queue_4_clock = clock; // @[:freechips.rocketchip.system.DefaultRV32Config.fir@24235.4]
  assign queue_4_reset = reset; // @[:freechips.rocketchip.system.DefaultRV32Config.fir@24236.4]
  assign queue_4_io_enq_valid = _T_52[4] & auto_out_r_valid; // @[Deinterleaver.scala 108:23:freechips.rocketchip.system.DefaultRV32Config.fir@25012.4]
  assign queue_4_io_enq_bits_id = auto_out_r_bits_id; // @[Deinterleaver.scala 109:22:freechips.rocketchip.system.DefaultRV32Config.fir@25018.4]
  assign queue_4_io_enq_bits_data = auto_out_r_bits_data; // @[Deinterleaver.scala 109:22:freechips.rocketchip.system.DefaultRV32Config.fir@25017.4]
  assign queue_4_io_enq_bits_resp = auto_out_r_bits_resp; // @[Deinterleaver.scala 109:22:freechips.rocketchip.system.DefaultRV32Config.fir@25016.4]
  assign queue_4_io_enq_bits_echo_tl_state_size = auto_out_r_bits_echo_tl_state_size; // @[Deinterleaver.scala 109:22:freechips.rocketchip.system.DefaultRV32Config.fir@25015.4]
  assign queue_4_io_enq_bits_echo_tl_state_source = auto_out_r_bits_echo_tl_state_source; // @[Deinterleaver.scala 109:22:freechips.rocketchip.system.DefaultRV32Config.fir@25014.4]
  assign queue_4_io_enq_bits_last = auto_out_r_bits_last; // @[Deinterleaver.scala 109:22:freechips.rocketchip.system.DefaultRV32Config.fir@25013.4]
  assign queue_4_io_deq_ready = _T_49[4] & _T_61; // @[Deinterleaver.scala 99:23:freechips.rocketchip.system.DefaultRV32Config.fir@24911.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_46 = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  _T_47 = _RAND_1[3:0];
  _RAND_2 = {1{`RANDOM}};
  _T_54 = _RAND_2[4:0];
  _RAND_3 = {1{`RANDOM}};
  _T_81 = _RAND_3[4:0];
  _RAND_4 = {1{`RANDOM}};
  _T_108 = _RAND_4[4:0];
  _RAND_5 = {1{`RANDOM}};
  _T_135 = _RAND_5[4:0];
  _RAND_6 = {1{`RANDOM}};
  _T_162 = _RAND_6[4:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      _T_46 <= 1'h0;
    end else if (_T_223) begin
      _T_46 <= _T_224;
    end
    _T_47 <= _GEN_1[3:0];
    if (reset) begin
      _T_54 <= 5'h0;
    end else begin
      _T_54 <= _T_67;
    end
    if (reset) begin
      _T_81 <= 5'h0;
    end else begin
      _T_81 <= _T_94;
    end
    if (reset) begin
      _T_108 <= 5'h0;
    end else begin
      _T_108 <= _T_121;
    end
    if (reset) begin
      _T_135 <= 5'h0;
    end else begin
      _T_135 <= _T_148;
    end
    if (reset) begin
      _T_162 <= 5'h0;
    end else begin
      _T_162 <= _T_175;
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_5) begin
          $fwrite(32'h80000002,"Assertion failed: ID 5 should not be used\n    at Deinterleaver.scala:53 assert(!q.enq.valid, s\"ID ${i} should not be used\")\n"); // @[Deinterleaver.scala 53:19:freechips.rocketchip.system.DefaultRV32Config.fir@24243.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_5) begin
          $fatal; // @[Deinterleaver.scala 53:19:freechips.rocketchip.system.DefaultRV32Config.fir@24244.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_9) begin
          $fwrite(32'h80000002,"Assertion failed: ID 6 should not be used\n    at Deinterleaver.scala:53 assert(!q.enq.valid, s\"ID ${i} should not be used\")\n"); // @[Deinterleaver.scala 53:19:freechips.rocketchip.system.DefaultRV32Config.fir@24269.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_9) begin
          $fatal; // @[Deinterleaver.scala 53:19:freechips.rocketchip.system.DefaultRV32Config.fir@24270.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_13) begin
          $fwrite(32'h80000002,"Assertion failed: ID 7 should not be used\n    at Deinterleaver.scala:53 assert(!q.enq.valid, s\"ID ${i} should not be used\")\n"); // @[Deinterleaver.scala 53:19:freechips.rocketchip.system.DefaultRV32Config.fir@24295.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_13) begin
          $fatal; // @[Deinterleaver.scala 53:19:freechips.rocketchip.system.DefaultRV32Config.fir@24296.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_17) begin
          $fwrite(32'h80000002,"Assertion failed: ID 8 should not be used\n    at Deinterleaver.scala:53 assert(!q.enq.valid, s\"ID ${i} should not be used\")\n"); // @[Deinterleaver.scala 53:19:freechips.rocketchip.system.DefaultRV32Config.fir@24321.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_17) begin
          $fatal; // @[Deinterleaver.scala 53:19:freechips.rocketchip.system.DefaultRV32Config.fir@24322.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_21) begin
          $fwrite(32'h80000002,"Assertion failed: ID 9 should not be used\n    at Deinterleaver.scala:53 assert(!q.enq.valid, s\"ID ${i} should not be used\")\n"); // @[Deinterleaver.scala 53:19:freechips.rocketchip.system.DefaultRV32Config.fir@24347.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_21) begin
          $fatal; // @[Deinterleaver.scala 53:19:freechips.rocketchip.system.DefaultRV32Config.fir@24348.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_25) begin
          $fwrite(32'h80000002,"Assertion failed: ID 10 should not be used\n    at Deinterleaver.scala:53 assert(!q.enq.valid, s\"ID ${i} should not be used\")\n"); // @[Deinterleaver.scala 53:19:freechips.rocketchip.system.DefaultRV32Config.fir@24373.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_25) begin
          $fatal; // @[Deinterleaver.scala 53:19:freechips.rocketchip.system.DefaultRV32Config.fir@24374.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_29) begin
          $fwrite(32'h80000002,"Assertion failed: ID 11 should not be used\n    at Deinterleaver.scala:53 assert(!q.enq.valid, s\"ID ${i} should not be used\")\n"); // @[Deinterleaver.scala 53:19:freechips.rocketchip.system.DefaultRV32Config.fir@24399.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_29) begin
          $fatal; // @[Deinterleaver.scala 53:19:freechips.rocketchip.system.DefaultRV32Config.fir@24400.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_33) begin
          $fwrite(32'h80000002,"Assertion failed: ID 12 should not be used\n    at Deinterleaver.scala:53 assert(!q.enq.valid, s\"ID ${i} should not be used\")\n"); // @[Deinterleaver.scala 53:19:freechips.rocketchip.system.DefaultRV32Config.fir@24425.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_33) begin
          $fatal; // @[Deinterleaver.scala 53:19:freechips.rocketchip.system.DefaultRV32Config.fir@24426.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_37) begin
          $fwrite(32'h80000002,"Assertion failed: ID 13 should not be used\n    at Deinterleaver.scala:53 assert(!q.enq.valid, s\"ID ${i} should not be used\")\n"); // @[Deinterleaver.scala 53:19:freechips.rocketchip.system.DefaultRV32Config.fir@24451.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_37) begin
          $fatal; // @[Deinterleaver.scala 53:19:freechips.rocketchip.system.DefaultRV32Config.fir@24452.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_41) begin
          $fwrite(32'h80000002,"Assertion failed: ID 14 should not be used\n    at Deinterleaver.scala:53 assert(!q.enq.valid, s\"ID ${i} should not be used\")\n"); // @[Deinterleaver.scala 53:19:freechips.rocketchip.system.DefaultRV32Config.fir@24477.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_41) begin
          $fatal; // @[Deinterleaver.scala 53:19:freechips.rocketchip.system.DefaultRV32Config.fir@24478.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_45) begin
          $fwrite(32'h80000002,"Assertion failed: ID 15 should not be used\n    at Deinterleaver.scala:53 assert(!q.enq.valid, s\"ID ${i} should not be used\")\n"); // @[Deinterleaver.scala 53:19:freechips.rocketchip.system.DefaultRV32Config.fir@24503.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_45) begin
          $fatal; // @[Deinterleaver.scala 53:19:freechips.rocketchip.system.DefaultRV32Config.fir@24504.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_73) begin
          $fwrite(32'h80000002,"Assertion failed\n    at Deinterleaver.scala:79 assert (!dec || count =/= 0.U)\n"); // @[Deinterleaver.scala 79:20:freechips.rocketchip.system.DefaultRV32Config.fir@24554.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_73) begin
          $fatal; // @[Deinterleaver.scala 79:20:freechips.rocketchip.system.DefaultRV32Config.fir@24555.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_79) begin
          $fwrite(32'h80000002,"Assertion failed\n    at Deinterleaver.scala:80 assert (!inc || count =/= beats.U)\n"); // @[Deinterleaver.scala 80:20:freechips.rocketchip.system.DefaultRV32Config.fir@24564.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_79) begin
          $fatal; // @[Deinterleaver.scala 80:20:freechips.rocketchip.system.DefaultRV32Config.fir@24565.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_100) begin
          $fwrite(32'h80000002,"Assertion failed\n    at Deinterleaver.scala:79 assert (!dec || count =/= 0.U)\n"); // @[Deinterleaver.scala 79:20:freechips.rocketchip.system.DefaultRV32Config.fir@24591.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_100) begin
          $fatal; // @[Deinterleaver.scala 79:20:freechips.rocketchip.system.DefaultRV32Config.fir@24592.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_106) begin
          $fwrite(32'h80000002,"Assertion failed\n    at Deinterleaver.scala:80 assert (!inc || count =/= beats.U)\n"); // @[Deinterleaver.scala 80:20:freechips.rocketchip.system.DefaultRV32Config.fir@24601.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_106) begin
          $fatal; // @[Deinterleaver.scala 80:20:freechips.rocketchip.system.DefaultRV32Config.fir@24602.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_127) begin
          $fwrite(32'h80000002,"Assertion failed\n    at Deinterleaver.scala:79 assert (!dec || count =/= 0.U)\n"); // @[Deinterleaver.scala 79:20:freechips.rocketchip.system.DefaultRV32Config.fir@24628.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_127) begin
          $fatal; // @[Deinterleaver.scala 79:20:freechips.rocketchip.system.DefaultRV32Config.fir@24629.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_133) begin
          $fwrite(32'h80000002,"Assertion failed\n    at Deinterleaver.scala:80 assert (!inc || count =/= beats.U)\n"); // @[Deinterleaver.scala 80:20:freechips.rocketchip.system.DefaultRV32Config.fir@24638.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_133) begin
          $fatal; // @[Deinterleaver.scala 80:20:freechips.rocketchip.system.DefaultRV32Config.fir@24639.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_154) begin
          $fwrite(32'h80000002,"Assertion failed\n    at Deinterleaver.scala:79 assert (!dec || count =/= 0.U)\n"); // @[Deinterleaver.scala 79:20:freechips.rocketchip.system.DefaultRV32Config.fir@24665.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_154) begin
          $fatal; // @[Deinterleaver.scala 79:20:freechips.rocketchip.system.DefaultRV32Config.fir@24666.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_160) begin
          $fwrite(32'h80000002,"Assertion failed\n    at Deinterleaver.scala:80 assert (!inc || count =/= beats.U)\n"); // @[Deinterleaver.scala 80:20:freechips.rocketchip.system.DefaultRV32Config.fir@24675.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_160) begin
          $fatal; // @[Deinterleaver.scala 80:20:freechips.rocketchip.system.DefaultRV32Config.fir@24676.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_181) begin
          $fwrite(32'h80000002,"Assertion failed\n    at Deinterleaver.scala:79 assert (!dec || count =/= 0.U)\n"); // @[Deinterleaver.scala 79:20:freechips.rocketchip.system.DefaultRV32Config.fir@24702.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_181) begin
          $fatal; // @[Deinterleaver.scala 79:20:freechips.rocketchip.system.DefaultRV32Config.fir@24703.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_187) begin
          $fwrite(32'h80000002,"Assertion failed\n    at Deinterleaver.scala:80 assert (!inc || count =/= beats.U)\n"); // @[Deinterleaver.scala 80:20:freechips.rocketchip.system.DefaultRV32Config.fir@24712.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_187) begin
          $fatal; // @[Deinterleaver.scala 80:20:freechips.rocketchip.system.DefaultRV32Config.fir@24713.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
  end
endmodule
