module OptimizationBarrier( // @[:freechips.rocketchip.system.DefaultRV32Config.fir@175626.2]
  input  [19:0] io_x_ppn, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@175629.4]
  input         io_x_u, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@175629.4]
  input         io_x_ae, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@175629.4]
  input         io_x_sw, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@175629.4]
  input         io_x_sx, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@175629.4]
  input         io_x_sr, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@175629.4]
  input         io_x_pw, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@175629.4]
  input         io_x_px, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@175629.4]
  input         io_x_pr, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@175629.4]
  input         io_x_ppp, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@175629.4]
  input         io_x_pal, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@175629.4]
  input         io_x_paa, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@175629.4]
  input         io_x_eff, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@175629.4]
  input         io_x_c, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@175629.4]
  output [19:0] io_y_ppn, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@175629.4]
  output        io_y_u, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@175629.4]
  output        io_y_ae, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@175629.4]
  output        io_y_sw, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@175629.4]
  output        io_y_sx, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@175629.4]
  output        io_y_sr, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@175629.4]
  output        io_y_pw, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@175629.4]
  output        io_y_px, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@175629.4]
  output        io_y_pr, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@175629.4]
  output        io_y_ppp, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@175629.4]
  output        io_y_pal, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@175629.4]
  output        io_y_paa, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@175629.4]
  output        io_y_eff, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@175629.4]
  output        io_y_c // @[:freechips.rocketchip.system.DefaultRV32Config.fir@175629.4]
);
  assign io_y_ppn = io_x_ppn; // @[package.scala 236:12:freechips.rocketchip.system.DefaultRV32Config.fir@175634.4]
  assign io_y_u = io_x_u; // @[package.scala 236:12:freechips.rocketchip.system.DefaultRV32Config.fir@175634.4]
  assign io_y_ae = io_x_ae; // @[package.scala 236:12:freechips.rocketchip.system.DefaultRV32Config.fir@175634.4]
  assign io_y_sw = io_x_sw; // @[package.scala 236:12:freechips.rocketchip.system.DefaultRV32Config.fir@175634.4]
  assign io_y_sx = io_x_sx; // @[package.scala 236:12:freechips.rocketchip.system.DefaultRV32Config.fir@175634.4]
  assign io_y_sr = io_x_sr; // @[package.scala 236:12:freechips.rocketchip.system.DefaultRV32Config.fir@175634.4]
  assign io_y_pw = io_x_pw; // @[package.scala 236:12:freechips.rocketchip.system.DefaultRV32Config.fir@175634.4]
  assign io_y_px = io_x_px; // @[package.scala 236:12:freechips.rocketchip.system.DefaultRV32Config.fir@175634.4]
  assign io_y_pr = io_x_pr; // @[package.scala 236:12:freechips.rocketchip.system.DefaultRV32Config.fir@175634.4]
  assign io_y_ppp = io_x_ppp; // @[package.scala 236:12:freechips.rocketchip.system.DefaultRV32Config.fir@175634.4]
  assign io_y_pal = io_x_pal; // @[package.scala 236:12:freechips.rocketchip.system.DefaultRV32Config.fir@175634.4]
  assign io_y_paa = io_x_paa; // @[package.scala 236:12:freechips.rocketchip.system.DefaultRV32Config.fir@175634.4]
  assign io_y_eff = io_x_eff; // @[package.scala 236:12:freechips.rocketchip.system.DefaultRV32Config.fir@175634.4]
  assign io_y_c = io_x_c; // @[package.scala 236:12:freechips.rocketchip.system.DefaultRV32Config.fir@175634.4]
endmodule
