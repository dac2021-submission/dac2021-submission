module IntXbar( // @[:freechips.rocketchip.system.DefaultRV32Config.fir@3.2]
  input   auto_int_in_0, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@6.4]
  input   auto_int_in_1, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@6.4]
  output  auto_int_out_0, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@6.4]
  output  auto_int_out_1 // @[:freechips.rocketchip.system.DefaultRV32Config.fir@6.4]
);
  assign auto_int_out_0 = auto_int_in_0; // @[LazyModule.scala 305:12:freechips.rocketchip.system.DefaultRV32Config.fir@15.4]
  assign auto_int_out_1 = auto_int_in_1; // @[LazyModule.scala 305:12:freechips.rocketchip.system.DefaultRV32Config.fir@15.4]
endmodule
