module FPUDecoder( // @[:freechips.rocketchip.system.DefaultRV32Config.fir@210598.2]
  input  [31:0] io_inst, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@210601.4]
  output        io_sigs_wen, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@210601.4]
  output        io_sigs_ren1, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@210601.4]
  output        io_sigs_ren2, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@210601.4]
  output        io_sigs_ren3, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@210601.4]
  output        io_sigs_swap12, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@210601.4]
  output        io_sigs_swap23, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@210601.4]
  output        io_sigs_singleOut, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@210601.4]
  output        io_sigs_fromint, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@210601.4]
  output        io_sigs_toint, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@210601.4]
  output        io_sigs_fastpipe, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@210601.4]
  output        io_sigs_fma, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@210601.4]
  output        io_sigs_div, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@210601.4]
  output        io_sigs_sqrt, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@210601.4]
  output        io_sigs_wflags // @[:freechips.rocketchip.system.DefaultRV32Config.fir@210601.4]
);
  wire [31:0] _T; // @[Decode.scala 14:65:freechips.rocketchip.system.DefaultRV32Config.fir@210606.4]
  wire [31:0] _T_2; // @[Decode.scala 14:65:freechips.rocketchip.system.DefaultRV32Config.fir@210609.4]
  wire  _T_3; // @[Decode.scala 14:121:freechips.rocketchip.system.DefaultRV32Config.fir@210610.4]
  wire [31:0] _T_4; // @[Decode.scala 14:65:freechips.rocketchip.system.DefaultRV32Config.fir@210611.4]
  wire  _T_5; // @[Decode.scala 14:121:freechips.rocketchip.system.DefaultRV32Config.fir@210612.4]
  wire [31:0] _T_6; // @[Decode.scala 14:65:freechips.rocketchip.system.DefaultRV32Config.fir@210613.4]
  wire  _T_7; // @[Decode.scala 14:121:freechips.rocketchip.system.DefaultRV32Config.fir@210614.4]
  wire  _T_9; // @[Decode.scala 15:30:freechips.rocketchip.system.DefaultRV32Config.fir@210616.4]
  wire [31:0] _T_10; // @[Decode.scala 14:65:freechips.rocketchip.system.DefaultRV32Config.fir@210618.4]
  wire  _T_11; // @[Decode.scala 14:121:freechips.rocketchip.system.DefaultRV32Config.fir@210619.4]
  wire [31:0] _T_12; // @[Decode.scala 14:65:freechips.rocketchip.system.DefaultRV32Config.fir@210620.4]
  wire  _T_13; // @[Decode.scala 14:121:freechips.rocketchip.system.DefaultRV32Config.fir@210621.4]
  wire [31:0] _T_14; // @[Decode.scala 14:65:freechips.rocketchip.system.DefaultRV32Config.fir@210622.4]
  wire  decoder_4; // @[Decode.scala 14:121:freechips.rocketchip.system.DefaultRV32Config.fir@210623.4]
  wire  _T_17; // @[Decode.scala 15:30:freechips.rocketchip.system.DefaultRV32Config.fir@210625.4]
  wire [31:0] _T_18; // @[Decode.scala 14:65:freechips.rocketchip.system.DefaultRV32Config.fir@210627.4]
  wire  _T_19; // @[Decode.scala 14:121:freechips.rocketchip.system.DefaultRV32Config.fir@210628.4]
  wire [31:0] _T_20; // @[Decode.scala 14:65:freechips.rocketchip.system.DefaultRV32Config.fir@210629.4]
  wire  _T_21; // @[Decode.scala 14:121:freechips.rocketchip.system.DefaultRV32Config.fir@210630.4]
  wire  _T_23; // @[Decode.scala 15:30:freechips.rocketchip.system.DefaultRV32Config.fir@210632.4]
  wire [31:0] _T_24; // @[Decode.scala 14:65:freechips.rocketchip.system.DefaultRV32Config.fir@210636.4]
  wire [31:0] _T_38; // @[Decode.scala 14:65:freechips.rocketchip.system.DefaultRV32Config.fir@210652.4]
  wire  _T_39; // @[Decode.scala 14:121:freechips.rocketchip.system.DefaultRV32Config.fir@210653.4]
  wire [31:0] _T_40; // @[Decode.scala 14:65:freechips.rocketchip.system.DefaultRV32Config.fir@210654.4]
  wire  _T_41; // @[Decode.scala 14:121:freechips.rocketchip.system.DefaultRV32Config.fir@210655.4]
  wire [31:0] _T_42; // @[Decode.scala 14:65:freechips.rocketchip.system.DefaultRV32Config.fir@210656.4]
  wire  _T_43; // @[Decode.scala 14:121:freechips.rocketchip.system.DefaultRV32Config.fir@210657.4]
  wire  _T_45; // @[Decode.scala 15:30:freechips.rocketchip.system.DefaultRV32Config.fir@210659.4]
  wire [31:0] _T_46; // @[Decode.scala 14:65:freechips.rocketchip.system.DefaultRV32Config.fir@210661.4]
  wire  _T_49; // @[Decode.scala 14:121:freechips.rocketchip.system.DefaultRV32Config.fir@210665.4]
  wire [31:0] _T_51; // @[Decode.scala 14:65:freechips.rocketchip.system.DefaultRV32Config.fir@210668.4]
  wire [31:0] _T_53; // @[Decode.scala 14:65:freechips.rocketchip.system.DefaultRV32Config.fir@210671.4]
  wire  _T_54; // @[Decode.scala 14:121:freechips.rocketchip.system.DefaultRV32Config.fir@210672.4]
  wire [31:0] _T_55; // @[Decode.scala 14:65:freechips.rocketchip.system.DefaultRV32Config.fir@210673.4]
  wire  _T_56; // @[Decode.scala 14:121:freechips.rocketchip.system.DefaultRV32Config.fir@210674.4]
  wire  _T_58; // @[Decode.scala 15:30:freechips.rocketchip.system.DefaultRV32Config.fir@210676.4]
  wire [31:0] _T_59; // @[Decode.scala 14:65:freechips.rocketchip.system.DefaultRV32Config.fir@210678.4]
  wire [31:0] _T_61; // @[Decode.scala 14:65:freechips.rocketchip.system.DefaultRV32Config.fir@210681.4]
  wire [31:0] _T_63; // @[Decode.scala 14:65:freechips.rocketchip.system.DefaultRV32Config.fir@210684.4]
  wire  _T_64; // @[Decode.scala 14:121:freechips.rocketchip.system.DefaultRV32Config.fir@210685.4]
  wire [31:0] _T_65; // @[Decode.scala 14:65:freechips.rocketchip.system.DefaultRV32Config.fir@210686.4]
  wire  _T_66; // @[Decode.scala 14:121:freechips.rocketchip.system.DefaultRV32Config.fir@210687.4]
  wire [31:0] _T_67; // @[Decode.scala 14:65:freechips.rocketchip.system.DefaultRV32Config.fir@210688.4]
  wire  _T_68; // @[Decode.scala 14:121:freechips.rocketchip.system.DefaultRV32Config.fir@210689.4]
  wire  _T_70; // @[Decode.scala 15:30:freechips.rocketchip.system.DefaultRV32Config.fir@210691.4]
  wire  _T_71; // @[Decode.scala 15:30:freechips.rocketchip.system.DefaultRV32Config.fir@210692.4]
  assign _T = io_inst & 32'h40; // @[Decode.scala 14:65:freechips.rocketchip.system.DefaultRV32Config.fir@210606.4]
  assign _T_2 = io_inst & 32'h80000020; // @[Decode.scala 14:65:freechips.rocketchip.system.DefaultRV32Config.fir@210609.4]
  assign _T_3 = _T_2 == 32'h0; // @[Decode.scala 14:121:freechips.rocketchip.system.DefaultRV32Config.fir@210610.4]
  assign _T_4 = io_inst & 32'h30; // @[Decode.scala 14:65:freechips.rocketchip.system.DefaultRV32Config.fir@210611.4]
  assign _T_5 = _T_4 == 32'h0; // @[Decode.scala 14:121:freechips.rocketchip.system.DefaultRV32Config.fir@210612.4]
  assign _T_6 = io_inst & 32'h10000020; // @[Decode.scala 14:65:freechips.rocketchip.system.DefaultRV32Config.fir@210613.4]
  assign _T_7 = _T_6 == 32'h10000000; // @[Decode.scala 14:121:freechips.rocketchip.system.DefaultRV32Config.fir@210614.4]
  assign _T_9 = _T_3 | _T_5; // @[Decode.scala 15:30:freechips.rocketchip.system.DefaultRV32Config.fir@210616.4]
  assign _T_10 = io_inst & 32'h80000004; // @[Decode.scala 14:65:freechips.rocketchip.system.DefaultRV32Config.fir@210618.4]
  assign _T_11 = _T_10 == 32'h0; // @[Decode.scala 14:121:freechips.rocketchip.system.DefaultRV32Config.fir@210619.4]
  assign _T_12 = io_inst & 32'h10000004; // @[Decode.scala 14:65:freechips.rocketchip.system.DefaultRV32Config.fir@210620.4]
  assign _T_13 = _T_12 == 32'h0; // @[Decode.scala 14:121:freechips.rocketchip.system.DefaultRV32Config.fir@210621.4]
  assign _T_14 = io_inst & 32'h50; // @[Decode.scala 14:65:freechips.rocketchip.system.DefaultRV32Config.fir@210622.4]
  assign decoder_4 = _T_14 == 32'h40; // @[Decode.scala 14:121:freechips.rocketchip.system.DefaultRV32Config.fir@210623.4]
  assign _T_17 = _T_11 | _T_13; // @[Decode.scala 15:30:freechips.rocketchip.system.DefaultRV32Config.fir@210625.4]
  assign _T_18 = io_inst & 32'h40000004; // @[Decode.scala 14:65:freechips.rocketchip.system.DefaultRV32Config.fir@210627.4]
  assign _T_19 = _T_18 == 32'h0; // @[Decode.scala 14:121:freechips.rocketchip.system.DefaultRV32Config.fir@210628.4]
  assign _T_20 = io_inst & 32'h20; // @[Decode.scala 14:65:freechips.rocketchip.system.DefaultRV32Config.fir@210629.4]
  assign _T_21 = _T_20 == 32'h20; // @[Decode.scala 14:121:freechips.rocketchip.system.DefaultRV32Config.fir@210630.4]
  assign _T_23 = _T_19 | _T_21; // @[Decode.scala 15:30:freechips.rocketchip.system.DefaultRV32Config.fir@210632.4]
  assign _T_24 = io_inst & 32'h30000010; // @[Decode.scala 14:65:freechips.rocketchip.system.DefaultRV32Config.fir@210636.4]
  assign _T_38 = io_inst & 32'h20000000; // @[Decode.scala 14:65:freechips.rocketchip.system.DefaultRV32Config.fir@210652.4]
  assign _T_39 = _T_38 == 32'h0; // @[Decode.scala 14:121:freechips.rocketchip.system.DefaultRV32Config.fir@210653.4]
  assign _T_40 = io_inst & 32'h10000000; // @[Decode.scala 14:65:freechips.rocketchip.system.DefaultRV32Config.fir@210654.4]
  assign _T_41 = _T_40 == 32'h0; // @[Decode.scala 14:121:freechips.rocketchip.system.DefaultRV32Config.fir@210655.4]
  assign _T_42 = io_inst & 32'h10; // @[Decode.scala 14:65:freechips.rocketchip.system.DefaultRV32Config.fir@210656.4]
  assign _T_43 = _T_42 == 32'h0; // @[Decode.scala 14:121:freechips.rocketchip.system.DefaultRV32Config.fir@210657.4]
  assign _T_45 = _T_39 | _T_41; // @[Decode.scala 15:30:freechips.rocketchip.system.DefaultRV32Config.fir@210659.4]
  assign _T_46 = io_inst & 32'h90000010; // @[Decode.scala 14:65:freechips.rocketchip.system.DefaultRV32Config.fir@210661.4]
  assign _T_49 = _T_46 == 32'h80000010; // @[Decode.scala 14:121:freechips.rocketchip.system.DefaultRV32Config.fir@210665.4]
  assign _T_51 = io_inst & 32'ha0000010; // @[Decode.scala 14:65:freechips.rocketchip.system.DefaultRV32Config.fir@210668.4]
  assign _T_53 = io_inst & 32'hb0000004; // @[Decode.scala 14:65:freechips.rocketchip.system.DefaultRV32Config.fir@210671.4]
  assign _T_54 = _T_53 == 32'h0; // @[Decode.scala 14:121:freechips.rocketchip.system.DefaultRV32Config.fir@210672.4]
  assign _T_55 = io_inst & 32'ha8000004; // @[Decode.scala 14:65:freechips.rocketchip.system.DefaultRV32Config.fir@210673.4]
  assign _T_56 = _T_55 == 32'h0; // @[Decode.scala 14:121:freechips.rocketchip.system.DefaultRV32Config.fir@210674.4]
  assign _T_58 = _T_54 | _T_56; // @[Decode.scala 15:30:freechips.rocketchip.system.DefaultRV32Config.fir@210676.4]
  assign _T_59 = io_inst & 32'h58000010; // @[Decode.scala 14:65:freechips.rocketchip.system.DefaultRV32Config.fir@210678.4]
  assign _T_61 = io_inst & 32'hc0000010; // @[Decode.scala 14:65:freechips.rocketchip.system.DefaultRV32Config.fir@210681.4]
  assign _T_63 = io_inst & 32'h20000004; // @[Decode.scala 14:65:freechips.rocketchip.system.DefaultRV32Config.fir@210684.4]
  assign _T_64 = _T_63 == 32'h0; // @[Decode.scala 14:121:freechips.rocketchip.system.DefaultRV32Config.fir@210685.4]
  assign _T_65 = io_inst & 32'h8002000; // @[Decode.scala 14:65:freechips.rocketchip.system.DefaultRV32Config.fir@210686.4]
  assign _T_66 = _T_65 == 32'h8000000; // @[Decode.scala 14:121:freechips.rocketchip.system.DefaultRV32Config.fir@210687.4]
  assign _T_67 = io_inst & 32'hc0000004; // @[Decode.scala 14:65:freechips.rocketchip.system.DefaultRV32Config.fir@210688.4]
  assign _T_68 = _T_67 == 32'h80000000; // @[Decode.scala 14:121:freechips.rocketchip.system.DefaultRV32Config.fir@210689.4]
  assign _T_70 = _T_64 | decoder_4; // @[Decode.scala 15:30:freechips.rocketchip.system.DefaultRV32Config.fir@210691.4]
  assign _T_71 = _T_70 | _T_66; // @[Decode.scala 15:30:freechips.rocketchip.system.DefaultRV32Config.fir@210692.4]
  assign io_sigs_wen = _T_9 | _T_7; // @[FPU.scala 135:40:freechips.rocketchip.system.DefaultRV32Config.fir@210695.4]
  assign io_sigs_ren1 = _T_17 | decoder_4; // @[FPU.scala 135:40:freechips.rocketchip.system.DefaultRV32Config.fir@210696.4]
  assign io_sigs_ren2 = _T_23 | decoder_4; // @[FPU.scala 135:40:freechips.rocketchip.system.DefaultRV32Config.fir@210697.4]
  assign io_sigs_ren3 = _T_14 == 32'h40; // @[FPU.scala 135:40:freechips.rocketchip.system.DefaultRV32Config.fir@210698.4]
  assign io_sigs_swap12 = _T == 32'h0; // @[FPU.scala 135:40:freechips.rocketchip.system.DefaultRV32Config.fir@210699.4]
  assign io_sigs_swap23 = _T_24 == 32'h10; // @[FPU.scala 135:40:freechips.rocketchip.system.DefaultRV32Config.fir@210700.4]
  assign io_sigs_singleOut = _T_45 | _T_43; // @[FPU.scala 135:40:freechips.rocketchip.system.DefaultRV32Config.fir@210702.4]
  assign io_sigs_fromint = _T_46 == 32'h90000010; // @[FPU.scala 135:40:freechips.rocketchip.system.DefaultRV32Config.fir@210703.4]
  assign io_sigs_toint = _T_21 | _T_49; // @[FPU.scala 135:40:freechips.rocketchip.system.DefaultRV32Config.fir@210704.4]
  assign io_sigs_fastpipe = _T_51 == 32'h20000010; // @[FPU.scala 135:40:freechips.rocketchip.system.DefaultRV32Config.fir@210705.4]
  assign io_sigs_fma = _T_58 | decoder_4; // @[FPU.scala 135:40:freechips.rocketchip.system.DefaultRV32Config.fir@210706.4]
  assign io_sigs_div = _T_59 == 32'h18000010; // @[FPU.scala 135:40:freechips.rocketchip.system.DefaultRV32Config.fir@210707.4]
  assign io_sigs_sqrt = _T_61 == 32'h40000010; // @[FPU.scala 135:40:freechips.rocketchip.system.DefaultRV32Config.fir@210708.4]
  assign io_sigs_wflags = _T_71 | _T_68; // @[FPU.scala 135:40:freechips.rocketchip.system.DefaultRV32Config.fir@210709.4]
endmodule
