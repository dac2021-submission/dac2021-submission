module TLMonitor_46( // @[:freechips.rocketchip.system.DefaultRV32Config.fir@169948.2]
  input         clock, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@169949.4]
  input         reset, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@169950.4]
  input         io_in_a_ready, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@169951.4]
  input         io_in_a_valid, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@169951.4]
  input  [2:0]  io_in_a_bits_opcode, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@169951.4]
  input  [2:0]  io_in_a_bits_param, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@169951.4]
  input  [3:0]  io_in_a_bits_size, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@169951.4]
  input         io_in_a_bits_source, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@169951.4]
  input  [31:0] io_in_a_bits_address, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@169951.4]
  input  [3:0]  io_in_a_bits_mask, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@169951.4]
  input         io_in_b_ready, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@169951.4]
  input         io_in_b_valid, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@169951.4]
  input  [2:0]  io_in_b_bits_opcode, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@169951.4]
  input  [1:0]  io_in_b_bits_param, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@169951.4]
  input  [3:0]  io_in_b_bits_size, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@169951.4]
  input         io_in_b_bits_source, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@169951.4]
  input  [31:0] io_in_b_bits_address, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@169951.4]
  input  [3:0]  io_in_b_bits_mask, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@169951.4]
  input         io_in_b_bits_corrupt, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@169951.4]
  input         io_in_c_ready, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@169951.4]
  input         io_in_c_valid, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@169951.4]
  input  [2:0]  io_in_c_bits_opcode, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@169951.4]
  input  [2:0]  io_in_c_bits_param, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@169951.4]
  input  [3:0]  io_in_c_bits_size, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@169951.4]
  input         io_in_c_bits_source, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@169951.4]
  input  [31:0] io_in_c_bits_address, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@169951.4]
  input         io_in_d_ready, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@169951.4]
  input         io_in_d_valid, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@169951.4]
  input  [2:0]  io_in_d_bits_opcode, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@169951.4]
  input  [1:0]  io_in_d_bits_param, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@169951.4]
  input  [3:0]  io_in_d_bits_size, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@169951.4]
  input         io_in_d_bits_source, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@169951.4]
  input  [1:0]  io_in_d_bits_sink, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@169951.4]
  input         io_in_d_bits_denied, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@169951.4]
  input         io_in_d_bits_corrupt, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@169951.4]
  input         io_in_e_ready, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@169951.4]
  input         io_in_e_valid, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@169951.4]
  input  [1:0]  io_in_e_bits_sink // @[:freechips.rocketchip.system.DefaultRV32Config.fir@169951.4]
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
`endif // RANDOMIZE_REG_INIT
  wire [31:0] plusarg_reader_out; // @[PlusArg.scala 80:11:freechips.rocketchip.system.DefaultRV32Config.fir@172754.4]
  wire  _T_4; // @[Parameters.scala 47:9:freechips.rocketchip.system.DefaultRV32Config.fir@169962.6]
  wire  _T_7; // @[Parameters.scala 924:46:freechips.rocketchip.system.DefaultRV32Config.fir@169968.6]
  wire [26:0] _T_9; // @[package.scala 207:77:freechips.rocketchip.system.DefaultRV32Config.fir@169970.6]
  wire [11:0] _T_11; // @[package.scala 207:46:freechips.rocketchip.system.DefaultRV32Config.fir@169972.6]
  wire [31:0] _GEN_71; // @[Edges.scala 22:16:freechips.rocketchip.system.DefaultRV32Config.fir@169973.6]
  wire [31:0] _T_12; // @[Edges.scala 22:16:freechips.rocketchip.system.DefaultRV32Config.fir@169973.6]
  wire  _T_13; // @[Edges.scala 22:24:freechips.rocketchip.system.DefaultRV32Config.fir@169974.6]
  wire [1:0] _T_16; // @[OneHot.scala 65:12:freechips.rocketchip.system.DefaultRV32Config.fir@169977.6]
  wire [1:0] _T_18; // @[Misc.scala 201:81:freechips.rocketchip.system.DefaultRV32Config.fir@169979.6]
  wire  _T_19; // @[Misc.scala 205:21:freechips.rocketchip.system.DefaultRV32Config.fir@169980.6]
  wire  _T_22; // @[Misc.scala 210:20:freechips.rocketchip.system.DefaultRV32Config.fir@169983.6]
  wire  _T_24; // @[Misc.scala 214:38:freechips.rocketchip.system.DefaultRV32Config.fir@169985.6]
  wire  _T_25; // @[Misc.scala 214:29:freechips.rocketchip.system.DefaultRV32Config.fir@169986.6]
  wire  _T_27; // @[Misc.scala 214:38:freechips.rocketchip.system.DefaultRV32Config.fir@169988.6]
  wire  _T_28; // @[Misc.scala 214:29:freechips.rocketchip.system.DefaultRV32Config.fir@169989.6]
  wire  _T_31; // @[Misc.scala 210:20:freechips.rocketchip.system.DefaultRV32Config.fir@169992.6]
  wire  _T_32; // @[Misc.scala 213:27:freechips.rocketchip.system.DefaultRV32Config.fir@169993.6]
  wire  _T_33; // @[Misc.scala 214:38:freechips.rocketchip.system.DefaultRV32Config.fir@169994.6]
  wire  _T_34; // @[Misc.scala 214:29:freechips.rocketchip.system.DefaultRV32Config.fir@169995.6]
  wire  _T_35; // @[Misc.scala 213:27:freechips.rocketchip.system.DefaultRV32Config.fir@169996.6]
  wire  _T_36; // @[Misc.scala 214:38:freechips.rocketchip.system.DefaultRV32Config.fir@169997.6]
  wire  _T_37; // @[Misc.scala 214:29:freechips.rocketchip.system.DefaultRV32Config.fir@169998.6]
  wire  _T_38; // @[Misc.scala 213:27:freechips.rocketchip.system.DefaultRV32Config.fir@169999.6]
  wire  _T_39; // @[Misc.scala 214:38:freechips.rocketchip.system.DefaultRV32Config.fir@170000.6]
  wire  _T_40; // @[Misc.scala 214:29:freechips.rocketchip.system.DefaultRV32Config.fir@170001.6]
  wire  _T_41; // @[Misc.scala 213:27:freechips.rocketchip.system.DefaultRV32Config.fir@170002.6]
  wire  _T_42; // @[Misc.scala 214:38:freechips.rocketchip.system.DefaultRV32Config.fir@170003.6]
  wire  _T_43; // @[Misc.scala 214:29:freechips.rocketchip.system.DefaultRV32Config.fir@170004.6]
  wire [3:0] _T_46; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@170007.6]
  wire [32:0] _T_50; // @[Parameters.scala 137:49:freechips.rocketchip.system.DefaultRV32Config.fir@170011.6]
  wire  _T_67; // @[Monitor.scala 79:25:freechips.rocketchip.system.DefaultRV32Config.fir@170032.6]
  wire [32:0] _T_72; // @[Parameters.scala 137:52:freechips.rocketchip.system.DefaultRV32Config.fir@170038.8]
  wire  _T_73; // @[Parameters.scala 137:67:freechips.rocketchip.system.DefaultRV32Config.fir@170039.8]
  wire [31:0] _T_74; // @[Parameters.scala 137:31:freechips.rocketchip.system.DefaultRV32Config.fir@170040.8]
  wire [32:0] _T_75; // @[Parameters.scala 137:49:freechips.rocketchip.system.DefaultRV32Config.fir@170041.8]
  wire [32:0] _T_77; // @[Parameters.scala 137:52:freechips.rocketchip.system.DefaultRV32Config.fir@170043.8]
  wire  _T_78; // @[Parameters.scala 137:67:freechips.rocketchip.system.DefaultRV32Config.fir@170044.8]
  wire [31:0] _T_79; // @[Parameters.scala 137:31:freechips.rocketchip.system.DefaultRV32Config.fir@170045.8]
  wire [32:0] _T_80; // @[Parameters.scala 137:49:freechips.rocketchip.system.DefaultRV32Config.fir@170046.8]
  wire [32:0] _T_82; // @[Parameters.scala 137:52:freechips.rocketchip.system.DefaultRV32Config.fir@170048.8]
  wire  _T_83; // @[Parameters.scala 137:67:freechips.rocketchip.system.DefaultRV32Config.fir@170049.8]
  wire [31:0] _T_84; // @[Parameters.scala 137:31:freechips.rocketchip.system.DefaultRV32Config.fir@170050.8]
  wire [32:0] _T_85; // @[Parameters.scala 137:49:freechips.rocketchip.system.DefaultRV32Config.fir@170051.8]
  wire [32:0] _T_87; // @[Parameters.scala 137:52:freechips.rocketchip.system.DefaultRV32Config.fir@170053.8]
  wire  _T_88; // @[Parameters.scala 137:67:freechips.rocketchip.system.DefaultRV32Config.fir@170054.8]
  wire [31:0] _T_89; // @[Parameters.scala 137:31:freechips.rocketchip.system.DefaultRV32Config.fir@170055.8]
  wire [32:0] _T_90; // @[Parameters.scala 137:49:freechips.rocketchip.system.DefaultRV32Config.fir@170056.8]
  wire [32:0] _T_92; // @[Parameters.scala 137:52:freechips.rocketchip.system.DefaultRV32Config.fir@170058.8]
  wire  _T_93; // @[Parameters.scala 137:67:freechips.rocketchip.system.DefaultRV32Config.fir@170059.8]
  wire [31:0] _T_94; // @[Parameters.scala 137:31:freechips.rocketchip.system.DefaultRV32Config.fir@170060.8]
  wire [32:0] _T_95; // @[Parameters.scala 137:49:freechips.rocketchip.system.DefaultRV32Config.fir@170061.8]
  wire [32:0] _T_97; // @[Parameters.scala 137:52:freechips.rocketchip.system.DefaultRV32Config.fir@170063.8]
  wire  _T_98; // @[Parameters.scala 137:67:freechips.rocketchip.system.DefaultRV32Config.fir@170064.8]
  wire  _T_99; // @[Parameters.scala 552:42:freechips.rocketchip.system.DefaultRV32Config.fir@170065.8]
  wire  _T_106; // @[Parameters.scala 93:42:freechips.rocketchip.system.DefaultRV32Config.fir@170072.8]
  wire [31:0] _T_109; // @[Parameters.scala 137:31:freechips.rocketchip.system.DefaultRV32Config.fir@170075.8]
  wire [32:0] _T_110; // @[Parameters.scala 137:49:freechips.rocketchip.system.DefaultRV32Config.fir@170076.8]
  wire [32:0] _T_112; // @[Parameters.scala 137:52:freechips.rocketchip.system.DefaultRV32Config.fir@170078.8]
  wire  _T_113; // @[Parameters.scala 137:67:freechips.rocketchip.system.DefaultRV32Config.fir@170079.8]
  wire  _T_114; // @[Parameters.scala 551:56:freechips.rocketchip.system.DefaultRV32Config.fir@170080.8]
  wire  _T_118; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@170084.8]
  wire  _T_119; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@170085.8]
  wire  _T_123; // @[Parameters.scala 92:48:freechips.rocketchip.system.DefaultRV32Config.fir@170096.8]
  wire  _T_124; // @[Mux.scala 27:72:freechips.rocketchip.system.DefaultRV32Config.fir@170097.8]
  wire  _T_129; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@170103.8]
  wire  _T_130; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@170104.8]
  wire  _T_132; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@170110.8]
  wire  _T_133; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@170111.8]
  wire  _T_136; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@170118.8]
  wire  _T_137; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@170119.8]
  wire  _T_139; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@170125.8]
  wire  _T_140; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@170126.8]
  wire  _T_141; // @[Bundles.scala 110:27:freechips.rocketchip.system.DefaultRV32Config.fir@170131.8]
  wire  _T_143; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@170133.8]
  wire  _T_144; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@170134.8]
  wire [3:0] _T_145; // @[Monitor.scala 86:18:freechips.rocketchip.system.DefaultRV32Config.fir@170139.8]
  wire  _T_146; // @[Monitor.scala 86:31:freechips.rocketchip.system.DefaultRV32Config.fir@170140.8]
  wire  _T_148; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@170142.8]
  wire  _T_149; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@170143.8]
  wire  _T_154; // @[Monitor.scala 90:25:freechips.rocketchip.system.DefaultRV32Config.fir@170157.6]
  wire  _T_232; // @[Monitor.scala 97:31:freechips.rocketchip.system.DefaultRV32Config.fir@170264.8]
  wire  _T_234; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@170266.8]
  wire  _T_235; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@170267.8]
  wire  _T_245; // @[Monitor.scala 102:25:freechips.rocketchip.system.DefaultRV32Config.fir@170290.6]
  wire  _T_247; // @[Parameters.scala 93:42:freechips.rocketchip.system.DefaultRV32Config.fir@170293.8]
  wire  _T_255; // @[Parameters.scala 551:56:freechips.rocketchip.system.DefaultRV32Config.fir@170301.8]
  wire  _T_290; // @[Parameters.scala 552:42:freechips.rocketchip.system.DefaultRV32Config.fir@170336.8]
  wire  _T_291; // @[Parameters.scala 552:42:freechips.rocketchip.system.DefaultRV32Config.fir@170337.8]
  wire  _T_292; // @[Parameters.scala 552:42:freechips.rocketchip.system.DefaultRV32Config.fir@170338.8]
  wire  _T_293; // @[Parameters.scala 552:42:freechips.rocketchip.system.DefaultRV32Config.fir@170339.8]
  wire  _T_294; // @[Parameters.scala 552:42:freechips.rocketchip.system.DefaultRV32Config.fir@170340.8]
  wire  _T_295; // @[Parameters.scala 551:56:freechips.rocketchip.system.DefaultRV32Config.fir@170341.8]
  wire  _T_297; // @[Parameters.scala 553:30:freechips.rocketchip.system.DefaultRV32Config.fir@170343.8]
  wire  _T_299; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@170345.8]
  wire  _T_300; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@170346.8]
  wire  _T_307; // @[Monitor.scala 106:31:freechips.rocketchip.system.DefaultRV32Config.fir@170365.8]
  wire  _T_309; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@170367.8]
  wire  _T_310; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@170368.8]
  wire  _T_311; // @[Monitor.scala 107:30:freechips.rocketchip.system.DefaultRV32Config.fir@170373.8]
  wire  _T_313; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@170375.8]
  wire  _T_314; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@170376.8]
  wire  _T_319; // @[Monitor.scala 111:25:freechips.rocketchip.system.DefaultRV32Config.fir@170390.6]
  wire  _T_354; // @[Parameters.scala 552:42:freechips.rocketchip.system.DefaultRV32Config.fir@170426.8]
  wire  _T_355; // @[Parameters.scala 552:42:freechips.rocketchip.system.DefaultRV32Config.fir@170427.8]
  wire  _T_356; // @[Parameters.scala 552:42:freechips.rocketchip.system.DefaultRV32Config.fir@170428.8]
  wire  _T_357; // @[Parameters.scala 551:56:freechips.rocketchip.system.DefaultRV32Config.fir@170429.8]
  wire  _T_366; // @[Parameters.scala 93:42:freechips.rocketchip.system.DefaultRV32Config.fir@170438.8]
  wire  _T_374; // @[Parameters.scala 551:56:freechips.rocketchip.system.DefaultRV32Config.fir@170446.8]
  wire  _T_376; // @[Parameters.scala 553:30:freechips.rocketchip.system.DefaultRV32Config.fir@170448.8]
  wire  _T_378; // @[Parameters.scala 553:30:freechips.rocketchip.system.DefaultRV32Config.fir@170450.8]
  wire  _T_380; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@170452.8]
  wire  _T_381; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@170453.8]
  wire  _T_396; // @[Monitor.scala 119:25:freechips.rocketchip.system.DefaultRV32Config.fir@170489.6]
  wire [3:0] _T_469; // @[Monitor.scala 124:33:freechips.rocketchip.system.DefaultRV32Config.fir@170579.8]
  wire [3:0] _T_470; // @[Monitor.scala 124:31:freechips.rocketchip.system.DefaultRV32Config.fir@170580.8]
  wire  _T_471; // @[Monitor.scala 124:40:freechips.rocketchip.system.DefaultRV32Config.fir@170581.8]
  wire  _T_473; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@170583.8]
  wire  _T_474; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@170584.8]
  wire  _T_475; // @[Monitor.scala 127:25:freechips.rocketchip.system.DefaultRV32Config.fir@170590.6]
  wire  _T_477; // @[Parameters.scala 93:42:freechips.rocketchip.system.DefaultRV32Config.fir@170593.8]
  wire  _T_501; // @[Parameters.scala 552:42:freechips.rocketchip.system.DefaultRV32Config.fir@170617.8]
  wire  _T_502; // @[Parameters.scala 552:42:freechips.rocketchip.system.DefaultRV32Config.fir@170618.8]
  wire  _T_503; // @[Parameters.scala 551:56:freechips.rocketchip.system.DefaultRV32Config.fir@170619.8]
  wire  _T_526; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@170642.8]
  wire  _T_527; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@170643.8]
  wire  _T_534; // @[Bundles.scala 140:33:freechips.rocketchip.system.DefaultRV32Config.fir@170662.8]
  wire  _T_536; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@170664.8]
  wire  _T_537; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@170665.8]
  wire  _T_542; // @[Monitor.scala 135:25:freechips.rocketchip.system.DefaultRV32Config.fir@170679.6]
  wire  _T_601; // @[Bundles.scala 147:30:freechips.rocketchip.system.DefaultRV32Config.fir@170751.8]
  wire  _T_603; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@170753.8]
  wire  _T_604; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@170754.8]
  wire  _T_609; // @[Monitor.scala 143:25:freechips.rocketchip.system.DefaultRV32Config.fir@170768.6]
  wire  _T_660; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@170820.8]
  wire  _T_661; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@170821.8]
  wire  _T_668; // @[Bundles.scala 160:28:freechips.rocketchip.system.DefaultRV32Config.fir@170840.8]
  wire  _T_670; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@170842.8]
  wire  _T_671; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@170843.8]
  wire  _T_680; // @[Bundles.scala 44:24:freechips.rocketchip.system.DefaultRV32Config.fir@170867.6]
  wire  _T_682; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@170869.6]
  wire  _T_683; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@170870.6]
  wire  _T_684; // @[Parameters.scala 47:9:freechips.rocketchip.system.DefaultRV32Config.fir@170875.6]
  wire  _T_687; // @[Parameters.scala 924:46:freechips.rocketchip.system.DefaultRV32Config.fir@170881.6]
  wire  _T_689; // @[Monitor.scala 307:25:freechips.rocketchip.system.DefaultRV32Config.fir@170883.6]
  wire  _T_691; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@170886.8]
  wire  _T_692; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@170887.8]
  wire  _T_693; // @[Monitor.scala 309:27:freechips.rocketchip.system.DefaultRV32Config.fir@170892.8]
  wire  _T_695; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@170894.8]
  wire  _T_696; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@170895.8]
  wire  _T_697; // @[Monitor.scala 310:28:freechips.rocketchip.system.DefaultRV32Config.fir@170900.8]
  wire  _T_699; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@170902.8]
  wire  _T_700; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@170903.8]
  wire  _T_701; // @[Monitor.scala 311:15:freechips.rocketchip.system.DefaultRV32Config.fir@170908.8]
  wire  _T_703; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@170910.8]
  wire  _T_704; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@170911.8]
  wire  _T_705; // @[Monitor.scala 312:15:freechips.rocketchip.system.DefaultRV32Config.fir@170916.8]
  wire  _T_707; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@170918.8]
  wire  _T_708; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@170919.8]
  wire  _T_709; // @[Monitor.scala 315:25:freechips.rocketchip.system.DefaultRV32Config.fir@170925.6]
  wire  _T_720; // @[Bundles.scala 104:26:freechips.rocketchip.system.DefaultRV32Config.fir@170949.8]
  wire  _T_722; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@170951.8]
  wire  _T_723; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@170952.8]
  wire  _T_724; // @[Monitor.scala 320:28:freechips.rocketchip.system.DefaultRV32Config.fir@170957.8]
  wire  _T_726; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@170959.8]
  wire  _T_727; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@170960.8]
  wire  _T_737; // @[Monitor.scala 325:25:freechips.rocketchip.system.DefaultRV32Config.fir@170983.6]
  wire  _T_757; // @[Monitor.scala 331:30:freechips.rocketchip.system.DefaultRV32Config.fir@171024.8]
  wire  _T_759; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@171026.8]
  wire  _T_760; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@171027.8]
  wire  _T_766; // @[Monitor.scala 335:25:freechips.rocketchip.system.DefaultRV32Config.fir@171042.6]
  wire  _T_783; // @[Monitor.scala 343:25:freechips.rocketchip.system.DefaultRV32Config.fir@171077.6]
  wire  _T_801; // @[Monitor.scala 351:25:freechips.rocketchip.system.DefaultRV32Config.fir@171113.6]
  wire  _T_818; // @[Bundles.scala 42:24:freechips.rocketchip.system.DefaultRV32Config.fir@171150.6]
  wire  _T_820; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@171152.6]
  wire  _T_821; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@171153.6]
  wire  _T_822; // @[Parameters.scala 47:9:freechips.rocketchip.system.DefaultRV32Config.fir@171158.6]
  wire [32:0] _T_825; // @[Parameters.scala 137:49:freechips.rocketchip.system.DefaultRV32Config.fir@171161.6]
  wire [31:0] _T_842; // @[Parameters.scala 137:31:freechips.rocketchip.system.DefaultRV32Config.fir@171182.6]
  wire [32:0] _T_843; // @[Parameters.scala 137:49:freechips.rocketchip.system.DefaultRV32Config.fir@171183.6]
  wire [32:0] _T_845; // @[Parameters.scala 137:52:freechips.rocketchip.system.DefaultRV32Config.fir@171185.6]
  wire  _T_846; // @[Parameters.scala 137:67:freechips.rocketchip.system.DefaultRV32Config.fir@171186.6]
  wire [31:0] _T_847; // @[Parameters.scala 137:31:freechips.rocketchip.system.DefaultRV32Config.fir@171187.6]
  wire [32:0] _T_848; // @[Parameters.scala 137:49:freechips.rocketchip.system.DefaultRV32Config.fir@171188.6]
  wire [32:0] _T_850; // @[Parameters.scala 137:52:freechips.rocketchip.system.DefaultRV32Config.fir@171190.6]
  wire  _T_851; // @[Parameters.scala 137:67:freechips.rocketchip.system.DefaultRV32Config.fir@171191.6]
  wire [31:0] _T_852; // @[Parameters.scala 137:31:freechips.rocketchip.system.DefaultRV32Config.fir@171192.6]
  wire [32:0] _T_853; // @[Parameters.scala 137:49:freechips.rocketchip.system.DefaultRV32Config.fir@171193.6]
  wire [32:0] _T_855; // @[Parameters.scala 137:52:freechips.rocketchip.system.DefaultRV32Config.fir@171195.6]
  wire  _T_856; // @[Parameters.scala 137:67:freechips.rocketchip.system.DefaultRV32Config.fir@171196.6]
  wire [32:0] _T_860; // @[Parameters.scala 137:52:freechips.rocketchip.system.DefaultRV32Config.fir@171200.6]
  wire  _T_861; // @[Parameters.scala 137:67:freechips.rocketchip.system.DefaultRV32Config.fir@171201.6]
  wire [31:0] _T_862; // @[Parameters.scala 137:31:freechips.rocketchip.system.DefaultRV32Config.fir@171202.6]
  wire [32:0] _T_863; // @[Parameters.scala 137:49:freechips.rocketchip.system.DefaultRV32Config.fir@171203.6]
  wire [32:0] _T_865; // @[Parameters.scala 137:52:freechips.rocketchip.system.DefaultRV32Config.fir@171205.6]
  wire  _T_866; // @[Parameters.scala 137:67:freechips.rocketchip.system.DefaultRV32Config.fir@171206.6]
  wire [31:0] _T_867; // @[Parameters.scala 137:31:freechips.rocketchip.system.DefaultRV32Config.fir@171207.6]
  wire [32:0] _T_868; // @[Parameters.scala 137:49:freechips.rocketchip.system.DefaultRV32Config.fir@171208.6]
  wire [32:0] _T_870; // @[Parameters.scala 137:52:freechips.rocketchip.system.DefaultRV32Config.fir@171210.6]
  wire  _T_871; // @[Parameters.scala 137:67:freechips.rocketchip.system.DefaultRV32Config.fir@171211.6]
  wire [31:0] _T_872; // @[Parameters.scala 137:31:freechips.rocketchip.system.DefaultRV32Config.fir@171212.6]
  wire [32:0] _T_873; // @[Parameters.scala 137:49:freechips.rocketchip.system.DefaultRV32Config.fir@171213.6]
  wire [32:0] _T_875; // @[Parameters.scala 137:52:freechips.rocketchip.system.DefaultRV32Config.fir@171215.6]
  wire  _T_876; // @[Parameters.scala 137:67:freechips.rocketchip.system.DefaultRV32Config.fir@171216.6]
  wire  _T_878; // @[Parameters.scala 535:64:freechips.rocketchip.system.DefaultRV32Config.fir@171226.6]
  wire  _T_879; // @[Parameters.scala 535:64:freechips.rocketchip.system.DefaultRV32Config.fir@171227.6]
  wire  _T_880; // @[Parameters.scala 535:64:freechips.rocketchip.system.DefaultRV32Config.fir@171228.6]
  wire  _T_881; // @[Parameters.scala 535:64:freechips.rocketchip.system.DefaultRV32Config.fir@171229.6]
  wire  _T_882; // @[Parameters.scala 535:64:freechips.rocketchip.system.DefaultRV32Config.fir@171230.6]
  wire  _T_883; // @[Parameters.scala 535:64:freechips.rocketchip.system.DefaultRV32Config.fir@171231.6]
  wire [26:0] _T_885; // @[package.scala 207:77:freechips.rocketchip.system.DefaultRV32Config.fir@171233.6]
  wire [11:0] _T_887; // @[package.scala 207:46:freechips.rocketchip.system.DefaultRV32Config.fir@171235.6]
  wire [31:0] _GEN_72; // @[Edges.scala 22:16:freechips.rocketchip.system.DefaultRV32Config.fir@171236.6]
  wire [31:0] _T_888; // @[Edges.scala 22:16:freechips.rocketchip.system.DefaultRV32Config.fir@171236.6]
  wire  _T_889; // @[Edges.scala 22:24:freechips.rocketchip.system.DefaultRV32Config.fir@171237.6]
  wire [1:0] _T_892; // @[OneHot.scala 65:12:freechips.rocketchip.system.DefaultRV32Config.fir@171240.6]
  wire [1:0] _T_894; // @[Misc.scala 201:81:freechips.rocketchip.system.DefaultRV32Config.fir@171242.6]
  wire  _T_895; // @[Misc.scala 205:21:freechips.rocketchip.system.DefaultRV32Config.fir@171243.6]
  wire  _T_898; // @[Misc.scala 210:20:freechips.rocketchip.system.DefaultRV32Config.fir@171246.6]
  wire  _T_900; // @[Misc.scala 214:38:freechips.rocketchip.system.DefaultRV32Config.fir@171248.6]
  wire  _T_901; // @[Misc.scala 214:29:freechips.rocketchip.system.DefaultRV32Config.fir@171249.6]
  wire  _T_903; // @[Misc.scala 214:38:freechips.rocketchip.system.DefaultRV32Config.fir@171251.6]
  wire  _T_904; // @[Misc.scala 214:29:freechips.rocketchip.system.DefaultRV32Config.fir@171252.6]
  wire  _T_907; // @[Misc.scala 210:20:freechips.rocketchip.system.DefaultRV32Config.fir@171255.6]
  wire  _T_908; // @[Misc.scala 213:27:freechips.rocketchip.system.DefaultRV32Config.fir@171256.6]
  wire  _T_909; // @[Misc.scala 214:38:freechips.rocketchip.system.DefaultRV32Config.fir@171257.6]
  wire  _T_910; // @[Misc.scala 214:29:freechips.rocketchip.system.DefaultRV32Config.fir@171258.6]
  wire  _T_911; // @[Misc.scala 213:27:freechips.rocketchip.system.DefaultRV32Config.fir@171259.6]
  wire  _T_912; // @[Misc.scala 214:38:freechips.rocketchip.system.DefaultRV32Config.fir@171260.6]
  wire  _T_913; // @[Misc.scala 214:29:freechips.rocketchip.system.DefaultRV32Config.fir@171261.6]
  wire  _T_914; // @[Misc.scala 213:27:freechips.rocketchip.system.DefaultRV32Config.fir@171262.6]
  wire  _T_915; // @[Misc.scala 214:38:freechips.rocketchip.system.DefaultRV32Config.fir@171263.6]
  wire  _T_916; // @[Misc.scala 214:29:freechips.rocketchip.system.DefaultRV32Config.fir@171264.6]
  wire  _T_917; // @[Misc.scala 213:27:freechips.rocketchip.system.DefaultRV32Config.fir@171265.6]
  wire  _T_918; // @[Misc.scala 214:38:freechips.rocketchip.system.DefaultRV32Config.fir@171266.6]
  wire  _T_919; // @[Misc.scala 214:29:freechips.rocketchip.system.DefaultRV32Config.fir@171267.6]
  wire [3:0] _T_922; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@171270.6]
  wire  _T_931; // @[Monitor.scala 164:25:freechips.rocketchip.system.DefaultRV32Config.fir@171283.6]
  wire  _T_935; // @[Parameters.scala 92:48:freechips.rocketchip.system.DefaultRV32Config.fir@171291.8]
  wire  _T_936; // @[Mux.scala 27:72:freechips.rocketchip.system.DefaultRV32Config.fir@171292.8]
  wire  _T_941; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@171298.8]
  wire  _T_942; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@171299.8]
  wire  _T_944; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@171305.8]
  wire  _T_945; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@171306.8]
  wire  _T_950; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@171319.8]
  wire  _T_951; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@171320.8]
  wire  _T_952; // @[Bundles.scala 104:26:freechips.rocketchip.system.DefaultRV32Config.fir@171325.8]
  wire  _T_954; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@171327.8]
  wire  _T_955; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@171328.8]
  wire  _T_956; // @[Monitor.scala 170:30:freechips.rocketchip.system.DefaultRV32Config.fir@171333.8]
  wire  _T_958; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@171335.8]
  wire  _T_959; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@171336.8]
  wire  _T_960; // @[Monitor.scala 171:18:freechips.rocketchip.system.DefaultRV32Config.fir@171341.8]
  wire  _T_962; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@171343.8]
  wire  _T_963; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@171344.8]
  wire  _T_964; // @[Monitor.scala 174:25:freechips.rocketchip.system.DefaultRV32Config.fir@171350.6]
  wire  _T_967; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@171354.8]
  wire  _T_977; // @[Monitor.scala 179:31:freechips.rocketchip.system.DefaultRV32Config.fir@171380.8]
  wire  _T_979; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@171382.8]
  wire  _T_980; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@171383.8]
  wire  _T_989; // @[Monitor.scala 184:25:freechips.rocketchip.system.DefaultRV32Config.fir@171405.6]
  wire  _T_1010; // @[Monitor.scala 193:25:freechips.rocketchip.system.DefaultRV32Config.fir@171452.6]
  wire [3:0] _T_1027; // @[Monitor.scala 199:33:freechips.rocketchip.system.DefaultRV32Config.fir@171490.8]
  wire [3:0] _T_1028; // @[Monitor.scala 199:31:freechips.rocketchip.system.DefaultRV32Config.fir@171491.8]
  wire  _T_1029; // @[Monitor.scala 199:40:freechips.rocketchip.system.DefaultRV32Config.fir@171492.8]
  wire  _T_1031; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@171494.8]
  wire  _T_1032; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@171495.8]
  wire  _T_1033; // @[Monitor.scala 202:25:freechips.rocketchip.system.DefaultRV32Config.fir@171501.6]
  wire  _T_1054; // @[Monitor.scala 211:25:freechips.rocketchip.system.DefaultRV32Config.fir@171548.6]
  wire  _T_1075; // @[Monitor.scala 220:25:freechips.rocketchip.system.DefaultRV32Config.fir@171595.6]
  wire  _T_1100; // @[Parameters.scala 47:9:freechips.rocketchip.system.DefaultRV32Config.fir@171652.6]
  wire  _T_1103; // @[Parameters.scala 924:46:freechips.rocketchip.system.DefaultRV32Config.fir@171658.6]
  wire [26:0] _T_1105; // @[package.scala 207:77:freechips.rocketchip.system.DefaultRV32Config.fir@171660.6]
  wire [11:0] _T_1107; // @[package.scala 207:46:freechips.rocketchip.system.DefaultRV32Config.fir@171662.6]
  wire [31:0] _GEN_73; // @[Edges.scala 22:16:freechips.rocketchip.system.DefaultRV32Config.fir@171663.6]
  wire [31:0] _T_1108; // @[Edges.scala 22:16:freechips.rocketchip.system.DefaultRV32Config.fir@171663.6]
  wire  _T_1109; // @[Edges.scala 22:24:freechips.rocketchip.system.DefaultRV32Config.fir@171664.6]
  wire [31:0] _T_1110; // @[Parameters.scala 137:31:freechips.rocketchip.system.DefaultRV32Config.fir@171665.6]
  wire [32:0] _T_1111; // @[Parameters.scala 137:49:freechips.rocketchip.system.DefaultRV32Config.fir@171666.6]
  wire [32:0] _T_1113; // @[Parameters.scala 137:52:freechips.rocketchip.system.DefaultRV32Config.fir@171668.6]
  wire  _T_1114; // @[Parameters.scala 137:67:freechips.rocketchip.system.DefaultRV32Config.fir@171669.6]
  wire [31:0] _T_1115; // @[Parameters.scala 137:31:freechips.rocketchip.system.DefaultRV32Config.fir@171670.6]
  wire [32:0] _T_1116; // @[Parameters.scala 137:49:freechips.rocketchip.system.DefaultRV32Config.fir@171671.6]
  wire [32:0] _T_1118; // @[Parameters.scala 137:52:freechips.rocketchip.system.DefaultRV32Config.fir@171673.6]
  wire  _T_1119; // @[Parameters.scala 137:67:freechips.rocketchip.system.DefaultRV32Config.fir@171674.6]
  wire [31:0] _T_1120; // @[Parameters.scala 137:31:freechips.rocketchip.system.DefaultRV32Config.fir@171675.6]
  wire [32:0] _T_1121; // @[Parameters.scala 137:49:freechips.rocketchip.system.DefaultRV32Config.fir@171676.6]
  wire [32:0] _T_1123; // @[Parameters.scala 137:52:freechips.rocketchip.system.DefaultRV32Config.fir@171678.6]
  wire  _T_1124; // @[Parameters.scala 137:67:freechips.rocketchip.system.DefaultRV32Config.fir@171679.6]
  wire [32:0] _T_1126; // @[Parameters.scala 137:49:freechips.rocketchip.system.DefaultRV32Config.fir@171681.6]
  wire [32:0] _T_1128; // @[Parameters.scala 137:52:freechips.rocketchip.system.DefaultRV32Config.fir@171683.6]
  wire  _T_1129; // @[Parameters.scala 137:67:freechips.rocketchip.system.DefaultRV32Config.fir@171684.6]
  wire [31:0] _T_1130; // @[Parameters.scala 137:31:freechips.rocketchip.system.DefaultRV32Config.fir@171685.6]
  wire [32:0] _T_1131; // @[Parameters.scala 137:49:freechips.rocketchip.system.DefaultRV32Config.fir@171686.6]
  wire [32:0] _T_1133; // @[Parameters.scala 137:52:freechips.rocketchip.system.DefaultRV32Config.fir@171688.6]
  wire  _T_1134; // @[Parameters.scala 137:67:freechips.rocketchip.system.DefaultRV32Config.fir@171689.6]
  wire [31:0] _T_1135; // @[Parameters.scala 137:31:freechips.rocketchip.system.DefaultRV32Config.fir@171690.6]
  wire [32:0] _T_1136; // @[Parameters.scala 137:49:freechips.rocketchip.system.DefaultRV32Config.fir@171691.6]
  wire [32:0] _T_1138; // @[Parameters.scala 137:52:freechips.rocketchip.system.DefaultRV32Config.fir@171693.6]
  wire  _T_1139; // @[Parameters.scala 137:67:freechips.rocketchip.system.DefaultRV32Config.fir@171694.6]
  wire [31:0] _T_1140; // @[Parameters.scala 137:31:freechips.rocketchip.system.DefaultRV32Config.fir@171695.6]
  wire [32:0] _T_1141; // @[Parameters.scala 137:49:freechips.rocketchip.system.DefaultRV32Config.fir@171696.6]
  wire [32:0] _T_1143; // @[Parameters.scala 137:52:freechips.rocketchip.system.DefaultRV32Config.fir@171698.6]
  wire  _T_1144; // @[Parameters.scala 137:67:freechips.rocketchip.system.DefaultRV32Config.fir@171699.6]
  wire  _T_1146; // @[Parameters.scala 535:64:freechips.rocketchip.system.DefaultRV32Config.fir@171709.6]
  wire  _T_1147; // @[Parameters.scala 535:64:freechips.rocketchip.system.DefaultRV32Config.fir@171710.6]
  wire  _T_1148; // @[Parameters.scala 535:64:freechips.rocketchip.system.DefaultRV32Config.fir@171711.6]
  wire  _T_1149; // @[Parameters.scala 535:64:freechips.rocketchip.system.DefaultRV32Config.fir@171712.6]
  wire  _T_1150; // @[Parameters.scala 535:64:freechips.rocketchip.system.DefaultRV32Config.fir@171713.6]
  wire  _T_1151; // @[Parameters.scala 535:64:freechips.rocketchip.system.DefaultRV32Config.fir@171714.6]
  wire  _T_1172; // @[Monitor.scala 239:25:freechips.rocketchip.system.DefaultRV32Config.fir@171739.6]
  wire  _T_1174; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@171742.8]
  wire  _T_1175; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@171743.8]
  wire  _T_1177; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@171749.8]
  wire  _T_1178; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@171750.8]
  wire  _T_1179; // @[Monitor.scala 242:30:freechips.rocketchip.system.DefaultRV32Config.fir@171755.8]
  wire  _T_1181; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@171757.8]
  wire  _T_1182; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@171758.8]
  wire  _T_1184; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@171764.8]
  wire  _T_1185; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@171765.8]
  wire  _T_1186; // @[Bundles.scala 122:29:freechips.rocketchip.system.DefaultRV32Config.fir@171770.8]
  wire  _T_1188; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@171772.8]
  wire  _T_1189; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@171773.8]
  wire  _T_1194; // @[Monitor.scala 248:25:freechips.rocketchip.system.DefaultRV32Config.fir@171787.6]
  wire  _T_1212; // @[Monitor.scala 256:25:freechips.rocketchip.system.DefaultRV32Config.fir@171827.6]
  wire  _T_1251; // @[Parameters.scala 93:42:freechips.rocketchip.system.DefaultRV32Config.fir@171867.8]
  wire  _T_1259; // @[Parameters.scala 551:56:freechips.rocketchip.system.DefaultRV32Config.fir@171875.8]
  wire  _T_1263; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@171879.8]
  wire  _T_1264; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@171880.8]
  wire  _T_1268; // @[Parameters.scala 92:48:freechips.rocketchip.system.DefaultRV32Config.fir@171891.8]
  wire  _T_1269; // @[Mux.scala 27:72:freechips.rocketchip.system.DefaultRV32Config.fir@171892.8]
  wire  _T_1274; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@171898.8]
  wire  _T_1275; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@171899.8]
  wire  _T_1286; // @[Bundles.scala 116:29:freechips.rocketchip.system.DefaultRV32Config.fir@171926.8]
  wire  _T_1288; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@171928.8]
  wire  _T_1289; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@171929.8]
  wire  _T_1294; // @[Monitor.scala 266:25:freechips.rocketchip.system.DefaultRV32Config.fir@171943.6]
  wire  _T_1372; // @[Monitor.scala 275:25:freechips.rocketchip.system.DefaultRV32Config.fir@172051.6]
  wire  _T_1382; // @[Monitor.scala 279:31:freechips.rocketchip.system.DefaultRV32Config.fir@172074.8]
  wire  _T_1384; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@172076.8]
  wire  _T_1385; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@172077.8]
  wire  _T_1390; // @[Monitor.scala 283:25:freechips.rocketchip.system.DefaultRV32Config.fir@172091.6]
  wire  _T_1404; // @[Monitor.scala 290:25:freechips.rocketchip.system.DefaultRV32Config.fir@172123.6]
  wire  _T_1426; // @[Decoupled.scala 40:37:freechips.rocketchip.system.DefaultRV32Config.fir@172174.4]
  wire  _T_1433; // @[Edges.scala 93:28:freechips.rocketchip.system.DefaultRV32Config.fir@172181.4]
  reg [9:0] _T_1435; // @[Edges.scala 230:27:freechips.rocketchip.system.DefaultRV32Config.fir@172183.4]
  wire [9:0] _T_1437; // @[Edges.scala 231:28:freechips.rocketchip.system.DefaultRV32Config.fir@172185.4]
  wire  _T_1438; // @[Edges.scala 232:25:freechips.rocketchip.system.DefaultRV32Config.fir@172186.4]
  reg [2:0] _T_1446; // @[Monitor.scala 381:22:freechips.rocketchip.system.DefaultRV32Config.fir@172197.4]
  reg [2:0] _T_1447; // @[Monitor.scala 382:22:freechips.rocketchip.system.DefaultRV32Config.fir@172198.4]
  reg [3:0] _T_1448; // @[Monitor.scala 383:22:freechips.rocketchip.system.DefaultRV32Config.fir@172199.4]
  reg  _T_1449; // @[Monitor.scala 384:22:freechips.rocketchip.system.DefaultRV32Config.fir@172200.4]
  reg [31:0] _T_1450; // @[Monitor.scala 385:22:freechips.rocketchip.system.DefaultRV32Config.fir@172201.4]
  wire  _T_1451; // @[Monitor.scala 386:22:freechips.rocketchip.system.DefaultRV32Config.fir@172202.4]
  wire  _T_1452; // @[Monitor.scala 386:19:freechips.rocketchip.system.DefaultRV32Config.fir@172203.4]
  wire  _T_1453; // @[Monitor.scala 387:32:freechips.rocketchip.system.DefaultRV32Config.fir@172205.6]
  wire  _T_1455; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@172207.6]
  wire  _T_1456; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@172208.6]
  wire  _T_1457; // @[Monitor.scala 388:32:freechips.rocketchip.system.DefaultRV32Config.fir@172213.6]
  wire  _T_1459; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@172215.6]
  wire  _T_1460; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@172216.6]
  wire  _T_1461; // @[Monitor.scala 389:32:freechips.rocketchip.system.DefaultRV32Config.fir@172221.6]
  wire  _T_1463; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@172223.6]
  wire  _T_1464; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@172224.6]
  wire  _T_1465; // @[Monitor.scala 390:32:freechips.rocketchip.system.DefaultRV32Config.fir@172229.6]
  wire  _T_1467; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@172231.6]
  wire  _T_1468; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@172232.6]
  wire  _T_1469; // @[Monitor.scala 391:32:freechips.rocketchip.system.DefaultRV32Config.fir@172237.6]
  wire  _T_1471; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@172239.6]
  wire  _T_1472; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@172240.6]
  wire  _T_1474; // @[Monitor.scala 393:20:freechips.rocketchip.system.DefaultRV32Config.fir@172247.4]
  wire  _T_1475; // @[Decoupled.scala 40:37:freechips.rocketchip.system.DefaultRV32Config.fir@172255.4]
  wire [26:0] _T_1477; // @[package.scala 207:77:freechips.rocketchip.system.DefaultRV32Config.fir@172257.4]
  wire [11:0] _T_1479; // @[package.scala 207:46:freechips.rocketchip.system.DefaultRV32Config.fir@172259.4]
  reg [9:0] _T_1483; // @[Edges.scala 230:27:freechips.rocketchip.system.DefaultRV32Config.fir@172263.4]
  wire [9:0] _T_1485; // @[Edges.scala 231:28:freechips.rocketchip.system.DefaultRV32Config.fir@172265.4]
  wire  _T_1486; // @[Edges.scala 232:25:freechips.rocketchip.system.DefaultRV32Config.fir@172266.4]
  reg [2:0] _T_1494; // @[Monitor.scala 532:22:freechips.rocketchip.system.DefaultRV32Config.fir@172277.4]
  reg [1:0] _T_1495; // @[Monitor.scala 533:22:freechips.rocketchip.system.DefaultRV32Config.fir@172278.4]
  reg [3:0] _T_1496; // @[Monitor.scala 534:22:freechips.rocketchip.system.DefaultRV32Config.fir@172279.4]
  reg  _T_1497; // @[Monitor.scala 535:22:freechips.rocketchip.system.DefaultRV32Config.fir@172280.4]
  reg [1:0] _T_1498; // @[Monitor.scala 536:22:freechips.rocketchip.system.DefaultRV32Config.fir@172281.4]
  reg  _T_1499; // @[Monitor.scala 537:22:freechips.rocketchip.system.DefaultRV32Config.fir@172282.4]
  wire  _T_1500; // @[Monitor.scala 538:22:freechips.rocketchip.system.DefaultRV32Config.fir@172283.4]
  wire  _T_1501; // @[Monitor.scala 538:19:freechips.rocketchip.system.DefaultRV32Config.fir@172284.4]
  wire  _T_1502; // @[Monitor.scala 539:29:freechips.rocketchip.system.DefaultRV32Config.fir@172286.6]
  wire  _T_1504; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@172288.6]
  wire  _T_1505; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@172289.6]
  wire  _T_1506; // @[Monitor.scala 540:29:freechips.rocketchip.system.DefaultRV32Config.fir@172294.6]
  wire  _T_1508; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@172296.6]
  wire  _T_1509; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@172297.6]
  wire  _T_1510; // @[Monitor.scala 541:29:freechips.rocketchip.system.DefaultRV32Config.fir@172302.6]
  wire  _T_1512; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@172304.6]
  wire  _T_1513; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@172305.6]
  wire  _T_1514; // @[Monitor.scala 542:29:freechips.rocketchip.system.DefaultRV32Config.fir@172310.6]
  wire  _T_1516; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@172312.6]
  wire  _T_1517; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@172313.6]
  wire  _T_1518; // @[Monitor.scala 543:29:freechips.rocketchip.system.DefaultRV32Config.fir@172318.6]
  wire  _T_1520; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@172320.6]
  wire  _T_1521; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@172321.6]
  wire  _T_1522; // @[Monitor.scala 544:29:freechips.rocketchip.system.DefaultRV32Config.fir@172326.6]
  wire  _T_1524; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@172328.6]
  wire  _T_1525; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@172329.6]
  wire  _T_1527; // @[Monitor.scala 546:20:freechips.rocketchip.system.DefaultRV32Config.fir@172336.4]
  wire  _T_1528; // @[Decoupled.scala 40:37:freechips.rocketchip.system.DefaultRV32Config.fir@172345.4]
  reg [9:0] _T_1537; // @[Edges.scala 230:27:freechips.rocketchip.system.DefaultRV32Config.fir@172354.4]
  wire [9:0] _T_1539; // @[Edges.scala 231:28:freechips.rocketchip.system.DefaultRV32Config.fir@172356.4]
  wire  _T_1540; // @[Edges.scala 232:25:freechips.rocketchip.system.DefaultRV32Config.fir@172357.4]
  reg [2:0] _T_1548; // @[Monitor.scala 404:22:freechips.rocketchip.system.DefaultRV32Config.fir@172368.4]
  reg [1:0] _T_1549; // @[Monitor.scala 405:22:freechips.rocketchip.system.DefaultRV32Config.fir@172369.4]
  reg [3:0] _T_1550; // @[Monitor.scala 406:22:freechips.rocketchip.system.DefaultRV32Config.fir@172370.4]
  reg  _T_1551; // @[Monitor.scala 407:22:freechips.rocketchip.system.DefaultRV32Config.fir@172371.4]
  reg [31:0] _T_1552; // @[Monitor.scala 408:22:freechips.rocketchip.system.DefaultRV32Config.fir@172372.4]
  wire  _T_1553; // @[Monitor.scala 409:22:freechips.rocketchip.system.DefaultRV32Config.fir@172373.4]
  wire  _T_1554; // @[Monitor.scala 409:19:freechips.rocketchip.system.DefaultRV32Config.fir@172374.4]
  wire  _T_1555; // @[Monitor.scala 410:32:freechips.rocketchip.system.DefaultRV32Config.fir@172376.6]
  wire  _T_1557; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@172378.6]
  wire  _T_1558; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@172379.6]
  wire  _T_1559; // @[Monitor.scala 411:32:freechips.rocketchip.system.DefaultRV32Config.fir@172384.6]
  wire  _T_1561; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@172386.6]
  wire  _T_1562; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@172387.6]
  wire  _T_1563; // @[Monitor.scala 412:32:freechips.rocketchip.system.DefaultRV32Config.fir@172392.6]
  wire  _T_1565; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@172394.6]
  wire  _T_1566; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@172395.6]
  wire  _T_1567; // @[Monitor.scala 413:32:freechips.rocketchip.system.DefaultRV32Config.fir@172400.6]
  wire  _T_1569; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@172402.6]
  wire  _T_1570; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@172403.6]
  wire  _T_1571; // @[Monitor.scala 414:32:freechips.rocketchip.system.DefaultRV32Config.fir@172408.6]
  wire  _T_1573; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@172410.6]
  wire  _T_1574; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@172411.6]
  wire  _T_1576; // @[Monitor.scala 416:20:freechips.rocketchip.system.DefaultRV32Config.fir@172418.4]
  wire  _T_1577; // @[Decoupled.scala 40:37:freechips.rocketchip.system.DefaultRV32Config.fir@172426.4]
  reg [9:0] _T_1585; // @[Edges.scala 230:27:freechips.rocketchip.system.DefaultRV32Config.fir@172434.4]
  wire [9:0] _T_1587; // @[Edges.scala 231:28:freechips.rocketchip.system.DefaultRV32Config.fir@172436.4]
  wire  _T_1588; // @[Edges.scala 232:25:freechips.rocketchip.system.DefaultRV32Config.fir@172437.4]
  reg [2:0] _T_1596; // @[Monitor.scala 509:22:freechips.rocketchip.system.DefaultRV32Config.fir@172448.4]
  reg [2:0] _T_1597; // @[Monitor.scala 510:22:freechips.rocketchip.system.DefaultRV32Config.fir@172449.4]
  reg [3:0] _T_1598; // @[Monitor.scala 511:22:freechips.rocketchip.system.DefaultRV32Config.fir@172450.4]
  reg  _T_1599; // @[Monitor.scala 512:22:freechips.rocketchip.system.DefaultRV32Config.fir@172451.4]
  reg [31:0] _T_1600; // @[Monitor.scala 513:22:freechips.rocketchip.system.DefaultRV32Config.fir@172452.4]
  wire  _T_1601; // @[Monitor.scala 514:22:freechips.rocketchip.system.DefaultRV32Config.fir@172453.4]
  wire  _T_1602; // @[Monitor.scala 514:19:freechips.rocketchip.system.DefaultRV32Config.fir@172454.4]
  wire  _T_1603; // @[Monitor.scala 515:32:freechips.rocketchip.system.DefaultRV32Config.fir@172456.6]
  wire  _T_1605; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@172458.6]
  wire  _T_1606; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@172459.6]
  wire  _T_1607; // @[Monitor.scala 516:32:freechips.rocketchip.system.DefaultRV32Config.fir@172464.6]
  wire  _T_1609; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@172466.6]
  wire  _T_1610; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@172467.6]
  wire  _T_1611; // @[Monitor.scala 517:32:freechips.rocketchip.system.DefaultRV32Config.fir@172472.6]
  wire  _T_1613; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@172474.6]
  wire  _T_1614; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@172475.6]
  wire  _T_1615; // @[Monitor.scala 518:32:freechips.rocketchip.system.DefaultRV32Config.fir@172480.6]
  wire  _T_1617; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@172482.6]
  wire  _T_1618; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@172483.6]
  wire  _T_1619; // @[Monitor.scala 519:32:freechips.rocketchip.system.DefaultRV32Config.fir@172488.6]
  wire  _T_1621; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@172490.6]
  wire  _T_1622; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@172491.6]
  wire  _T_1624; // @[Monitor.scala 521:20:freechips.rocketchip.system.DefaultRV32Config.fir@172498.4]
  reg [1:0] inflight; // @[Monitor.scala 608:27:freechips.rocketchip.system.DefaultRV32Config.fir@172506.4]
  reg [7:0] inflight_opcodes; // @[Monitor.scala 610:35:freechips.rocketchip.system.DefaultRV32Config.fir@172507.4]
  reg [15:0] inflight_sizes; // @[Monitor.scala 612:33:freechips.rocketchip.system.DefaultRV32Config.fir@172508.4]
  reg [9:0] _T_1634; // @[Edges.scala 230:27:freechips.rocketchip.system.DefaultRV32Config.fir@172518.4]
  wire [9:0] _T_1636; // @[Edges.scala 231:28:freechips.rocketchip.system.DefaultRV32Config.fir@172520.4]
  wire  a_first; // @[Edges.scala 232:25:freechips.rocketchip.system.DefaultRV32Config.fir@172521.4]
  reg [9:0] _T_1652; // @[Edges.scala 230:27:freechips.rocketchip.system.DefaultRV32Config.fir@172540.4]
  wire [9:0] _T_1654; // @[Edges.scala 231:28:freechips.rocketchip.system.DefaultRV32Config.fir@172542.4]
  wire  d_first; // @[Edges.scala 232:25:freechips.rocketchip.system.DefaultRV32Config.fir@172543.4]
  wire [2:0] _GEN_74; // @[Monitor.scala 629:69:freechips.rocketchip.system.DefaultRV32Config.fir@172562.4]
  wire [3:0] _T_1662; // @[Monitor.scala 629:69:freechips.rocketchip.system.DefaultRV32Config.fir@172562.4]
  wire [7:0] _T_1663; // @[Monitor.scala 629:44:freechips.rocketchip.system.DefaultRV32Config.fir@172563.4]
  wire [15:0] _T_1667; // @[Monitor.scala 606:57:freechips.rocketchip.system.DefaultRV32Config.fir@172567.4]
  wire [15:0] _GEN_75; // @[Monitor.scala 629:97:freechips.rocketchip.system.DefaultRV32Config.fir@172568.4]
  wire [15:0] _T_1668; // @[Monitor.scala 629:97:freechips.rocketchip.system.DefaultRV32Config.fir@172568.4]
  wire [15:0] _T_1669; // @[Monitor.scala 629:152:freechips.rocketchip.system.DefaultRV32Config.fir@172569.4]
  wire [3:0] _T_1670; // @[Monitor.scala 633:65:freechips.rocketchip.system.DefaultRV32Config.fir@172573.4]
  wire [15:0] _T_1671; // @[Monitor.scala 633:40:freechips.rocketchip.system.DefaultRV32Config.fir@172574.4]
  wire [15:0] _T_1675; // @[Monitor.scala 606:57:freechips.rocketchip.system.DefaultRV32Config.fir@172578.4]
  wire [15:0] _T_1676; // @[Monitor.scala 633:91:freechips.rocketchip.system.DefaultRV32Config.fir@172579.4]
  wire [15:0] _T_1677; // @[Monitor.scala 633:144:freechips.rocketchip.system.DefaultRV32Config.fir@172580.4]
  wire  _T_1681; // @[Monitor.scala 643:27:freechips.rocketchip.system.DefaultRV32Config.fir@172605.4]
  wire [1:0] _T_1683; // @[OneHot.scala 58:35:freechips.rocketchip.system.DefaultRV32Config.fir@172608.6]
  wire [3:0] _T_1684; // @[Monitor.scala 645:53:freechips.rocketchip.system.DefaultRV32Config.fir@172610.6]
  wire [3:0] _T_1685; // @[Monitor.scala 645:61:freechips.rocketchip.system.DefaultRV32Config.fir@172611.6]
  wire [4:0] _T_1686; // @[Monitor.scala 646:49:freechips.rocketchip.system.DefaultRV32Config.fir@172613.6]
  wire [4:0] _T_1687; // @[Monitor.scala 646:57:freechips.rocketchip.system.DefaultRV32Config.fir@172614.6]
  wire [2:0] _GEN_78; // @[Monitor.scala 647:72:freechips.rocketchip.system.DefaultRV32Config.fir@172616.6]
  wire [3:0] _T_1688; // @[Monitor.scala 647:72:freechips.rocketchip.system.DefaultRV32Config.fir@172616.6]
  wire [3:0] a_opcodes_set_interm; // @[Monitor.scala 643:72:freechips.rocketchip.system.DefaultRV32Config.fir@172607.4]
  wire [18:0] _GEN_79; // @[Monitor.scala 647:47:freechips.rocketchip.system.DefaultRV32Config.fir@172617.6]
  wire [18:0] _T_1689; // @[Monitor.scala 647:47:freechips.rocketchip.system.DefaultRV32Config.fir@172617.6]
  wire [3:0] _T_1690; // @[Monitor.scala 648:68:freechips.rocketchip.system.DefaultRV32Config.fir@172619.6]
  wire [4:0] a_sizes_set_interm; // @[Monitor.scala 643:72:freechips.rocketchip.system.DefaultRV32Config.fir@172607.4]
  wire [19:0] _GEN_80; // @[Monitor.scala 648:43:freechips.rocketchip.system.DefaultRV32Config.fir@172620.6]
  wire [19:0] _T_1691; // @[Monitor.scala 648:43:freechips.rocketchip.system.DefaultRV32Config.fir@172620.6]
  wire [1:0] _T_1692; // @[Monitor.scala 649:26:freechips.rocketchip.system.DefaultRV32Config.fir@172622.6]
  wire  _T_1694; // @[Monitor.scala 649:17:freechips.rocketchip.system.DefaultRV32Config.fir@172624.6]
  wire  _T_1696; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@172626.6]
  wire  _T_1697; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@172627.6]
  wire [1:0] a_set; // @[Monitor.scala 643:72:freechips.rocketchip.system.DefaultRV32Config.fir@172607.4]
  wire [18:0] _GEN_30; // @[Monitor.scala 643:72:freechips.rocketchip.system.DefaultRV32Config.fir@172607.4]
  wire [19:0] _GEN_31; // @[Monitor.scala 643:72:freechips.rocketchip.system.DefaultRV32Config.fir@172607.4]
  wire  _T_1700; // @[Monitor.scala 660:27:freechips.rocketchip.system.DefaultRV32Config.fir@172641.4]
  wire  _T_1702; // @[Monitor.scala 660:75:freechips.rocketchip.system.DefaultRV32Config.fir@172643.4]
  wire  _T_1703; // @[Monitor.scala 660:72:freechips.rocketchip.system.DefaultRV32Config.fir@172644.4]
  wire [1:0] _T_1704; // @[OneHot.scala 58:35:freechips.rocketchip.system.DefaultRV32Config.fir@172646.6]
  wire [30:0] _GEN_82; // @[Monitor.scala 662:76:freechips.rocketchip.system.DefaultRV32Config.fir@172653.6]
  wire [30:0] _T_1710; // @[Monitor.scala 662:76:freechips.rocketchip.system.DefaultRV32Config.fir@172653.6]
  wire [30:0] _GEN_83; // @[Monitor.scala 663:72:freechips.rocketchip.system.DefaultRV32Config.fir@172660.6]
  wire [30:0] _T_1716; // @[Monitor.scala 663:72:freechips.rocketchip.system.DefaultRV32Config.fir@172660.6]
  wire [1:0] d_clr; // @[Monitor.scala 660:91:freechips.rocketchip.system.DefaultRV32Config.fir@172645.4]
  wire [30:0] _GEN_33; // @[Monitor.scala 660:91:freechips.rocketchip.system.DefaultRV32Config.fir@172645.4]
  wire [30:0] _GEN_34; // @[Monitor.scala 660:91:freechips.rocketchip.system.DefaultRV32Config.fir@172645.4]
  wire  _T_1717; // @[Monitor.scala 665:26:freechips.rocketchip.system.DefaultRV32Config.fir@172663.4]
  wire  _T_1720; // @[Monitor.scala 665:71:freechips.rocketchip.system.DefaultRV32Config.fir@172666.4]
  wire [1:0] _T_1721; // @[Monitor.scala 666:25:freechips.rocketchip.system.DefaultRV32Config.fir@172668.6]
  wire  _T_1723; // @[Monitor.scala 666:93:freechips.rocketchip.system.DefaultRV32Config.fir@172670.6]
  wire  _T_1724; // @[Monitor.scala 666:68:freechips.rocketchip.system.DefaultRV32Config.fir@172671.6]
  wire  _T_1725; // @[Monitor.scala 666:142:freechips.rocketchip.system.DefaultRV32Config.fir@172672.6]
  wire  _T_1726; // @[Monitor.scala 666:119:freechips.rocketchip.system.DefaultRV32Config.fir@172673.6]
  wire  _T_1727; // @[Monitor.scala 666:166:freechips.rocketchip.system.DefaultRV32Config.fir@172674.6]
  wire  _T_1728; // @[Monitor.scala 666:49:freechips.rocketchip.system.DefaultRV32Config.fir@172675.6]
  wire  _T_1730; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@172677.6]
  wire  _T_1731; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@172678.6]
  wire [3:0] a_opcode_lookup; // @[:freechips.rocketchip.system.DefaultRV32Config.fir@172560.4 :freechips.rocketchip.system.DefaultRV32Config.fir@172561.4 Monitor.scala 629:21:freechips.rocketchip.system.DefaultRV32Config.fir@172570.4]
  wire [2:0] _GEN_37; // @[Monitor.scala 667:37:freechips.rocketchip.system.DefaultRV32Config.fir@172684.6]
  wire [2:0] _GEN_38; // @[Monitor.scala 667:37:freechips.rocketchip.system.DefaultRV32Config.fir@172684.6]
  wire [2:0] _GEN_39; // @[Monitor.scala 667:37:freechips.rocketchip.system.DefaultRV32Config.fir@172684.6]
  wire [2:0] _GEN_40; // @[Monitor.scala 667:37:freechips.rocketchip.system.DefaultRV32Config.fir@172684.6]
  wire [2:0] _GEN_41; // @[Monitor.scala 667:37:freechips.rocketchip.system.DefaultRV32Config.fir@172684.6]
  wire [2:0] _GEN_42; // @[Monitor.scala 667:37:freechips.rocketchip.system.DefaultRV32Config.fir@172684.6]
  wire  _T_1733; // @[Monitor.scala 667:37:freechips.rocketchip.system.DefaultRV32Config.fir@172684.6]
  wire [2:0] _GEN_49; // @[Monitor.scala 667:96:freechips.rocketchip.system.DefaultRV32Config.fir@172686.6]
  wire [2:0] _GEN_50; // @[Monitor.scala 667:96:freechips.rocketchip.system.DefaultRV32Config.fir@172686.6]
  wire  _T_1735; // @[Monitor.scala 667:96:freechips.rocketchip.system.DefaultRV32Config.fir@172686.6]
  wire  _T_1736; // @[Monitor.scala 667:71:freechips.rocketchip.system.DefaultRV32Config.fir@172687.6]
  wire [2:0] _GEN_53; // @[Monitor.scala 668:60:freechips.rocketchip.system.DefaultRV32Config.fir@172688.6]
  wire [2:0] _GEN_54; // @[Monitor.scala 668:60:freechips.rocketchip.system.DefaultRV32Config.fir@172688.6]
  wire [2:0] _GEN_55; // @[Monitor.scala 668:60:freechips.rocketchip.system.DefaultRV32Config.fir@172688.6]
  wire [2:0] _GEN_56; // @[Monitor.scala 668:60:freechips.rocketchip.system.DefaultRV32Config.fir@172688.6]
  wire [2:0] _GEN_57; // @[Monitor.scala 668:60:freechips.rocketchip.system.DefaultRV32Config.fir@172688.6]
  wire [2:0] _GEN_58; // @[Monitor.scala 668:60:freechips.rocketchip.system.DefaultRV32Config.fir@172688.6]
  wire  _T_1737; // @[Monitor.scala 668:60:freechips.rocketchip.system.DefaultRV32Config.fir@172688.6]
  wire [2:0] _GEN_65; // @[Monitor.scala 668:124:freechips.rocketchip.system.DefaultRV32Config.fir@172689.6]
  wire [2:0] _GEN_66; // @[Monitor.scala 668:124:freechips.rocketchip.system.DefaultRV32Config.fir@172689.6]
  wire  _T_1738; // @[Monitor.scala 668:124:freechips.rocketchip.system.DefaultRV32Config.fir@172689.6]
  wire  _T_1739; // @[Monitor.scala 668:99:freechips.rocketchip.system.DefaultRV32Config.fir@172690.6]
  wire  _T_1740; // @[Monitor.scala 668:34:freechips.rocketchip.system.DefaultRV32Config.fir@172691.6]
  wire  _T_1741; // @[Monitor.scala 668:15:freechips.rocketchip.system.DefaultRV32Config.fir@172692.6]
  wire  _T_1743; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@172694.6]
  wire  _T_1744; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@172695.6]
  wire [7:0] a_size_lookup; // @[:freechips.rocketchip.system.DefaultRV32Config.fir@172571.4 :freechips.rocketchip.system.DefaultRV32Config.fir@172572.4 Monitor.scala 633:19:freechips.rocketchip.system.DefaultRV32Config.fir@172581.4]
  wire [7:0] _GEN_84; // @[Monitor.scala 670:34:freechips.rocketchip.system.DefaultRV32Config.fir@172700.6]
  wire  _T_1745; // @[Monitor.scala 670:34:freechips.rocketchip.system.DefaultRV32Config.fir@172700.6]
  wire  _T_1747; // @[Monitor.scala 670:72:freechips.rocketchip.system.DefaultRV32Config.fir@172702.6]
  wire  _T_1748; // @[Monitor.scala 670:53:freechips.rocketchip.system.DefaultRV32Config.fir@172703.6]
  wire  _T_1750; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@172705.6]
  wire  _T_1751; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@172706.6]
  wire  _T_1753; // @[Monitor.scala 672:36:freechips.rocketchip.system.DefaultRV32Config.fir@172713.4]
  wire  _T_1754; // @[Monitor.scala 672:47:freechips.rocketchip.system.DefaultRV32Config.fir@172714.4]
  wire  _T_1756; // @[Monitor.scala 672:65:freechips.rocketchip.system.DefaultRV32Config.fir@172716.4]
  wire  _T_1758; // @[Monitor.scala 672:116:freechips.rocketchip.system.DefaultRV32Config.fir@172718.4]
  wire  _T_1759; // @[Monitor.scala 673:15:freechips.rocketchip.system.DefaultRV32Config.fir@172720.6]
  wire  _T_1760; // @[Monitor.scala 673:32:freechips.rocketchip.system.DefaultRV32Config.fir@172721.6]
  wire  _T_1762; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@172723.6]
  wire  _T_1763; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@172724.6]
  wire  _T_1764; // @[Monitor.scala 677:20:freechips.rocketchip.system.DefaultRV32Config.fir@172730.4]
  wire  _T_1765; // @[Monitor.scala 677:40:freechips.rocketchip.system.DefaultRV32Config.fir@172731.4]
  wire  _T_1766; // @[Monitor.scala 677:33:freechips.rocketchip.system.DefaultRV32Config.fir@172732.4]
  wire  _T_1767; // @[Monitor.scala 677:30:freechips.rocketchip.system.DefaultRV32Config.fir@172733.4]
  wire  _T_1769; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@172735.4]
  wire  _T_1770; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@172736.4]
  wire [1:0] _T_1771; // @[Monitor.scala 680:27:freechips.rocketchip.system.DefaultRV32Config.fir@172741.4]
  wire [1:0] _T_1772; // @[Monitor.scala 680:38:freechips.rocketchip.system.DefaultRV32Config.fir@172742.4]
  wire [1:0] _T_1773; // @[Monitor.scala 680:36:freechips.rocketchip.system.DefaultRV32Config.fir@172743.4]
  wire [7:0] a_opcodes_set; // @[:freechips.rocketchip.system.DefaultRV32Config.fir@172556.4 :freechips.rocketchip.system.DefaultRV32Config.fir@172557.4 Monitor.scala 647:21:freechips.rocketchip.system.DefaultRV32Config.fir@172618.6]
  wire [7:0] _T_1774; // @[Monitor.scala 681:43:freechips.rocketchip.system.DefaultRV32Config.fir@172745.4]
  wire [7:0] d_opcodes_clr; // @[:freechips.rocketchip.system.DefaultRV32Config.fir@172635.4 :freechips.rocketchip.system.DefaultRV32Config.fir@172636.4 Monitor.scala 662:21:freechips.rocketchip.system.DefaultRV32Config.fir@172654.6]
  wire [7:0] _T_1775; // @[Monitor.scala 681:62:freechips.rocketchip.system.DefaultRV32Config.fir@172746.4]
  wire [7:0] _T_1776; // @[Monitor.scala 681:60:freechips.rocketchip.system.DefaultRV32Config.fir@172747.4]
  wire [15:0] a_sizes_set; // @[:freechips.rocketchip.system.DefaultRV32Config.fir@172558.4 :freechips.rocketchip.system.DefaultRV32Config.fir@172559.4 Monitor.scala 648:19:freechips.rocketchip.system.DefaultRV32Config.fir@172621.6]
  wire [15:0] _T_1777; // @[Monitor.scala 682:39:freechips.rocketchip.system.DefaultRV32Config.fir@172749.4]
  wire [15:0] d_sizes_clr; // @[:freechips.rocketchip.system.DefaultRV32Config.fir@172637.4 :freechips.rocketchip.system.DefaultRV32Config.fir@172638.4 Monitor.scala 663:19:freechips.rocketchip.system.DefaultRV32Config.fir@172661.6]
  wire [15:0] _T_1778; // @[Monitor.scala 682:56:freechips.rocketchip.system.DefaultRV32Config.fir@172750.4]
  wire [15:0] _T_1779; // @[Monitor.scala 682:54:freechips.rocketchip.system.DefaultRV32Config.fir@172751.4]
  reg [31:0] _T_1780; // @[Monitor.scala 684:27:freechips.rocketchip.system.DefaultRV32Config.fir@172753.4]
  wire  _T_1781; // @[Monitor.scala 687:26:freechips.rocketchip.system.DefaultRV32Config.fir@172756.4]
  wire  _T_1782; // @[Monitor.scala 687:16:freechips.rocketchip.system.DefaultRV32Config.fir@172757.4]
  wire  _T_1783; // @[Monitor.scala 687:39:freechips.rocketchip.system.DefaultRV32Config.fir@172758.4]
  wire  _T_1784; // @[Monitor.scala 687:30:freechips.rocketchip.system.DefaultRV32Config.fir@172759.4]
  wire  _T_1785; // @[Monitor.scala 687:59:freechips.rocketchip.system.DefaultRV32Config.fir@172760.4]
  wire  _T_1786; // @[Monitor.scala 687:47:freechips.rocketchip.system.DefaultRV32Config.fir@172761.4]
  wire  _T_1788; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@172763.4]
  wire  _T_1789; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@172764.4]
  wire [31:0] _T_1791; // @[Monitor.scala 689:26:freechips.rocketchip.system.DefaultRV32Config.fir@172770.4]
  wire  _T_1794; // @[Monitor.scala 690:27:freechips.rocketchip.system.DefaultRV32Config.fir@172774.4]
  reg [3:0] _T_1795; // @[Monitor.scala 694:27:freechips.rocketchip.system.DefaultRV32Config.fir@172778.4]
  reg [9:0] _T_1804; // @[Edges.scala 230:27:freechips.rocketchip.system.DefaultRV32Config.fir@172787.4]
  wire [9:0] _T_1806; // @[Edges.scala 231:28:freechips.rocketchip.system.DefaultRV32Config.fir@172789.4]
  wire  _T_1807; // @[Edges.scala 232:25:freechips.rocketchip.system.DefaultRV32Config.fir@172790.4]
  wire  _T_1817; // @[Monitor.scala 700:27:freechips.rocketchip.system.DefaultRV32Config.fir@172804.4]
  wire  _T_1820; // @[Edges.scala 72:43:freechips.rocketchip.system.DefaultRV32Config.fir@172807.4]
  wire  _T_1821; // @[Edges.scala 72:40:freechips.rocketchip.system.DefaultRV32Config.fir@172808.4]
  wire  _T_1822; // @[Monitor.scala 700:38:freechips.rocketchip.system.DefaultRV32Config.fir@172809.4]
  wire [3:0] _T_1823; // @[OneHot.scala 58:35:freechips.rocketchip.system.DefaultRV32Config.fir@172811.6]
  wire [3:0] _T_1824; // @[Monitor.scala 702:23:freechips.rocketchip.system.DefaultRV32Config.fir@172813.6]
  wire  _T_1826; // @[Monitor.scala 702:14:freechips.rocketchip.system.DefaultRV32Config.fir@172815.6]
  wire  _T_1828; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@172817.6]
  wire  _T_1829; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@172818.6]
  wire [3:0] _GEN_69; // @[Monitor.scala 700:72:freechips.rocketchip.system.DefaultRV32Config.fir@172810.4]
  wire  _T_1831; // @[Decoupled.scala 40:37:freechips.rocketchip.system.DefaultRV32Config.fir@172826.4]
  wire [3:0] _T_1834; // @[OneHot.scala 58:35:freechips.rocketchip.system.DefaultRV32Config.fir@172830.6]
  wire [3:0] _T_1835; // @[Monitor.scala 708:24:freechips.rocketchip.system.DefaultRV32Config.fir@172832.6]
  wire [3:0] _T_1836; // @[Monitor.scala 708:35:freechips.rocketchip.system.DefaultRV32Config.fir@172833.6]
  wire  _T_1839; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@172836.6]
  wire  _T_1840; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@172837.6]
  wire [3:0] _GEN_70; // @[Monitor.scala 706:73:freechips.rocketchip.system.DefaultRV32Config.fir@172829.4]
  wire [3:0] _T_1841; // @[Monitor.scala 713:27:freechips.rocketchip.system.DefaultRV32Config.fir@172843.4]
  wire [3:0] _T_1842; // @[Monitor.scala 713:38:freechips.rocketchip.system.DefaultRV32Config.fir@172844.4]
  wire [3:0] _T_1843; // @[Monitor.scala 713:36:freechips.rocketchip.system.DefaultRV32Config.fir@172845.4]
  wire  _GEN_85; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@170087.10]
  wire  _GEN_99; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@170212.10]
  wire  _GEN_115; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@170348.10]
  wire  _GEN_125; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@170455.10]
  wire  _GEN_135; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@170554.10]
  wire  _GEN_145; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@170645.10]
  wire  _GEN_155; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@170734.10]
  wire  _GEN_165; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@170823.10]
  wire  _GEN_175; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@170889.10]
  wire  _GEN_185; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@170931.10]
  wire  _GEN_195; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@170989.10]
  wire  _GEN_205; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@171048.10]
  wire  _GEN_211; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@171083.10]
  wire  _GEN_217; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@171119.10]
  wire  _GEN_223; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@171301.10]
  wire  _GEN_235; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@171356.10]
  wire  _GEN_247; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@171411.10]
  wire  _GEN_257; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@171458.10]
  wire  _GEN_267; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@171507.10]
  wire  _GEN_275; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@171554.10]
  wire  _GEN_283; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@171601.10]
  wire  _GEN_293; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@171745.10]
  wire  _GEN_303; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@171793.10]
  wire  _GEN_313; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@171882.10]
  wire  _GEN_325; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@171998.10]
  wire  _GEN_337; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@172057.10]
  wire  _GEN_345; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@172097.10]
  wire  _GEN_353; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@172129.10]
  plusarg_reader #(.FORMAT("tilelink_timeout=%d"), .DEFAULT(0), .WIDTH(32)) plusarg_reader ( // @[PlusArg.scala 80:11:freechips.rocketchip.system.DefaultRV32Config.fir@172754.4]
    .out(plusarg_reader_out)
  );
  assign _T_4 = ~io_in_a_bits_source; // @[Parameters.scala 47:9:freechips.rocketchip.system.DefaultRV32Config.fir@169962.6]
  assign _T_7 = _T_4 | io_in_a_bits_source; // @[Parameters.scala 924:46:freechips.rocketchip.system.DefaultRV32Config.fir@169968.6]
  assign _T_9 = 27'hfff << io_in_a_bits_size; // @[package.scala 207:77:freechips.rocketchip.system.DefaultRV32Config.fir@169970.6]
  assign _T_11 = ~_T_9[11:0]; // @[package.scala 207:46:freechips.rocketchip.system.DefaultRV32Config.fir@169972.6]
  assign _GEN_71 = {{20'd0}, _T_11}; // @[Edges.scala 22:16:freechips.rocketchip.system.DefaultRV32Config.fir@169973.6]
  assign _T_12 = io_in_a_bits_address & _GEN_71; // @[Edges.scala 22:16:freechips.rocketchip.system.DefaultRV32Config.fir@169973.6]
  assign _T_13 = _T_12 == 32'h0; // @[Edges.scala 22:24:freechips.rocketchip.system.DefaultRV32Config.fir@169974.6]
  assign _T_16 = 2'h1 << io_in_a_bits_size[0]; // @[OneHot.scala 65:12:freechips.rocketchip.system.DefaultRV32Config.fir@169977.6]
  assign _T_18 = _T_16 | 2'h1; // @[Misc.scala 201:81:freechips.rocketchip.system.DefaultRV32Config.fir@169979.6]
  assign _T_19 = io_in_a_bits_size >= 4'h2; // @[Misc.scala 205:21:freechips.rocketchip.system.DefaultRV32Config.fir@169980.6]
  assign _T_22 = ~io_in_a_bits_address[1]; // @[Misc.scala 210:20:freechips.rocketchip.system.DefaultRV32Config.fir@169983.6]
  assign _T_24 = _T_18[1] & _T_22; // @[Misc.scala 214:38:freechips.rocketchip.system.DefaultRV32Config.fir@169985.6]
  assign _T_25 = _T_19 | _T_24; // @[Misc.scala 214:29:freechips.rocketchip.system.DefaultRV32Config.fir@169986.6]
  assign _T_27 = _T_18[1] & io_in_a_bits_address[1]; // @[Misc.scala 214:38:freechips.rocketchip.system.DefaultRV32Config.fir@169988.6]
  assign _T_28 = _T_19 | _T_27; // @[Misc.scala 214:29:freechips.rocketchip.system.DefaultRV32Config.fir@169989.6]
  assign _T_31 = ~io_in_a_bits_address[0]; // @[Misc.scala 210:20:freechips.rocketchip.system.DefaultRV32Config.fir@169992.6]
  assign _T_32 = _T_22 & _T_31; // @[Misc.scala 213:27:freechips.rocketchip.system.DefaultRV32Config.fir@169993.6]
  assign _T_33 = _T_18[0] & _T_32; // @[Misc.scala 214:38:freechips.rocketchip.system.DefaultRV32Config.fir@169994.6]
  assign _T_34 = _T_25 | _T_33; // @[Misc.scala 214:29:freechips.rocketchip.system.DefaultRV32Config.fir@169995.6]
  assign _T_35 = _T_22 & io_in_a_bits_address[0]; // @[Misc.scala 213:27:freechips.rocketchip.system.DefaultRV32Config.fir@169996.6]
  assign _T_36 = _T_18[0] & _T_35; // @[Misc.scala 214:38:freechips.rocketchip.system.DefaultRV32Config.fir@169997.6]
  assign _T_37 = _T_25 | _T_36; // @[Misc.scala 214:29:freechips.rocketchip.system.DefaultRV32Config.fir@169998.6]
  assign _T_38 = io_in_a_bits_address[1] & _T_31; // @[Misc.scala 213:27:freechips.rocketchip.system.DefaultRV32Config.fir@169999.6]
  assign _T_39 = _T_18[0] & _T_38; // @[Misc.scala 214:38:freechips.rocketchip.system.DefaultRV32Config.fir@170000.6]
  assign _T_40 = _T_28 | _T_39; // @[Misc.scala 214:29:freechips.rocketchip.system.DefaultRV32Config.fir@170001.6]
  assign _T_41 = io_in_a_bits_address[1] & io_in_a_bits_address[0]; // @[Misc.scala 213:27:freechips.rocketchip.system.DefaultRV32Config.fir@170002.6]
  assign _T_42 = _T_18[0] & _T_41; // @[Misc.scala 214:38:freechips.rocketchip.system.DefaultRV32Config.fir@170003.6]
  assign _T_43 = _T_28 | _T_42; // @[Misc.scala 214:29:freechips.rocketchip.system.DefaultRV32Config.fir@170004.6]
  assign _T_46 = {_T_43,_T_40,_T_37,_T_34}; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@170007.6]
  assign _T_50 = {1'b0,$signed(io_in_a_bits_address)}; // @[Parameters.scala 137:49:freechips.rocketchip.system.DefaultRV32Config.fir@170011.6]
  assign _T_67 = io_in_a_bits_opcode == 3'h6; // @[Monitor.scala 79:25:freechips.rocketchip.system.DefaultRV32Config.fir@170032.6]
  assign _T_72 = $signed(_T_50) & -33'sh1000; // @[Parameters.scala 137:52:freechips.rocketchip.system.DefaultRV32Config.fir@170038.8]
  assign _T_73 = $signed(_T_72) == 33'sh0; // @[Parameters.scala 137:67:freechips.rocketchip.system.DefaultRV32Config.fir@170039.8]
  assign _T_74 = io_in_a_bits_address ^ 32'h3000; // @[Parameters.scala 137:31:freechips.rocketchip.system.DefaultRV32Config.fir@170040.8]
  assign _T_75 = {1'b0,$signed(_T_74)}; // @[Parameters.scala 137:49:freechips.rocketchip.system.DefaultRV32Config.fir@170041.8]
  assign _T_77 = $signed(_T_75) & -33'sh1000; // @[Parameters.scala 137:52:freechips.rocketchip.system.DefaultRV32Config.fir@170043.8]
  assign _T_78 = $signed(_T_77) == 33'sh0; // @[Parameters.scala 137:67:freechips.rocketchip.system.DefaultRV32Config.fir@170044.8]
  assign _T_79 = io_in_a_bits_address ^ 32'h10000; // @[Parameters.scala 137:31:freechips.rocketchip.system.DefaultRV32Config.fir@170045.8]
  assign _T_80 = {1'b0,$signed(_T_79)}; // @[Parameters.scala 137:49:freechips.rocketchip.system.DefaultRV32Config.fir@170046.8]
  assign _T_82 = $signed(_T_80) & -33'sh10000; // @[Parameters.scala 137:52:freechips.rocketchip.system.DefaultRV32Config.fir@170048.8]
  assign _T_83 = $signed(_T_82) == 33'sh0; // @[Parameters.scala 137:67:freechips.rocketchip.system.DefaultRV32Config.fir@170049.8]
  assign _T_84 = io_in_a_bits_address ^ 32'h2000000; // @[Parameters.scala 137:31:freechips.rocketchip.system.DefaultRV32Config.fir@170050.8]
  assign _T_85 = {1'b0,$signed(_T_84)}; // @[Parameters.scala 137:49:freechips.rocketchip.system.DefaultRV32Config.fir@170051.8]
  assign _T_87 = $signed(_T_85) & -33'sh10000; // @[Parameters.scala 137:52:freechips.rocketchip.system.DefaultRV32Config.fir@170053.8]
  assign _T_88 = $signed(_T_87) == 33'sh0; // @[Parameters.scala 137:67:freechips.rocketchip.system.DefaultRV32Config.fir@170054.8]
  assign _T_89 = io_in_a_bits_address ^ 32'hc000000; // @[Parameters.scala 137:31:freechips.rocketchip.system.DefaultRV32Config.fir@170055.8]
  assign _T_90 = {1'b0,$signed(_T_89)}; // @[Parameters.scala 137:49:freechips.rocketchip.system.DefaultRV32Config.fir@170056.8]
  assign _T_92 = $signed(_T_90) & -33'sh4000000; // @[Parameters.scala 137:52:freechips.rocketchip.system.DefaultRV32Config.fir@170058.8]
  assign _T_93 = $signed(_T_92) == 33'sh0; // @[Parameters.scala 137:67:freechips.rocketchip.system.DefaultRV32Config.fir@170059.8]
  assign _T_94 = io_in_a_bits_address ^ 32'h60000000; // @[Parameters.scala 137:31:freechips.rocketchip.system.DefaultRV32Config.fir@170060.8]
  assign _T_95 = {1'b0,$signed(_T_94)}; // @[Parameters.scala 137:49:freechips.rocketchip.system.DefaultRV32Config.fir@170061.8]
  assign _T_97 = $signed(_T_95) & -33'sh20000000; // @[Parameters.scala 137:52:freechips.rocketchip.system.DefaultRV32Config.fir@170063.8]
  assign _T_98 = $signed(_T_97) == 33'sh0; // @[Parameters.scala 137:67:freechips.rocketchip.system.DefaultRV32Config.fir@170064.8]
  assign _T_99 = _T_73 | _T_78; // @[Parameters.scala 552:42:freechips.rocketchip.system.DefaultRV32Config.fir@170065.8]
  assign _T_106 = io_in_a_bits_size <= 4'h6; // @[Parameters.scala 93:42:freechips.rocketchip.system.DefaultRV32Config.fir@170072.8]
  assign _T_109 = io_in_a_bits_address ^ 32'h80000000; // @[Parameters.scala 137:31:freechips.rocketchip.system.DefaultRV32Config.fir@170075.8]
  assign _T_110 = {1'b0,$signed(_T_109)}; // @[Parameters.scala 137:49:freechips.rocketchip.system.DefaultRV32Config.fir@170076.8]
  assign _T_112 = $signed(_T_110) & -33'sh10000000; // @[Parameters.scala 137:52:freechips.rocketchip.system.DefaultRV32Config.fir@170078.8]
  assign _T_113 = $signed(_T_112) == 33'sh0; // @[Parameters.scala 137:67:freechips.rocketchip.system.DefaultRV32Config.fir@170079.8]
  assign _T_114 = _T_106 & _T_113; // @[Parameters.scala 551:56:freechips.rocketchip.system.DefaultRV32Config.fir@170080.8]
  assign _T_118 = _T_114 | reset; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@170084.8]
  assign _T_119 = ~_T_118; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@170085.8]
  assign _T_123 = 4'h6 == io_in_a_bits_size; // @[Parameters.scala 92:48:freechips.rocketchip.system.DefaultRV32Config.fir@170096.8]
  assign _T_124 = _T_4 & _T_123; // @[Mux.scala 27:72:freechips.rocketchip.system.DefaultRV32Config.fir@170097.8]
  assign _T_129 = _T_124 | reset; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@170103.8]
  assign _T_130 = ~_T_129; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@170104.8]
  assign _T_132 = _T_7 | reset; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@170110.8]
  assign _T_133 = ~_T_132; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@170111.8]
  assign _T_136 = _T_19 | reset; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@170118.8]
  assign _T_137 = ~_T_136; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@170119.8]
  assign _T_139 = _T_13 | reset; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@170125.8]
  assign _T_140 = ~_T_139; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@170126.8]
  assign _T_141 = io_in_a_bits_param <= 3'h2; // @[Bundles.scala 110:27:freechips.rocketchip.system.DefaultRV32Config.fir@170131.8]
  assign _T_143 = _T_141 | reset; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@170133.8]
  assign _T_144 = ~_T_143; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@170134.8]
  assign _T_145 = ~io_in_a_bits_mask; // @[Monitor.scala 86:18:freechips.rocketchip.system.DefaultRV32Config.fir@170139.8]
  assign _T_146 = _T_145 == 4'h0; // @[Monitor.scala 86:31:freechips.rocketchip.system.DefaultRV32Config.fir@170140.8]
  assign _T_148 = _T_146 | reset; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@170142.8]
  assign _T_149 = ~_T_148; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@170143.8]
  assign _T_154 = io_in_a_bits_opcode == 3'h7; // @[Monitor.scala 90:25:freechips.rocketchip.system.DefaultRV32Config.fir@170157.6]
  assign _T_232 = io_in_a_bits_param != 3'h0; // @[Monitor.scala 97:31:freechips.rocketchip.system.DefaultRV32Config.fir@170264.8]
  assign _T_234 = _T_232 | reset; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@170266.8]
  assign _T_235 = ~_T_234; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@170267.8]
  assign _T_245 = io_in_a_bits_opcode == 3'h4; // @[Monitor.scala 102:25:freechips.rocketchip.system.DefaultRV32Config.fir@170290.6]
  assign _T_247 = io_in_a_bits_size <= 4'hc; // @[Parameters.scala 93:42:freechips.rocketchip.system.DefaultRV32Config.fir@170293.8]
  assign _T_255 = _T_247 & _T_78; // @[Parameters.scala 551:56:freechips.rocketchip.system.DefaultRV32Config.fir@170301.8]
  assign _T_290 = _T_73 | _T_83; // @[Parameters.scala 552:42:freechips.rocketchip.system.DefaultRV32Config.fir@170336.8]
  assign _T_291 = _T_290 | _T_88; // @[Parameters.scala 552:42:freechips.rocketchip.system.DefaultRV32Config.fir@170337.8]
  assign _T_292 = _T_291 | _T_93; // @[Parameters.scala 552:42:freechips.rocketchip.system.DefaultRV32Config.fir@170338.8]
  assign _T_293 = _T_292 | _T_98; // @[Parameters.scala 552:42:freechips.rocketchip.system.DefaultRV32Config.fir@170339.8]
  assign _T_294 = _T_293 | _T_113; // @[Parameters.scala 552:42:freechips.rocketchip.system.DefaultRV32Config.fir@170340.8]
  assign _T_295 = _T_106 & _T_294; // @[Parameters.scala 551:56:freechips.rocketchip.system.DefaultRV32Config.fir@170341.8]
  assign _T_297 = _T_255 | _T_295; // @[Parameters.scala 553:30:freechips.rocketchip.system.DefaultRV32Config.fir@170343.8]
  assign _T_299 = _T_297 | reset; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@170345.8]
  assign _T_300 = ~_T_299; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@170346.8]
  assign _T_307 = io_in_a_bits_param == 3'h0; // @[Monitor.scala 106:31:freechips.rocketchip.system.DefaultRV32Config.fir@170365.8]
  assign _T_309 = _T_307 | reset; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@170367.8]
  assign _T_310 = ~_T_309; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@170368.8]
  assign _T_311 = io_in_a_bits_mask == _T_46; // @[Monitor.scala 107:30:freechips.rocketchip.system.DefaultRV32Config.fir@170373.8]
  assign _T_313 = _T_311 | reset; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@170375.8]
  assign _T_314 = ~_T_313; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@170376.8]
  assign _T_319 = io_in_a_bits_opcode == 3'h0; // @[Monitor.scala 111:25:freechips.rocketchip.system.DefaultRV32Config.fir@170390.6]
  assign _T_354 = _T_73 | _T_88; // @[Parameters.scala 552:42:freechips.rocketchip.system.DefaultRV32Config.fir@170426.8]
  assign _T_355 = _T_354 | _T_93; // @[Parameters.scala 552:42:freechips.rocketchip.system.DefaultRV32Config.fir@170427.8]
  assign _T_356 = _T_355 | _T_113; // @[Parameters.scala 552:42:freechips.rocketchip.system.DefaultRV32Config.fir@170428.8]
  assign _T_357 = _T_106 & _T_356; // @[Parameters.scala 551:56:freechips.rocketchip.system.DefaultRV32Config.fir@170429.8]
  assign _T_366 = io_in_a_bits_size <= 4'h8; // @[Parameters.scala 93:42:freechips.rocketchip.system.DefaultRV32Config.fir@170438.8]
  assign _T_374 = _T_366 & _T_98; // @[Parameters.scala 551:56:freechips.rocketchip.system.DefaultRV32Config.fir@170446.8]
  assign _T_376 = _T_255 | _T_357; // @[Parameters.scala 553:30:freechips.rocketchip.system.DefaultRV32Config.fir@170448.8]
  assign _T_378 = _T_376 | _T_374; // @[Parameters.scala 553:30:freechips.rocketchip.system.DefaultRV32Config.fir@170450.8]
  assign _T_380 = _T_378 | reset; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@170452.8]
  assign _T_381 = ~_T_380; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@170453.8]
  assign _T_396 = io_in_a_bits_opcode == 3'h1; // @[Monitor.scala 119:25:freechips.rocketchip.system.DefaultRV32Config.fir@170489.6]
  assign _T_469 = ~_T_46; // @[Monitor.scala 124:33:freechips.rocketchip.system.DefaultRV32Config.fir@170579.8]
  assign _T_470 = io_in_a_bits_mask & _T_469; // @[Monitor.scala 124:31:freechips.rocketchip.system.DefaultRV32Config.fir@170580.8]
  assign _T_471 = _T_470 == 4'h0; // @[Monitor.scala 124:40:freechips.rocketchip.system.DefaultRV32Config.fir@170581.8]
  assign _T_473 = _T_471 | reset; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@170583.8]
  assign _T_474 = ~_T_473; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@170584.8]
  assign _T_475 = io_in_a_bits_opcode == 3'h2; // @[Monitor.scala 127:25:freechips.rocketchip.system.DefaultRV32Config.fir@170590.6]
  assign _T_477 = io_in_a_bits_size <= 4'h2; // @[Parameters.scala 93:42:freechips.rocketchip.system.DefaultRV32Config.fir@170593.8]
  assign _T_501 = _T_99 | _T_88; // @[Parameters.scala 552:42:freechips.rocketchip.system.DefaultRV32Config.fir@170617.8]
  assign _T_502 = _T_501 | _T_93; // @[Parameters.scala 552:42:freechips.rocketchip.system.DefaultRV32Config.fir@170618.8]
  assign _T_503 = _T_477 & _T_502; // @[Parameters.scala 551:56:freechips.rocketchip.system.DefaultRV32Config.fir@170619.8]
  assign _T_526 = _T_503 | reset; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@170642.8]
  assign _T_527 = ~_T_526; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@170643.8]
  assign _T_534 = io_in_a_bits_param <= 3'h4; // @[Bundles.scala 140:33:freechips.rocketchip.system.DefaultRV32Config.fir@170662.8]
  assign _T_536 = _T_534 | reset; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@170664.8]
  assign _T_537 = ~_T_536; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@170665.8]
  assign _T_542 = io_in_a_bits_opcode == 3'h3; // @[Monitor.scala 135:25:freechips.rocketchip.system.DefaultRV32Config.fir@170679.6]
  assign _T_601 = io_in_a_bits_param <= 3'h3; // @[Bundles.scala 147:30:freechips.rocketchip.system.DefaultRV32Config.fir@170751.8]
  assign _T_603 = _T_601 | reset; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@170753.8]
  assign _T_604 = ~_T_603; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@170754.8]
  assign _T_609 = io_in_a_bits_opcode == 3'h5; // @[Monitor.scala 143:25:freechips.rocketchip.system.DefaultRV32Config.fir@170768.6]
  assign _T_660 = _T_255 | reset; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@170820.8]
  assign _T_661 = ~_T_660; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@170821.8]
  assign _T_668 = io_in_a_bits_param <= 3'h1; // @[Bundles.scala 160:28:freechips.rocketchip.system.DefaultRV32Config.fir@170840.8]
  assign _T_670 = _T_668 | reset; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@170842.8]
  assign _T_671 = ~_T_670; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@170843.8]
  assign _T_680 = io_in_d_bits_opcode <= 3'h6; // @[Bundles.scala 44:24:freechips.rocketchip.system.DefaultRV32Config.fir@170867.6]
  assign _T_682 = _T_680 | reset; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@170869.6]
  assign _T_683 = ~_T_682; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@170870.6]
  assign _T_684 = ~io_in_d_bits_source; // @[Parameters.scala 47:9:freechips.rocketchip.system.DefaultRV32Config.fir@170875.6]
  assign _T_687 = _T_684 | io_in_d_bits_source; // @[Parameters.scala 924:46:freechips.rocketchip.system.DefaultRV32Config.fir@170881.6]
  assign _T_689 = io_in_d_bits_opcode == 3'h6; // @[Monitor.scala 307:25:freechips.rocketchip.system.DefaultRV32Config.fir@170883.6]
  assign _T_691 = _T_687 | reset; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@170886.8]
  assign _T_692 = ~_T_691; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@170887.8]
  assign _T_693 = io_in_d_bits_size >= 4'h2; // @[Monitor.scala 309:27:freechips.rocketchip.system.DefaultRV32Config.fir@170892.8]
  assign _T_695 = _T_693 | reset; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@170894.8]
  assign _T_696 = ~_T_695; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@170895.8]
  assign _T_697 = io_in_d_bits_param == 2'h0; // @[Monitor.scala 310:28:freechips.rocketchip.system.DefaultRV32Config.fir@170900.8]
  assign _T_699 = _T_697 | reset; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@170902.8]
  assign _T_700 = ~_T_699; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@170903.8]
  assign _T_701 = ~io_in_d_bits_corrupt; // @[Monitor.scala 311:15:freechips.rocketchip.system.DefaultRV32Config.fir@170908.8]
  assign _T_703 = _T_701 | reset; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@170910.8]
  assign _T_704 = ~_T_703; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@170911.8]
  assign _T_705 = ~io_in_d_bits_denied; // @[Monitor.scala 312:15:freechips.rocketchip.system.DefaultRV32Config.fir@170916.8]
  assign _T_707 = _T_705 | reset; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@170918.8]
  assign _T_708 = ~_T_707; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@170919.8]
  assign _T_709 = io_in_d_bits_opcode == 3'h4; // @[Monitor.scala 315:25:freechips.rocketchip.system.DefaultRV32Config.fir@170925.6]
  assign _T_720 = io_in_d_bits_param <= 2'h2; // @[Bundles.scala 104:26:freechips.rocketchip.system.DefaultRV32Config.fir@170949.8]
  assign _T_722 = _T_720 | reset; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@170951.8]
  assign _T_723 = ~_T_722; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@170952.8]
  assign _T_724 = io_in_d_bits_param != 2'h2; // @[Monitor.scala 320:28:freechips.rocketchip.system.DefaultRV32Config.fir@170957.8]
  assign _T_726 = _T_724 | reset; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@170959.8]
  assign _T_727 = ~_T_726; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@170960.8]
  assign _T_737 = io_in_d_bits_opcode == 3'h5; // @[Monitor.scala 325:25:freechips.rocketchip.system.DefaultRV32Config.fir@170983.6]
  assign _T_757 = _T_705 | io_in_d_bits_corrupt; // @[Monitor.scala 331:30:freechips.rocketchip.system.DefaultRV32Config.fir@171024.8]
  assign _T_759 = _T_757 | reset; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@171026.8]
  assign _T_760 = ~_T_759; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@171027.8]
  assign _T_766 = io_in_d_bits_opcode == 3'h0; // @[Monitor.scala 335:25:freechips.rocketchip.system.DefaultRV32Config.fir@171042.6]
  assign _T_783 = io_in_d_bits_opcode == 3'h1; // @[Monitor.scala 343:25:freechips.rocketchip.system.DefaultRV32Config.fir@171077.6]
  assign _T_801 = io_in_d_bits_opcode == 3'h2; // @[Monitor.scala 351:25:freechips.rocketchip.system.DefaultRV32Config.fir@171113.6]
  assign _T_818 = io_in_b_bits_opcode <= 3'h6; // @[Bundles.scala 42:24:freechips.rocketchip.system.DefaultRV32Config.fir@171150.6]
  assign _T_820 = _T_818 | reset; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@171152.6]
  assign _T_821 = ~_T_820; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@171153.6]
  assign _T_822 = ~io_in_b_bits_source; // @[Parameters.scala 47:9:freechips.rocketchip.system.DefaultRV32Config.fir@171158.6]
  assign _T_825 = {1'b0,$signed(io_in_b_bits_address)}; // @[Parameters.scala 137:49:freechips.rocketchip.system.DefaultRV32Config.fir@171161.6]
  assign _T_842 = io_in_b_bits_address ^ 32'h3000; // @[Parameters.scala 137:31:freechips.rocketchip.system.DefaultRV32Config.fir@171182.6]
  assign _T_843 = {1'b0,$signed(_T_842)}; // @[Parameters.scala 137:49:freechips.rocketchip.system.DefaultRV32Config.fir@171183.6]
  assign _T_845 = $signed(_T_843) & -33'sh1000; // @[Parameters.scala 137:52:freechips.rocketchip.system.DefaultRV32Config.fir@171185.6]
  assign _T_846 = $signed(_T_845) == 33'sh0; // @[Parameters.scala 137:67:freechips.rocketchip.system.DefaultRV32Config.fir@171186.6]
  assign _T_847 = io_in_b_bits_address ^ 32'hc000000; // @[Parameters.scala 137:31:freechips.rocketchip.system.DefaultRV32Config.fir@171187.6]
  assign _T_848 = {1'b0,$signed(_T_847)}; // @[Parameters.scala 137:49:freechips.rocketchip.system.DefaultRV32Config.fir@171188.6]
  assign _T_850 = $signed(_T_848) & -33'sh4000000; // @[Parameters.scala 137:52:freechips.rocketchip.system.DefaultRV32Config.fir@171190.6]
  assign _T_851 = $signed(_T_850) == 33'sh0; // @[Parameters.scala 137:67:freechips.rocketchip.system.DefaultRV32Config.fir@171191.6]
  assign _T_852 = io_in_b_bits_address ^ 32'h2000000; // @[Parameters.scala 137:31:freechips.rocketchip.system.DefaultRV32Config.fir@171192.6]
  assign _T_853 = {1'b0,$signed(_T_852)}; // @[Parameters.scala 137:49:freechips.rocketchip.system.DefaultRV32Config.fir@171193.6]
  assign _T_855 = $signed(_T_853) & -33'sh10000; // @[Parameters.scala 137:52:freechips.rocketchip.system.DefaultRV32Config.fir@171195.6]
  assign _T_856 = $signed(_T_855) == 33'sh0; // @[Parameters.scala 137:67:freechips.rocketchip.system.DefaultRV32Config.fir@171196.6]
  assign _T_860 = $signed(_T_825) & -33'sh1000; // @[Parameters.scala 137:52:freechips.rocketchip.system.DefaultRV32Config.fir@171200.6]
  assign _T_861 = $signed(_T_860) == 33'sh0; // @[Parameters.scala 137:67:freechips.rocketchip.system.DefaultRV32Config.fir@171201.6]
  assign _T_862 = io_in_b_bits_address ^ 32'h10000; // @[Parameters.scala 137:31:freechips.rocketchip.system.DefaultRV32Config.fir@171202.6]
  assign _T_863 = {1'b0,$signed(_T_862)}; // @[Parameters.scala 137:49:freechips.rocketchip.system.DefaultRV32Config.fir@171203.6]
  assign _T_865 = $signed(_T_863) & -33'sh10000; // @[Parameters.scala 137:52:freechips.rocketchip.system.DefaultRV32Config.fir@171205.6]
  assign _T_866 = $signed(_T_865) == 33'sh0; // @[Parameters.scala 137:67:freechips.rocketchip.system.DefaultRV32Config.fir@171206.6]
  assign _T_867 = io_in_b_bits_address ^ 32'h80000000; // @[Parameters.scala 137:31:freechips.rocketchip.system.DefaultRV32Config.fir@171207.6]
  assign _T_868 = {1'b0,$signed(_T_867)}; // @[Parameters.scala 137:49:freechips.rocketchip.system.DefaultRV32Config.fir@171208.6]
  assign _T_870 = $signed(_T_868) & -33'sh10000000; // @[Parameters.scala 137:52:freechips.rocketchip.system.DefaultRV32Config.fir@171210.6]
  assign _T_871 = $signed(_T_870) == 33'sh0; // @[Parameters.scala 137:67:freechips.rocketchip.system.DefaultRV32Config.fir@171211.6]
  assign _T_872 = io_in_b_bits_address ^ 32'h60000000; // @[Parameters.scala 137:31:freechips.rocketchip.system.DefaultRV32Config.fir@171212.6]
  assign _T_873 = {1'b0,$signed(_T_872)}; // @[Parameters.scala 137:49:freechips.rocketchip.system.DefaultRV32Config.fir@171213.6]
  assign _T_875 = $signed(_T_873) & -33'sh20000000; // @[Parameters.scala 137:52:freechips.rocketchip.system.DefaultRV32Config.fir@171215.6]
  assign _T_876 = $signed(_T_875) == 33'sh0; // @[Parameters.scala 137:67:freechips.rocketchip.system.DefaultRV32Config.fir@171216.6]
  assign _T_878 = _T_846 | _T_851; // @[Parameters.scala 535:64:freechips.rocketchip.system.DefaultRV32Config.fir@171226.6]
  assign _T_879 = _T_878 | _T_856; // @[Parameters.scala 535:64:freechips.rocketchip.system.DefaultRV32Config.fir@171227.6]
  assign _T_880 = _T_879 | _T_861; // @[Parameters.scala 535:64:freechips.rocketchip.system.DefaultRV32Config.fir@171228.6]
  assign _T_881 = _T_880 | _T_866; // @[Parameters.scala 535:64:freechips.rocketchip.system.DefaultRV32Config.fir@171229.6]
  assign _T_882 = _T_881 | _T_871; // @[Parameters.scala 535:64:freechips.rocketchip.system.DefaultRV32Config.fir@171230.6]
  assign _T_883 = _T_882 | _T_876; // @[Parameters.scala 535:64:freechips.rocketchip.system.DefaultRV32Config.fir@171231.6]
  assign _T_885 = 27'hfff << io_in_b_bits_size; // @[package.scala 207:77:freechips.rocketchip.system.DefaultRV32Config.fir@171233.6]
  assign _T_887 = ~_T_885[11:0]; // @[package.scala 207:46:freechips.rocketchip.system.DefaultRV32Config.fir@171235.6]
  assign _GEN_72 = {{20'd0}, _T_887}; // @[Edges.scala 22:16:freechips.rocketchip.system.DefaultRV32Config.fir@171236.6]
  assign _T_888 = io_in_b_bits_address & _GEN_72; // @[Edges.scala 22:16:freechips.rocketchip.system.DefaultRV32Config.fir@171236.6]
  assign _T_889 = _T_888 == 32'h0; // @[Edges.scala 22:24:freechips.rocketchip.system.DefaultRV32Config.fir@171237.6]
  assign _T_892 = 2'h1 << io_in_b_bits_size[0]; // @[OneHot.scala 65:12:freechips.rocketchip.system.DefaultRV32Config.fir@171240.6]
  assign _T_894 = _T_892 | 2'h1; // @[Misc.scala 201:81:freechips.rocketchip.system.DefaultRV32Config.fir@171242.6]
  assign _T_895 = io_in_b_bits_size >= 4'h2; // @[Misc.scala 205:21:freechips.rocketchip.system.DefaultRV32Config.fir@171243.6]
  assign _T_898 = ~io_in_b_bits_address[1]; // @[Misc.scala 210:20:freechips.rocketchip.system.DefaultRV32Config.fir@171246.6]
  assign _T_900 = _T_894[1] & _T_898; // @[Misc.scala 214:38:freechips.rocketchip.system.DefaultRV32Config.fir@171248.6]
  assign _T_901 = _T_895 | _T_900; // @[Misc.scala 214:29:freechips.rocketchip.system.DefaultRV32Config.fir@171249.6]
  assign _T_903 = _T_894[1] & io_in_b_bits_address[1]; // @[Misc.scala 214:38:freechips.rocketchip.system.DefaultRV32Config.fir@171251.6]
  assign _T_904 = _T_895 | _T_903; // @[Misc.scala 214:29:freechips.rocketchip.system.DefaultRV32Config.fir@171252.6]
  assign _T_907 = ~io_in_b_bits_address[0]; // @[Misc.scala 210:20:freechips.rocketchip.system.DefaultRV32Config.fir@171255.6]
  assign _T_908 = _T_898 & _T_907; // @[Misc.scala 213:27:freechips.rocketchip.system.DefaultRV32Config.fir@171256.6]
  assign _T_909 = _T_894[0] & _T_908; // @[Misc.scala 214:38:freechips.rocketchip.system.DefaultRV32Config.fir@171257.6]
  assign _T_910 = _T_901 | _T_909; // @[Misc.scala 214:29:freechips.rocketchip.system.DefaultRV32Config.fir@171258.6]
  assign _T_911 = _T_898 & io_in_b_bits_address[0]; // @[Misc.scala 213:27:freechips.rocketchip.system.DefaultRV32Config.fir@171259.6]
  assign _T_912 = _T_894[0] & _T_911; // @[Misc.scala 214:38:freechips.rocketchip.system.DefaultRV32Config.fir@171260.6]
  assign _T_913 = _T_901 | _T_912; // @[Misc.scala 214:29:freechips.rocketchip.system.DefaultRV32Config.fir@171261.6]
  assign _T_914 = io_in_b_bits_address[1] & _T_907; // @[Misc.scala 213:27:freechips.rocketchip.system.DefaultRV32Config.fir@171262.6]
  assign _T_915 = _T_894[0] & _T_914; // @[Misc.scala 214:38:freechips.rocketchip.system.DefaultRV32Config.fir@171263.6]
  assign _T_916 = _T_904 | _T_915; // @[Misc.scala 214:29:freechips.rocketchip.system.DefaultRV32Config.fir@171264.6]
  assign _T_917 = io_in_b_bits_address[1] & io_in_b_bits_address[0]; // @[Misc.scala 213:27:freechips.rocketchip.system.DefaultRV32Config.fir@171265.6]
  assign _T_918 = _T_894[0] & _T_917; // @[Misc.scala 214:38:freechips.rocketchip.system.DefaultRV32Config.fir@171266.6]
  assign _T_919 = _T_904 | _T_918; // @[Misc.scala 214:29:freechips.rocketchip.system.DefaultRV32Config.fir@171267.6]
  assign _T_922 = {_T_919,_T_916,_T_913,_T_910}; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@171270.6]
  assign _T_931 = io_in_b_bits_opcode == 3'h6; // @[Monitor.scala 164:25:freechips.rocketchip.system.DefaultRV32Config.fir@171283.6]
  assign _T_935 = 4'h6 == io_in_b_bits_size; // @[Parameters.scala 92:48:freechips.rocketchip.system.DefaultRV32Config.fir@171291.8]
  assign _T_936 = _T_822 & _T_935; // @[Mux.scala 27:72:freechips.rocketchip.system.DefaultRV32Config.fir@171292.8]
  assign _T_941 = _T_936 | reset; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@171298.8]
  assign _T_942 = ~_T_941; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@171299.8]
  assign _T_944 = _T_883 | reset; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@171305.8]
  assign _T_945 = ~_T_944; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@171306.8]
  assign _T_950 = _T_889 | reset; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@171319.8]
  assign _T_951 = ~_T_950; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@171320.8]
  assign _T_952 = io_in_b_bits_param <= 2'h2; // @[Bundles.scala 104:26:freechips.rocketchip.system.DefaultRV32Config.fir@171325.8]
  assign _T_954 = _T_952 | reset; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@171327.8]
  assign _T_955 = ~_T_954; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@171328.8]
  assign _T_956 = io_in_b_bits_mask == _T_922; // @[Monitor.scala 170:30:freechips.rocketchip.system.DefaultRV32Config.fir@171333.8]
  assign _T_958 = _T_956 | reset; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@171335.8]
  assign _T_959 = ~_T_958; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@171336.8]
  assign _T_960 = ~io_in_b_bits_corrupt; // @[Monitor.scala 171:18:freechips.rocketchip.system.DefaultRV32Config.fir@171341.8]
  assign _T_962 = _T_960 | reset; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@171343.8]
  assign _T_963 = ~_T_962; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@171344.8]
  assign _T_964 = io_in_b_bits_opcode == 3'h4; // @[Monitor.scala 174:25:freechips.rocketchip.system.DefaultRV32Config.fir@171350.6]
  assign _T_967 = ~reset; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@171354.8]
  assign _T_977 = io_in_b_bits_param == 2'h0; // @[Monitor.scala 179:31:freechips.rocketchip.system.DefaultRV32Config.fir@171380.8]
  assign _T_979 = _T_977 | reset; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@171382.8]
  assign _T_980 = ~_T_979; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@171383.8]
  assign _T_989 = io_in_b_bits_opcode == 3'h0; // @[Monitor.scala 184:25:freechips.rocketchip.system.DefaultRV32Config.fir@171405.6]
  assign _T_1010 = io_in_b_bits_opcode == 3'h1; // @[Monitor.scala 193:25:freechips.rocketchip.system.DefaultRV32Config.fir@171452.6]
  assign _T_1027 = ~_T_922; // @[Monitor.scala 199:33:freechips.rocketchip.system.DefaultRV32Config.fir@171490.8]
  assign _T_1028 = io_in_b_bits_mask & _T_1027; // @[Monitor.scala 199:31:freechips.rocketchip.system.DefaultRV32Config.fir@171491.8]
  assign _T_1029 = _T_1028 == 4'h0; // @[Monitor.scala 199:40:freechips.rocketchip.system.DefaultRV32Config.fir@171492.8]
  assign _T_1031 = _T_1029 | reset; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@171494.8]
  assign _T_1032 = ~_T_1031; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@171495.8]
  assign _T_1033 = io_in_b_bits_opcode == 3'h2; // @[Monitor.scala 202:25:freechips.rocketchip.system.DefaultRV32Config.fir@171501.6]
  assign _T_1054 = io_in_b_bits_opcode == 3'h3; // @[Monitor.scala 211:25:freechips.rocketchip.system.DefaultRV32Config.fir@171548.6]
  assign _T_1075 = io_in_b_bits_opcode == 3'h5; // @[Monitor.scala 220:25:freechips.rocketchip.system.DefaultRV32Config.fir@171595.6]
  assign _T_1100 = ~io_in_c_bits_source; // @[Parameters.scala 47:9:freechips.rocketchip.system.DefaultRV32Config.fir@171652.6]
  assign _T_1103 = _T_1100 | io_in_c_bits_source; // @[Parameters.scala 924:46:freechips.rocketchip.system.DefaultRV32Config.fir@171658.6]
  assign _T_1105 = 27'hfff << io_in_c_bits_size; // @[package.scala 207:77:freechips.rocketchip.system.DefaultRV32Config.fir@171660.6]
  assign _T_1107 = ~_T_1105[11:0]; // @[package.scala 207:46:freechips.rocketchip.system.DefaultRV32Config.fir@171662.6]
  assign _GEN_73 = {{20'd0}, _T_1107}; // @[Edges.scala 22:16:freechips.rocketchip.system.DefaultRV32Config.fir@171663.6]
  assign _T_1108 = io_in_c_bits_address & _GEN_73; // @[Edges.scala 22:16:freechips.rocketchip.system.DefaultRV32Config.fir@171663.6]
  assign _T_1109 = _T_1108 == 32'h0; // @[Edges.scala 22:24:freechips.rocketchip.system.DefaultRV32Config.fir@171664.6]
  assign _T_1110 = io_in_c_bits_address ^ 32'h3000; // @[Parameters.scala 137:31:freechips.rocketchip.system.DefaultRV32Config.fir@171665.6]
  assign _T_1111 = {1'b0,$signed(_T_1110)}; // @[Parameters.scala 137:49:freechips.rocketchip.system.DefaultRV32Config.fir@171666.6]
  assign _T_1113 = $signed(_T_1111) & -33'sh1000; // @[Parameters.scala 137:52:freechips.rocketchip.system.DefaultRV32Config.fir@171668.6]
  assign _T_1114 = $signed(_T_1113) == 33'sh0; // @[Parameters.scala 137:67:freechips.rocketchip.system.DefaultRV32Config.fir@171669.6]
  assign _T_1115 = io_in_c_bits_address ^ 32'hc000000; // @[Parameters.scala 137:31:freechips.rocketchip.system.DefaultRV32Config.fir@171670.6]
  assign _T_1116 = {1'b0,$signed(_T_1115)}; // @[Parameters.scala 137:49:freechips.rocketchip.system.DefaultRV32Config.fir@171671.6]
  assign _T_1118 = $signed(_T_1116) & -33'sh4000000; // @[Parameters.scala 137:52:freechips.rocketchip.system.DefaultRV32Config.fir@171673.6]
  assign _T_1119 = $signed(_T_1118) == 33'sh0; // @[Parameters.scala 137:67:freechips.rocketchip.system.DefaultRV32Config.fir@171674.6]
  assign _T_1120 = io_in_c_bits_address ^ 32'h2000000; // @[Parameters.scala 137:31:freechips.rocketchip.system.DefaultRV32Config.fir@171675.6]
  assign _T_1121 = {1'b0,$signed(_T_1120)}; // @[Parameters.scala 137:49:freechips.rocketchip.system.DefaultRV32Config.fir@171676.6]
  assign _T_1123 = $signed(_T_1121) & -33'sh10000; // @[Parameters.scala 137:52:freechips.rocketchip.system.DefaultRV32Config.fir@171678.6]
  assign _T_1124 = $signed(_T_1123) == 33'sh0; // @[Parameters.scala 137:67:freechips.rocketchip.system.DefaultRV32Config.fir@171679.6]
  assign _T_1126 = {1'b0,$signed(io_in_c_bits_address)}; // @[Parameters.scala 137:49:freechips.rocketchip.system.DefaultRV32Config.fir@171681.6]
  assign _T_1128 = $signed(_T_1126) & -33'sh1000; // @[Parameters.scala 137:52:freechips.rocketchip.system.DefaultRV32Config.fir@171683.6]
  assign _T_1129 = $signed(_T_1128) == 33'sh0; // @[Parameters.scala 137:67:freechips.rocketchip.system.DefaultRV32Config.fir@171684.6]
  assign _T_1130 = io_in_c_bits_address ^ 32'h10000; // @[Parameters.scala 137:31:freechips.rocketchip.system.DefaultRV32Config.fir@171685.6]
  assign _T_1131 = {1'b0,$signed(_T_1130)}; // @[Parameters.scala 137:49:freechips.rocketchip.system.DefaultRV32Config.fir@171686.6]
  assign _T_1133 = $signed(_T_1131) & -33'sh10000; // @[Parameters.scala 137:52:freechips.rocketchip.system.DefaultRV32Config.fir@171688.6]
  assign _T_1134 = $signed(_T_1133) == 33'sh0; // @[Parameters.scala 137:67:freechips.rocketchip.system.DefaultRV32Config.fir@171689.6]
  assign _T_1135 = io_in_c_bits_address ^ 32'h80000000; // @[Parameters.scala 137:31:freechips.rocketchip.system.DefaultRV32Config.fir@171690.6]
  assign _T_1136 = {1'b0,$signed(_T_1135)}; // @[Parameters.scala 137:49:freechips.rocketchip.system.DefaultRV32Config.fir@171691.6]
  assign _T_1138 = $signed(_T_1136) & -33'sh10000000; // @[Parameters.scala 137:52:freechips.rocketchip.system.DefaultRV32Config.fir@171693.6]
  assign _T_1139 = $signed(_T_1138) == 33'sh0; // @[Parameters.scala 137:67:freechips.rocketchip.system.DefaultRV32Config.fir@171694.6]
  assign _T_1140 = io_in_c_bits_address ^ 32'h60000000; // @[Parameters.scala 137:31:freechips.rocketchip.system.DefaultRV32Config.fir@171695.6]
  assign _T_1141 = {1'b0,$signed(_T_1140)}; // @[Parameters.scala 137:49:freechips.rocketchip.system.DefaultRV32Config.fir@171696.6]
  assign _T_1143 = $signed(_T_1141) & -33'sh20000000; // @[Parameters.scala 137:52:freechips.rocketchip.system.DefaultRV32Config.fir@171698.6]
  assign _T_1144 = $signed(_T_1143) == 33'sh0; // @[Parameters.scala 137:67:freechips.rocketchip.system.DefaultRV32Config.fir@171699.6]
  assign _T_1146 = _T_1114 | _T_1119; // @[Parameters.scala 535:64:freechips.rocketchip.system.DefaultRV32Config.fir@171709.6]
  assign _T_1147 = _T_1146 | _T_1124; // @[Parameters.scala 535:64:freechips.rocketchip.system.DefaultRV32Config.fir@171710.6]
  assign _T_1148 = _T_1147 | _T_1129; // @[Parameters.scala 535:64:freechips.rocketchip.system.DefaultRV32Config.fir@171711.6]
  assign _T_1149 = _T_1148 | _T_1134; // @[Parameters.scala 535:64:freechips.rocketchip.system.DefaultRV32Config.fir@171712.6]
  assign _T_1150 = _T_1149 | _T_1139; // @[Parameters.scala 535:64:freechips.rocketchip.system.DefaultRV32Config.fir@171713.6]
  assign _T_1151 = _T_1150 | _T_1144; // @[Parameters.scala 535:64:freechips.rocketchip.system.DefaultRV32Config.fir@171714.6]
  assign _T_1172 = io_in_c_bits_opcode == 3'h4; // @[Monitor.scala 239:25:freechips.rocketchip.system.DefaultRV32Config.fir@171739.6]
  assign _T_1174 = _T_1151 | reset; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@171742.8]
  assign _T_1175 = ~_T_1174; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@171743.8]
  assign _T_1177 = _T_1103 | reset; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@171749.8]
  assign _T_1178 = ~_T_1177; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@171750.8]
  assign _T_1179 = io_in_c_bits_size >= 4'h2; // @[Monitor.scala 242:30:freechips.rocketchip.system.DefaultRV32Config.fir@171755.8]
  assign _T_1181 = _T_1179 | reset; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@171757.8]
  assign _T_1182 = ~_T_1181; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@171758.8]
  assign _T_1184 = _T_1109 | reset; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@171764.8]
  assign _T_1185 = ~_T_1184; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@171765.8]
  assign _T_1186 = io_in_c_bits_param <= 3'h5; // @[Bundles.scala 122:29:freechips.rocketchip.system.DefaultRV32Config.fir@171770.8]
  assign _T_1188 = _T_1186 | reset; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@171772.8]
  assign _T_1189 = ~_T_1188; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@171773.8]
  assign _T_1194 = io_in_c_bits_opcode == 3'h5; // @[Monitor.scala 248:25:freechips.rocketchip.system.DefaultRV32Config.fir@171787.6]
  assign _T_1212 = io_in_c_bits_opcode == 3'h6; // @[Monitor.scala 256:25:freechips.rocketchip.system.DefaultRV32Config.fir@171827.6]
  assign _T_1251 = io_in_c_bits_size <= 4'h6; // @[Parameters.scala 93:42:freechips.rocketchip.system.DefaultRV32Config.fir@171867.8]
  assign _T_1259 = _T_1251 & _T_1139; // @[Parameters.scala 551:56:freechips.rocketchip.system.DefaultRV32Config.fir@171875.8]
  assign _T_1263 = _T_1259 | reset; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@171879.8]
  assign _T_1264 = ~_T_1263; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@171880.8]
  assign _T_1268 = 4'h6 == io_in_c_bits_size; // @[Parameters.scala 92:48:freechips.rocketchip.system.DefaultRV32Config.fir@171891.8]
  assign _T_1269 = _T_1100 & _T_1268; // @[Mux.scala 27:72:freechips.rocketchip.system.DefaultRV32Config.fir@171892.8]
  assign _T_1274 = _T_1269 | reset; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@171898.8]
  assign _T_1275 = ~_T_1274; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@171899.8]
  assign _T_1286 = io_in_c_bits_param <= 3'h2; // @[Bundles.scala 116:29:freechips.rocketchip.system.DefaultRV32Config.fir@171926.8]
  assign _T_1288 = _T_1286 | reset; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@171928.8]
  assign _T_1289 = ~_T_1288; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@171929.8]
  assign _T_1294 = io_in_c_bits_opcode == 3'h7; // @[Monitor.scala 266:25:freechips.rocketchip.system.DefaultRV32Config.fir@171943.6]
  assign _T_1372 = io_in_c_bits_opcode == 3'h0; // @[Monitor.scala 275:25:freechips.rocketchip.system.DefaultRV32Config.fir@172051.6]
  assign _T_1382 = io_in_c_bits_param == 3'h0; // @[Monitor.scala 279:31:freechips.rocketchip.system.DefaultRV32Config.fir@172074.8]
  assign _T_1384 = _T_1382 | reset; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@172076.8]
  assign _T_1385 = ~_T_1384; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@172077.8]
  assign _T_1390 = io_in_c_bits_opcode == 3'h1; // @[Monitor.scala 283:25:freechips.rocketchip.system.DefaultRV32Config.fir@172091.6]
  assign _T_1404 = io_in_c_bits_opcode == 3'h2; // @[Monitor.scala 290:25:freechips.rocketchip.system.DefaultRV32Config.fir@172123.6]
  assign _T_1426 = io_in_a_ready & io_in_a_valid; // @[Decoupled.scala 40:37:freechips.rocketchip.system.DefaultRV32Config.fir@172174.4]
  assign _T_1433 = ~io_in_a_bits_opcode[2]; // @[Edges.scala 93:28:freechips.rocketchip.system.DefaultRV32Config.fir@172181.4]
  assign _T_1437 = _T_1435 - 10'h1; // @[Edges.scala 231:28:freechips.rocketchip.system.DefaultRV32Config.fir@172185.4]
  assign _T_1438 = _T_1435 == 10'h0; // @[Edges.scala 232:25:freechips.rocketchip.system.DefaultRV32Config.fir@172186.4]
  assign _T_1451 = ~_T_1438; // @[Monitor.scala 386:22:freechips.rocketchip.system.DefaultRV32Config.fir@172202.4]
  assign _T_1452 = io_in_a_valid & _T_1451; // @[Monitor.scala 386:19:freechips.rocketchip.system.DefaultRV32Config.fir@172203.4]
  assign _T_1453 = io_in_a_bits_opcode == _T_1446; // @[Monitor.scala 387:32:freechips.rocketchip.system.DefaultRV32Config.fir@172205.6]
  assign _T_1455 = _T_1453 | reset; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@172207.6]
  assign _T_1456 = ~_T_1455; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@172208.6]
  assign _T_1457 = io_in_a_bits_param == _T_1447; // @[Monitor.scala 388:32:freechips.rocketchip.system.DefaultRV32Config.fir@172213.6]
  assign _T_1459 = _T_1457 | reset; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@172215.6]
  assign _T_1460 = ~_T_1459; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@172216.6]
  assign _T_1461 = io_in_a_bits_size == _T_1448; // @[Monitor.scala 389:32:freechips.rocketchip.system.DefaultRV32Config.fir@172221.6]
  assign _T_1463 = _T_1461 | reset; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@172223.6]
  assign _T_1464 = ~_T_1463; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@172224.6]
  assign _T_1465 = io_in_a_bits_source == _T_1449; // @[Monitor.scala 390:32:freechips.rocketchip.system.DefaultRV32Config.fir@172229.6]
  assign _T_1467 = _T_1465 | reset; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@172231.6]
  assign _T_1468 = ~_T_1467; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@172232.6]
  assign _T_1469 = io_in_a_bits_address == _T_1450; // @[Monitor.scala 391:32:freechips.rocketchip.system.DefaultRV32Config.fir@172237.6]
  assign _T_1471 = _T_1469 | reset; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@172239.6]
  assign _T_1472 = ~_T_1471; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@172240.6]
  assign _T_1474 = _T_1426 & _T_1438; // @[Monitor.scala 393:20:freechips.rocketchip.system.DefaultRV32Config.fir@172247.4]
  assign _T_1475 = io_in_d_ready & io_in_d_valid; // @[Decoupled.scala 40:37:freechips.rocketchip.system.DefaultRV32Config.fir@172255.4]
  assign _T_1477 = 27'hfff << io_in_d_bits_size; // @[package.scala 207:77:freechips.rocketchip.system.DefaultRV32Config.fir@172257.4]
  assign _T_1479 = ~_T_1477[11:0]; // @[package.scala 207:46:freechips.rocketchip.system.DefaultRV32Config.fir@172259.4]
  assign _T_1485 = _T_1483 - 10'h1; // @[Edges.scala 231:28:freechips.rocketchip.system.DefaultRV32Config.fir@172265.4]
  assign _T_1486 = _T_1483 == 10'h0; // @[Edges.scala 232:25:freechips.rocketchip.system.DefaultRV32Config.fir@172266.4]
  assign _T_1500 = ~_T_1486; // @[Monitor.scala 538:22:freechips.rocketchip.system.DefaultRV32Config.fir@172283.4]
  assign _T_1501 = io_in_d_valid & _T_1500; // @[Monitor.scala 538:19:freechips.rocketchip.system.DefaultRV32Config.fir@172284.4]
  assign _T_1502 = io_in_d_bits_opcode == _T_1494; // @[Monitor.scala 539:29:freechips.rocketchip.system.DefaultRV32Config.fir@172286.6]
  assign _T_1504 = _T_1502 | reset; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@172288.6]
  assign _T_1505 = ~_T_1504; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@172289.6]
  assign _T_1506 = io_in_d_bits_param == _T_1495; // @[Monitor.scala 540:29:freechips.rocketchip.system.DefaultRV32Config.fir@172294.6]
  assign _T_1508 = _T_1506 | reset; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@172296.6]
  assign _T_1509 = ~_T_1508; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@172297.6]
  assign _T_1510 = io_in_d_bits_size == _T_1496; // @[Monitor.scala 541:29:freechips.rocketchip.system.DefaultRV32Config.fir@172302.6]
  assign _T_1512 = _T_1510 | reset; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@172304.6]
  assign _T_1513 = ~_T_1512; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@172305.6]
  assign _T_1514 = io_in_d_bits_source == _T_1497; // @[Monitor.scala 542:29:freechips.rocketchip.system.DefaultRV32Config.fir@172310.6]
  assign _T_1516 = _T_1514 | reset; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@172312.6]
  assign _T_1517 = ~_T_1516; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@172313.6]
  assign _T_1518 = io_in_d_bits_sink == _T_1498; // @[Monitor.scala 543:29:freechips.rocketchip.system.DefaultRV32Config.fir@172318.6]
  assign _T_1520 = _T_1518 | reset; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@172320.6]
  assign _T_1521 = ~_T_1520; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@172321.6]
  assign _T_1522 = io_in_d_bits_denied == _T_1499; // @[Monitor.scala 544:29:freechips.rocketchip.system.DefaultRV32Config.fir@172326.6]
  assign _T_1524 = _T_1522 | reset; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@172328.6]
  assign _T_1525 = ~_T_1524; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@172329.6]
  assign _T_1527 = _T_1475 & _T_1486; // @[Monitor.scala 546:20:freechips.rocketchip.system.DefaultRV32Config.fir@172336.4]
  assign _T_1528 = io_in_b_ready & io_in_b_valid; // @[Decoupled.scala 40:37:freechips.rocketchip.system.DefaultRV32Config.fir@172345.4]
  assign _T_1539 = _T_1537 - 10'h1; // @[Edges.scala 231:28:freechips.rocketchip.system.DefaultRV32Config.fir@172356.4]
  assign _T_1540 = _T_1537 == 10'h0; // @[Edges.scala 232:25:freechips.rocketchip.system.DefaultRV32Config.fir@172357.4]
  assign _T_1553 = ~_T_1540; // @[Monitor.scala 409:22:freechips.rocketchip.system.DefaultRV32Config.fir@172373.4]
  assign _T_1554 = io_in_b_valid & _T_1553; // @[Monitor.scala 409:19:freechips.rocketchip.system.DefaultRV32Config.fir@172374.4]
  assign _T_1555 = io_in_b_bits_opcode == _T_1548; // @[Monitor.scala 410:32:freechips.rocketchip.system.DefaultRV32Config.fir@172376.6]
  assign _T_1557 = _T_1555 | reset; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@172378.6]
  assign _T_1558 = ~_T_1557; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@172379.6]
  assign _T_1559 = io_in_b_bits_param == _T_1549; // @[Monitor.scala 411:32:freechips.rocketchip.system.DefaultRV32Config.fir@172384.6]
  assign _T_1561 = _T_1559 | reset; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@172386.6]
  assign _T_1562 = ~_T_1561; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@172387.6]
  assign _T_1563 = io_in_b_bits_size == _T_1550; // @[Monitor.scala 412:32:freechips.rocketchip.system.DefaultRV32Config.fir@172392.6]
  assign _T_1565 = _T_1563 | reset; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@172394.6]
  assign _T_1566 = ~_T_1565; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@172395.6]
  assign _T_1567 = io_in_b_bits_source == _T_1551; // @[Monitor.scala 413:32:freechips.rocketchip.system.DefaultRV32Config.fir@172400.6]
  assign _T_1569 = _T_1567 | reset; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@172402.6]
  assign _T_1570 = ~_T_1569; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@172403.6]
  assign _T_1571 = io_in_b_bits_address == _T_1552; // @[Monitor.scala 414:32:freechips.rocketchip.system.DefaultRV32Config.fir@172408.6]
  assign _T_1573 = _T_1571 | reset; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@172410.6]
  assign _T_1574 = ~_T_1573; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@172411.6]
  assign _T_1576 = _T_1528 & _T_1540; // @[Monitor.scala 416:20:freechips.rocketchip.system.DefaultRV32Config.fir@172418.4]
  assign _T_1577 = io_in_c_ready & io_in_c_valid; // @[Decoupled.scala 40:37:freechips.rocketchip.system.DefaultRV32Config.fir@172426.4]
  assign _T_1587 = _T_1585 - 10'h1; // @[Edges.scala 231:28:freechips.rocketchip.system.DefaultRV32Config.fir@172436.4]
  assign _T_1588 = _T_1585 == 10'h0; // @[Edges.scala 232:25:freechips.rocketchip.system.DefaultRV32Config.fir@172437.4]
  assign _T_1601 = ~_T_1588; // @[Monitor.scala 514:22:freechips.rocketchip.system.DefaultRV32Config.fir@172453.4]
  assign _T_1602 = io_in_c_valid & _T_1601; // @[Monitor.scala 514:19:freechips.rocketchip.system.DefaultRV32Config.fir@172454.4]
  assign _T_1603 = io_in_c_bits_opcode == _T_1596; // @[Monitor.scala 515:32:freechips.rocketchip.system.DefaultRV32Config.fir@172456.6]
  assign _T_1605 = _T_1603 | reset; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@172458.6]
  assign _T_1606 = ~_T_1605; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@172459.6]
  assign _T_1607 = io_in_c_bits_param == _T_1597; // @[Monitor.scala 516:32:freechips.rocketchip.system.DefaultRV32Config.fir@172464.6]
  assign _T_1609 = _T_1607 | reset; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@172466.6]
  assign _T_1610 = ~_T_1609; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@172467.6]
  assign _T_1611 = io_in_c_bits_size == _T_1598; // @[Monitor.scala 517:32:freechips.rocketchip.system.DefaultRV32Config.fir@172472.6]
  assign _T_1613 = _T_1611 | reset; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@172474.6]
  assign _T_1614 = ~_T_1613; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@172475.6]
  assign _T_1615 = io_in_c_bits_source == _T_1599; // @[Monitor.scala 518:32:freechips.rocketchip.system.DefaultRV32Config.fir@172480.6]
  assign _T_1617 = _T_1615 | reset; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@172482.6]
  assign _T_1618 = ~_T_1617; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@172483.6]
  assign _T_1619 = io_in_c_bits_address == _T_1600; // @[Monitor.scala 519:32:freechips.rocketchip.system.DefaultRV32Config.fir@172488.6]
  assign _T_1621 = _T_1619 | reset; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@172490.6]
  assign _T_1622 = ~_T_1621; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@172491.6]
  assign _T_1624 = _T_1577 & _T_1588; // @[Monitor.scala 521:20:freechips.rocketchip.system.DefaultRV32Config.fir@172498.4]
  assign _T_1636 = _T_1634 - 10'h1; // @[Edges.scala 231:28:freechips.rocketchip.system.DefaultRV32Config.fir@172520.4]
  assign a_first = _T_1634 == 10'h0; // @[Edges.scala 232:25:freechips.rocketchip.system.DefaultRV32Config.fir@172521.4]
  assign _T_1654 = _T_1652 - 10'h1; // @[Edges.scala 231:28:freechips.rocketchip.system.DefaultRV32Config.fir@172542.4]
  assign d_first = _T_1652 == 10'h0; // @[Edges.scala 232:25:freechips.rocketchip.system.DefaultRV32Config.fir@172543.4]
  assign _GEN_74 = {io_in_d_bits_source, 2'h0}; // @[Monitor.scala 629:69:freechips.rocketchip.system.DefaultRV32Config.fir@172562.4]
  assign _T_1662 = {{1'd0}, _GEN_74}; // @[Monitor.scala 629:69:freechips.rocketchip.system.DefaultRV32Config.fir@172562.4]
  assign _T_1663 = inflight_opcodes >> _T_1662; // @[Monitor.scala 629:44:freechips.rocketchip.system.DefaultRV32Config.fir@172563.4]
  assign _T_1667 = 16'h10 - 16'h1; // @[Monitor.scala 606:57:freechips.rocketchip.system.DefaultRV32Config.fir@172567.4]
  assign _GEN_75 = {{8'd0}, _T_1663}; // @[Monitor.scala 629:97:freechips.rocketchip.system.DefaultRV32Config.fir@172568.4]
  assign _T_1668 = _GEN_75 & _T_1667; // @[Monitor.scala 629:97:freechips.rocketchip.system.DefaultRV32Config.fir@172568.4]
  assign _T_1669 = {{1'd0}, _T_1668[15:1]}; // @[Monitor.scala 629:152:freechips.rocketchip.system.DefaultRV32Config.fir@172569.4]
  assign _T_1670 = {io_in_d_bits_source, 3'h0}; // @[Monitor.scala 633:65:freechips.rocketchip.system.DefaultRV32Config.fir@172573.4]
  assign _T_1671 = inflight_sizes >> _T_1670; // @[Monitor.scala 633:40:freechips.rocketchip.system.DefaultRV32Config.fir@172574.4]
  assign _T_1675 = 16'h100 - 16'h1; // @[Monitor.scala 606:57:freechips.rocketchip.system.DefaultRV32Config.fir@172578.4]
  assign _T_1676 = _T_1671 & _T_1675; // @[Monitor.scala 633:91:freechips.rocketchip.system.DefaultRV32Config.fir@172579.4]
  assign _T_1677 = {{1'd0}, _T_1676[15:1]}; // @[Monitor.scala 633:144:freechips.rocketchip.system.DefaultRV32Config.fir@172580.4]
  assign _T_1681 = _T_1426 & a_first; // @[Monitor.scala 643:27:freechips.rocketchip.system.DefaultRV32Config.fir@172605.4]
  assign _T_1683 = 2'h1 << io_in_a_bits_source; // @[OneHot.scala 58:35:freechips.rocketchip.system.DefaultRV32Config.fir@172608.6]
  assign _T_1684 = {io_in_a_bits_opcode, 1'h0}; // @[Monitor.scala 645:53:freechips.rocketchip.system.DefaultRV32Config.fir@172610.6]
  assign _T_1685 = _T_1684 | 4'h1; // @[Monitor.scala 645:61:freechips.rocketchip.system.DefaultRV32Config.fir@172611.6]
  assign _T_1686 = {io_in_a_bits_size, 1'h0}; // @[Monitor.scala 646:49:freechips.rocketchip.system.DefaultRV32Config.fir@172613.6]
  assign _T_1687 = _T_1686 | 5'h1; // @[Monitor.scala 646:57:freechips.rocketchip.system.DefaultRV32Config.fir@172614.6]
  assign _GEN_78 = {io_in_a_bits_source, 2'h0}; // @[Monitor.scala 647:72:freechips.rocketchip.system.DefaultRV32Config.fir@172616.6]
  assign _T_1688 = {{1'd0}, _GEN_78}; // @[Monitor.scala 647:72:freechips.rocketchip.system.DefaultRV32Config.fir@172616.6]
  assign a_opcodes_set_interm = _T_1681 ? _T_1685 : 4'h0; // @[Monitor.scala 643:72:freechips.rocketchip.system.DefaultRV32Config.fir@172607.4]
  assign _GEN_79 = {{15'd0}, a_opcodes_set_interm}; // @[Monitor.scala 647:47:freechips.rocketchip.system.DefaultRV32Config.fir@172617.6]
  assign _T_1689 = _GEN_79 << _T_1688; // @[Monitor.scala 647:47:freechips.rocketchip.system.DefaultRV32Config.fir@172617.6]
  assign _T_1690 = {io_in_a_bits_source, 3'h0}; // @[Monitor.scala 648:68:freechips.rocketchip.system.DefaultRV32Config.fir@172619.6]
  assign a_sizes_set_interm = _T_1681 ? _T_1687 : 5'h0; // @[Monitor.scala 643:72:freechips.rocketchip.system.DefaultRV32Config.fir@172607.4]
  assign _GEN_80 = {{15'd0}, a_sizes_set_interm}; // @[Monitor.scala 648:43:freechips.rocketchip.system.DefaultRV32Config.fir@172620.6]
  assign _T_1691 = _GEN_80 << _T_1690; // @[Monitor.scala 648:43:freechips.rocketchip.system.DefaultRV32Config.fir@172620.6]
  assign _T_1692 = inflight >> io_in_a_bits_source; // @[Monitor.scala 649:26:freechips.rocketchip.system.DefaultRV32Config.fir@172622.6]
  assign _T_1694 = ~_T_1692[0]; // @[Monitor.scala 649:17:freechips.rocketchip.system.DefaultRV32Config.fir@172624.6]
  assign _T_1696 = _T_1694 | reset; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@172626.6]
  assign _T_1697 = ~_T_1696; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@172627.6]
  assign a_set = _T_1681 ? _T_1683 : 2'h0; // @[Monitor.scala 643:72:freechips.rocketchip.system.DefaultRV32Config.fir@172607.4]
  assign _GEN_30 = _T_1681 ? _T_1689 : 19'h0; // @[Monitor.scala 643:72:freechips.rocketchip.system.DefaultRV32Config.fir@172607.4]
  assign _GEN_31 = _T_1681 ? _T_1691 : 20'h0; // @[Monitor.scala 643:72:freechips.rocketchip.system.DefaultRV32Config.fir@172607.4]
  assign _T_1700 = _T_1475 & d_first; // @[Monitor.scala 660:27:freechips.rocketchip.system.DefaultRV32Config.fir@172641.4]
  assign _T_1702 = ~_T_689; // @[Monitor.scala 660:75:freechips.rocketchip.system.DefaultRV32Config.fir@172643.4]
  assign _T_1703 = _T_1700 & _T_1702; // @[Monitor.scala 660:72:freechips.rocketchip.system.DefaultRV32Config.fir@172644.4]
  assign _T_1704 = 2'h1 << io_in_d_bits_source; // @[OneHot.scala 58:35:freechips.rocketchip.system.DefaultRV32Config.fir@172646.6]
  assign _GEN_82 = {{15'd0}, _T_1667}; // @[Monitor.scala 662:76:freechips.rocketchip.system.DefaultRV32Config.fir@172653.6]
  assign _T_1710 = _GEN_82 << _T_1662; // @[Monitor.scala 662:76:freechips.rocketchip.system.DefaultRV32Config.fir@172653.6]
  assign _GEN_83 = {{15'd0}, _T_1675}; // @[Monitor.scala 663:72:freechips.rocketchip.system.DefaultRV32Config.fir@172660.6]
  assign _T_1716 = _GEN_83 << _T_1670; // @[Monitor.scala 663:72:freechips.rocketchip.system.DefaultRV32Config.fir@172660.6]
  assign d_clr = _T_1703 ? _T_1704 : 2'h0; // @[Monitor.scala 660:91:freechips.rocketchip.system.DefaultRV32Config.fir@172645.4]
  assign _GEN_33 = _T_1703 ? _T_1710 : 31'h0; // @[Monitor.scala 660:91:freechips.rocketchip.system.DefaultRV32Config.fir@172645.4]
  assign _GEN_34 = _T_1703 ? _T_1716 : 31'h0; // @[Monitor.scala 660:91:freechips.rocketchip.system.DefaultRV32Config.fir@172645.4]
  assign _T_1717 = io_in_d_valid & d_first; // @[Monitor.scala 665:26:freechips.rocketchip.system.DefaultRV32Config.fir@172663.4]
  assign _T_1720 = _T_1717 & _T_1702; // @[Monitor.scala 665:71:freechips.rocketchip.system.DefaultRV32Config.fir@172666.4]
  assign _T_1721 = inflight >> io_in_d_bits_source; // @[Monitor.scala 666:25:freechips.rocketchip.system.DefaultRV32Config.fir@172668.6]
  assign _T_1723 = io_in_a_bits_source == io_in_d_bits_source; // @[Monitor.scala 666:93:freechips.rocketchip.system.DefaultRV32Config.fir@172670.6]
  assign _T_1724 = io_in_a_valid & _T_1723; // @[Monitor.scala 666:68:freechips.rocketchip.system.DefaultRV32Config.fir@172671.6]
  assign _T_1725 = io_in_a_bits_size == io_in_d_bits_size; // @[Monitor.scala 666:142:freechips.rocketchip.system.DefaultRV32Config.fir@172672.6]
  assign _T_1726 = _T_1724 & _T_1725; // @[Monitor.scala 666:119:freechips.rocketchip.system.DefaultRV32Config.fir@172673.6]
  assign _T_1727 = _T_1726 & a_first; // @[Monitor.scala 666:166:freechips.rocketchip.system.DefaultRV32Config.fir@172674.6]
  assign _T_1728 = _T_1721[0] | _T_1727; // @[Monitor.scala 666:49:freechips.rocketchip.system.DefaultRV32Config.fir@172675.6]
  assign _T_1730 = _T_1728 | reset; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@172677.6]
  assign _T_1731 = ~_T_1730; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@172678.6]
  assign a_opcode_lookup = _T_1669[3:0]; // @[:freechips.rocketchip.system.DefaultRV32Config.fir@172560.4 :freechips.rocketchip.system.DefaultRV32Config.fir@172561.4 Monitor.scala 629:21:freechips.rocketchip.system.DefaultRV32Config.fir@172570.4]
  assign _GEN_37 = 3'h2 == a_opcode_lookup[2:0] ? 3'h1 : 3'h0; // @[Monitor.scala 667:37:freechips.rocketchip.system.DefaultRV32Config.fir@172684.6]
  assign _GEN_38 = 3'h3 == a_opcode_lookup[2:0] ? 3'h1 : _GEN_37; // @[Monitor.scala 667:37:freechips.rocketchip.system.DefaultRV32Config.fir@172684.6]
  assign _GEN_39 = 3'h4 == a_opcode_lookup[2:0] ? 3'h1 : _GEN_38; // @[Monitor.scala 667:37:freechips.rocketchip.system.DefaultRV32Config.fir@172684.6]
  assign _GEN_40 = 3'h5 == a_opcode_lookup[2:0] ? 3'h2 : _GEN_39; // @[Monitor.scala 667:37:freechips.rocketchip.system.DefaultRV32Config.fir@172684.6]
  assign _GEN_41 = 3'h6 == a_opcode_lookup[2:0] ? 3'h4 : _GEN_40; // @[Monitor.scala 667:37:freechips.rocketchip.system.DefaultRV32Config.fir@172684.6]
  assign _GEN_42 = 3'h7 == a_opcode_lookup[2:0] ? 3'h4 : _GEN_41; // @[Monitor.scala 667:37:freechips.rocketchip.system.DefaultRV32Config.fir@172684.6]
  assign _T_1733 = io_in_d_bits_opcode == _GEN_42; // @[Monitor.scala 667:37:freechips.rocketchip.system.DefaultRV32Config.fir@172684.6]
  assign _GEN_49 = 3'h6 == a_opcode_lookup[2:0] ? 3'h5 : _GEN_40; // @[Monitor.scala 667:96:freechips.rocketchip.system.DefaultRV32Config.fir@172686.6]
  assign _GEN_50 = 3'h7 == a_opcode_lookup[2:0] ? 3'h4 : _GEN_49; // @[Monitor.scala 667:96:freechips.rocketchip.system.DefaultRV32Config.fir@172686.6]
  assign _T_1735 = io_in_d_bits_opcode == _GEN_50; // @[Monitor.scala 667:96:freechips.rocketchip.system.DefaultRV32Config.fir@172686.6]
  assign _T_1736 = _T_1733 | _T_1735; // @[Monitor.scala 667:71:freechips.rocketchip.system.DefaultRV32Config.fir@172687.6]
  assign _GEN_53 = 3'h2 == io_in_a_bits_opcode ? 3'h1 : 3'h0; // @[Monitor.scala 668:60:freechips.rocketchip.system.DefaultRV32Config.fir@172688.6]
  assign _GEN_54 = 3'h3 == io_in_a_bits_opcode ? 3'h1 : _GEN_53; // @[Monitor.scala 668:60:freechips.rocketchip.system.DefaultRV32Config.fir@172688.6]
  assign _GEN_55 = 3'h4 == io_in_a_bits_opcode ? 3'h1 : _GEN_54; // @[Monitor.scala 668:60:freechips.rocketchip.system.DefaultRV32Config.fir@172688.6]
  assign _GEN_56 = 3'h5 == io_in_a_bits_opcode ? 3'h2 : _GEN_55; // @[Monitor.scala 668:60:freechips.rocketchip.system.DefaultRV32Config.fir@172688.6]
  assign _GEN_57 = 3'h6 == io_in_a_bits_opcode ? 3'h4 : _GEN_56; // @[Monitor.scala 668:60:freechips.rocketchip.system.DefaultRV32Config.fir@172688.6]
  assign _GEN_58 = 3'h7 == io_in_a_bits_opcode ? 3'h4 : _GEN_57; // @[Monitor.scala 668:60:freechips.rocketchip.system.DefaultRV32Config.fir@172688.6]
  assign _T_1737 = io_in_d_bits_opcode == _GEN_58; // @[Monitor.scala 668:60:freechips.rocketchip.system.DefaultRV32Config.fir@172688.6]
  assign _GEN_65 = 3'h6 == io_in_a_bits_opcode ? 3'h5 : _GEN_56; // @[Monitor.scala 668:124:freechips.rocketchip.system.DefaultRV32Config.fir@172689.6]
  assign _GEN_66 = 3'h7 == io_in_a_bits_opcode ? 3'h4 : _GEN_65; // @[Monitor.scala 668:124:freechips.rocketchip.system.DefaultRV32Config.fir@172689.6]
  assign _T_1738 = io_in_d_bits_opcode == _GEN_66; // @[Monitor.scala 668:124:freechips.rocketchip.system.DefaultRV32Config.fir@172689.6]
  assign _T_1739 = _T_1737 | _T_1738; // @[Monitor.scala 668:99:freechips.rocketchip.system.DefaultRV32Config.fir@172690.6]
  assign _T_1740 = io_in_a_valid & _T_1739; // @[Monitor.scala 668:34:freechips.rocketchip.system.DefaultRV32Config.fir@172691.6]
  assign _T_1741 = _T_1736 | _T_1740; // @[Monitor.scala 668:15:freechips.rocketchip.system.DefaultRV32Config.fir@172692.6]
  assign _T_1743 = _T_1741 | reset; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@172694.6]
  assign _T_1744 = ~_T_1743; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@172695.6]
  assign a_size_lookup = _T_1677[7:0]; // @[:freechips.rocketchip.system.DefaultRV32Config.fir@172571.4 :freechips.rocketchip.system.DefaultRV32Config.fir@172572.4 Monitor.scala 633:19:freechips.rocketchip.system.DefaultRV32Config.fir@172581.4]
  assign _GEN_84 = {{4'd0}, io_in_d_bits_size}; // @[Monitor.scala 670:34:freechips.rocketchip.system.DefaultRV32Config.fir@172700.6]
  assign _T_1745 = _GEN_84 == a_size_lookup; // @[Monitor.scala 670:34:freechips.rocketchip.system.DefaultRV32Config.fir@172700.6]
  assign _T_1747 = io_in_a_valid & _T_1725; // @[Monitor.scala 670:72:freechips.rocketchip.system.DefaultRV32Config.fir@172702.6]
  assign _T_1748 = _T_1745 | _T_1747; // @[Monitor.scala 670:53:freechips.rocketchip.system.DefaultRV32Config.fir@172703.6]
  assign _T_1750 = _T_1748 | reset; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@172705.6]
  assign _T_1751 = ~_T_1750; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@172706.6]
  assign _T_1753 = _T_1717 & a_first; // @[Monitor.scala 672:36:freechips.rocketchip.system.DefaultRV32Config.fir@172713.4]
  assign _T_1754 = _T_1753 & io_in_a_valid; // @[Monitor.scala 672:47:freechips.rocketchip.system.DefaultRV32Config.fir@172714.4]
  assign _T_1756 = _T_1754 & _T_1723; // @[Monitor.scala 672:65:freechips.rocketchip.system.DefaultRV32Config.fir@172716.4]
  assign _T_1758 = _T_1756 & _T_1702; // @[Monitor.scala 672:116:freechips.rocketchip.system.DefaultRV32Config.fir@172718.4]
  assign _T_1759 = ~io_in_d_ready; // @[Monitor.scala 673:15:freechips.rocketchip.system.DefaultRV32Config.fir@172720.6]
  assign _T_1760 = _T_1759 | io_in_a_ready; // @[Monitor.scala 673:32:freechips.rocketchip.system.DefaultRV32Config.fir@172721.6]
  assign _T_1762 = _T_1760 | reset; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@172723.6]
  assign _T_1763 = ~_T_1762; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@172724.6]
  assign _T_1764 = a_set != d_clr; // @[Monitor.scala 677:20:freechips.rocketchip.system.DefaultRV32Config.fir@172730.4]
  assign _T_1765 = |a_set; // @[Monitor.scala 677:40:freechips.rocketchip.system.DefaultRV32Config.fir@172731.4]
  assign _T_1766 = ~_T_1765; // @[Monitor.scala 677:33:freechips.rocketchip.system.DefaultRV32Config.fir@172732.4]
  assign _T_1767 = _T_1764 | _T_1766; // @[Monitor.scala 677:30:freechips.rocketchip.system.DefaultRV32Config.fir@172733.4]
  assign _T_1769 = _T_1767 | reset; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@172735.4]
  assign _T_1770 = ~_T_1769; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@172736.4]
  assign _T_1771 = inflight | a_set; // @[Monitor.scala 680:27:freechips.rocketchip.system.DefaultRV32Config.fir@172741.4]
  assign _T_1772 = ~d_clr; // @[Monitor.scala 680:38:freechips.rocketchip.system.DefaultRV32Config.fir@172742.4]
  assign _T_1773 = _T_1771 & _T_1772; // @[Monitor.scala 680:36:freechips.rocketchip.system.DefaultRV32Config.fir@172743.4]
  assign a_opcodes_set = _GEN_30[7:0]; // @[:freechips.rocketchip.system.DefaultRV32Config.fir@172556.4 :freechips.rocketchip.system.DefaultRV32Config.fir@172557.4 Monitor.scala 647:21:freechips.rocketchip.system.DefaultRV32Config.fir@172618.6]
  assign _T_1774 = inflight_opcodes | a_opcodes_set; // @[Monitor.scala 681:43:freechips.rocketchip.system.DefaultRV32Config.fir@172745.4]
  assign d_opcodes_clr = _GEN_33[7:0]; // @[:freechips.rocketchip.system.DefaultRV32Config.fir@172635.4 :freechips.rocketchip.system.DefaultRV32Config.fir@172636.4 Monitor.scala 662:21:freechips.rocketchip.system.DefaultRV32Config.fir@172654.6]
  assign _T_1775 = ~d_opcodes_clr; // @[Monitor.scala 681:62:freechips.rocketchip.system.DefaultRV32Config.fir@172746.4]
  assign _T_1776 = _T_1774 & _T_1775; // @[Monitor.scala 681:60:freechips.rocketchip.system.DefaultRV32Config.fir@172747.4]
  assign a_sizes_set = _GEN_31[15:0]; // @[:freechips.rocketchip.system.DefaultRV32Config.fir@172558.4 :freechips.rocketchip.system.DefaultRV32Config.fir@172559.4 Monitor.scala 648:19:freechips.rocketchip.system.DefaultRV32Config.fir@172621.6]
  assign _T_1777 = inflight_sizes | a_sizes_set; // @[Monitor.scala 682:39:freechips.rocketchip.system.DefaultRV32Config.fir@172749.4]
  assign d_sizes_clr = _GEN_34[15:0]; // @[:freechips.rocketchip.system.DefaultRV32Config.fir@172637.4 :freechips.rocketchip.system.DefaultRV32Config.fir@172638.4 Monitor.scala 663:19:freechips.rocketchip.system.DefaultRV32Config.fir@172661.6]
  assign _T_1778 = ~d_sizes_clr; // @[Monitor.scala 682:56:freechips.rocketchip.system.DefaultRV32Config.fir@172750.4]
  assign _T_1779 = _T_1777 & _T_1778; // @[Monitor.scala 682:54:freechips.rocketchip.system.DefaultRV32Config.fir@172751.4]
  assign _T_1781 = |inflight; // @[Monitor.scala 687:26:freechips.rocketchip.system.DefaultRV32Config.fir@172756.4]
  assign _T_1782 = ~_T_1781; // @[Monitor.scala 687:16:freechips.rocketchip.system.DefaultRV32Config.fir@172757.4]
  assign _T_1783 = plusarg_reader_out == 32'h0; // @[Monitor.scala 687:39:freechips.rocketchip.system.DefaultRV32Config.fir@172758.4]
  assign _T_1784 = _T_1782 | _T_1783; // @[Monitor.scala 687:30:freechips.rocketchip.system.DefaultRV32Config.fir@172759.4]
  assign _T_1785 = _T_1780 < plusarg_reader_out; // @[Monitor.scala 687:59:freechips.rocketchip.system.DefaultRV32Config.fir@172760.4]
  assign _T_1786 = _T_1784 | _T_1785; // @[Monitor.scala 687:47:freechips.rocketchip.system.DefaultRV32Config.fir@172761.4]
  assign _T_1788 = _T_1786 | reset; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@172763.4]
  assign _T_1789 = ~_T_1788; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@172764.4]
  assign _T_1791 = _T_1780 + 32'h1; // @[Monitor.scala 689:26:freechips.rocketchip.system.DefaultRV32Config.fir@172770.4]
  assign _T_1794 = _T_1426 | _T_1475; // @[Monitor.scala 690:27:freechips.rocketchip.system.DefaultRV32Config.fir@172774.4]
  assign _T_1806 = _T_1804 - 10'h1; // @[Edges.scala 231:28:freechips.rocketchip.system.DefaultRV32Config.fir@172789.4]
  assign _T_1807 = _T_1804 == 10'h0; // @[Edges.scala 232:25:freechips.rocketchip.system.DefaultRV32Config.fir@172790.4]
  assign _T_1817 = _T_1475 & _T_1807; // @[Monitor.scala 700:27:freechips.rocketchip.system.DefaultRV32Config.fir@172804.4]
  assign _T_1820 = ~io_in_d_bits_opcode[1]; // @[Edges.scala 72:43:freechips.rocketchip.system.DefaultRV32Config.fir@172807.4]
  assign _T_1821 = io_in_d_bits_opcode[2] & _T_1820; // @[Edges.scala 72:40:freechips.rocketchip.system.DefaultRV32Config.fir@172808.4]
  assign _T_1822 = _T_1817 & _T_1821; // @[Monitor.scala 700:38:freechips.rocketchip.system.DefaultRV32Config.fir@172809.4]
  assign _T_1823 = 4'h1 << io_in_d_bits_sink; // @[OneHot.scala 58:35:freechips.rocketchip.system.DefaultRV32Config.fir@172811.6]
  assign _T_1824 = _T_1795 >> io_in_d_bits_sink; // @[Monitor.scala 702:23:freechips.rocketchip.system.DefaultRV32Config.fir@172813.6]
  assign _T_1826 = ~_T_1824[0]; // @[Monitor.scala 702:14:freechips.rocketchip.system.DefaultRV32Config.fir@172815.6]
  assign _T_1828 = _T_1826 | reset; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@172817.6]
  assign _T_1829 = ~_T_1828; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@172818.6]
  assign _GEN_69 = _T_1822 ? _T_1823 : 4'h0; // @[Monitor.scala 700:72:freechips.rocketchip.system.DefaultRV32Config.fir@172810.4]
  assign _T_1831 = io_in_e_ready & io_in_e_valid; // @[Decoupled.scala 40:37:freechips.rocketchip.system.DefaultRV32Config.fir@172826.4]
  assign _T_1834 = 4'h1 << io_in_e_bits_sink; // @[OneHot.scala 58:35:freechips.rocketchip.system.DefaultRV32Config.fir@172830.6]
  assign _T_1835 = _GEN_69 | _T_1795; // @[Monitor.scala 708:24:freechips.rocketchip.system.DefaultRV32Config.fir@172832.6]
  assign _T_1836 = _T_1835 >> io_in_e_bits_sink; // @[Monitor.scala 708:35:freechips.rocketchip.system.DefaultRV32Config.fir@172833.6]
  assign _T_1839 = _T_1836[0] | reset; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@172836.6]
  assign _T_1840 = ~_T_1839; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@172837.6]
  assign _GEN_70 = _T_1831 ? _T_1834 : 4'h0; // @[Monitor.scala 706:73:freechips.rocketchip.system.DefaultRV32Config.fir@172829.4]
  assign _T_1841 = _T_1795 | _GEN_69; // @[Monitor.scala 713:27:freechips.rocketchip.system.DefaultRV32Config.fir@172843.4]
  assign _T_1842 = ~_GEN_70; // @[Monitor.scala 713:38:freechips.rocketchip.system.DefaultRV32Config.fir@172844.4]
  assign _T_1843 = _T_1841 & _T_1842; // @[Monitor.scala 713:36:freechips.rocketchip.system.DefaultRV32Config.fir@172845.4]
  assign _GEN_85 = io_in_a_valid & _T_67; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@170087.10]
  assign _GEN_99 = io_in_a_valid & _T_154; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@170212.10]
  assign _GEN_115 = io_in_a_valid & _T_245; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@170348.10]
  assign _GEN_125 = io_in_a_valid & _T_319; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@170455.10]
  assign _GEN_135 = io_in_a_valid & _T_396; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@170554.10]
  assign _GEN_145 = io_in_a_valid & _T_475; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@170645.10]
  assign _GEN_155 = io_in_a_valid & _T_542; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@170734.10]
  assign _GEN_165 = io_in_a_valid & _T_609; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@170823.10]
  assign _GEN_175 = io_in_d_valid & _T_689; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@170889.10]
  assign _GEN_185 = io_in_d_valid & _T_709; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@170931.10]
  assign _GEN_195 = io_in_d_valid & _T_737; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@170989.10]
  assign _GEN_205 = io_in_d_valid & _T_766; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@171048.10]
  assign _GEN_211 = io_in_d_valid & _T_783; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@171083.10]
  assign _GEN_217 = io_in_d_valid & _T_801; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@171119.10]
  assign _GEN_223 = io_in_b_valid & _T_931; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@171301.10]
  assign _GEN_235 = io_in_b_valid & _T_964; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@171356.10]
  assign _GEN_247 = io_in_b_valid & _T_989; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@171411.10]
  assign _GEN_257 = io_in_b_valid & _T_1010; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@171458.10]
  assign _GEN_267 = io_in_b_valid & _T_1033; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@171507.10]
  assign _GEN_275 = io_in_b_valid & _T_1054; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@171554.10]
  assign _GEN_283 = io_in_b_valid & _T_1075; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@171601.10]
  assign _GEN_293 = io_in_c_valid & _T_1172; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@171745.10]
  assign _GEN_303 = io_in_c_valid & _T_1194; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@171793.10]
  assign _GEN_313 = io_in_c_valid & _T_1212; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@171882.10]
  assign _GEN_325 = io_in_c_valid & _T_1294; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@171998.10]
  assign _GEN_337 = io_in_c_valid & _T_1372; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@172057.10]
  assign _GEN_345 = io_in_c_valid & _T_1390; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@172097.10]
  assign _GEN_353 = io_in_c_valid & _T_1404; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@172129.10]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_1435 = _RAND_0[9:0];
  _RAND_1 = {1{`RANDOM}};
  _T_1446 = _RAND_1[2:0];
  _RAND_2 = {1{`RANDOM}};
  _T_1447 = _RAND_2[2:0];
  _RAND_3 = {1{`RANDOM}};
  _T_1448 = _RAND_3[3:0];
  _RAND_4 = {1{`RANDOM}};
  _T_1449 = _RAND_4[0:0];
  _RAND_5 = {1{`RANDOM}};
  _T_1450 = _RAND_5[31:0];
  _RAND_6 = {1{`RANDOM}};
  _T_1483 = _RAND_6[9:0];
  _RAND_7 = {1{`RANDOM}};
  _T_1494 = _RAND_7[2:0];
  _RAND_8 = {1{`RANDOM}};
  _T_1495 = _RAND_8[1:0];
  _RAND_9 = {1{`RANDOM}};
  _T_1496 = _RAND_9[3:0];
  _RAND_10 = {1{`RANDOM}};
  _T_1497 = _RAND_10[0:0];
  _RAND_11 = {1{`RANDOM}};
  _T_1498 = _RAND_11[1:0];
  _RAND_12 = {1{`RANDOM}};
  _T_1499 = _RAND_12[0:0];
  _RAND_13 = {1{`RANDOM}};
  _T_1537 = _RAND_13[9:0];
  _RAND_14 = {1{`RANDOM}};
  _T_1548 = _RAND_14[2:0];
  _RAND_15 = {1{`RANDOM}};
  _T_1549 = _RAND_15[1:0];
  _RAND_16 = {1{`RANDOM}};
  _T_1550 = _RAND_16[3:0];
  _RAND_17 = {1{`RANDOM}};
  _T_1551 = _RAND_17[0:0];
  _RAND_18 = {1{`RANDOM}};
  _T_1552 = _RAND_18[31:0];
  _RAND_19 = {1{`RANDOM}};
  _T_1585 = _RAND_19[9:0];
  _RAND_20 = {1{`RANDOM}};
  _T_1596 = _RAND_20[2:0];
  _RAND_21 = {1{`RANDOM}};
  _T_1597 = _RAND_21[2:0];
  _RAND_22 = {1{`RANDOM}};
  _T_1598 = _RAND_22[3:0];
  _RAND_23 = {1{`RANDOM}};
  _T_1599 = _RAND_23[0:0];
  _RAND_24 = {1{`RANDOM}};
  _T_1600 = _RAND_24[31:0];
  _RAND_25 = {1{`RANDOM}};
  inflight = _RAND_25[1:0];
  _RAND_26 = {1{`RANDOM}};
  inflight_opcodes = _RAND_26[7:0];
  _RAND_27 = {1{`RANDOM}};
  inflight_sizes = _RAND_27[15:0];
  _RAND_28 = {1{`RANDOM}};
  _T_1634 = _RAND_28[9:0];
  _RAND_29 = {1{`RANDOM}};
  _T_1652 = _RAND_29[9:0];
  _RAND_30 = {1{`RANDOM}};
  _T_1780 = _RAND_30[31:0];
  _RAND_31 = {1{`RANDOM}};
  _T_1795 = _RAND_31[3:0];
  _RAND_32 = {1{`RANDOM}};
  _T_1804 = _RAND_32[9:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      _T_1435 <= 10'h0;
    end else if (_T_1426) begin
      if (_T_1438) begin
        if (_T_1433) begin
          _T_1435 <= _T_11[11:2];
        end else begin
          _T_1435 <= 10'h0;
        end
      end else begin
        _T_1435 <= _T_1437;
      end
    end
    if (_T_1474) begin
      _T_1446 <= io_in_a_bits_opcode;
    end
    if (_T_1474) begin
      _T_1447 <= io_in_a_bits_param;
    end
    if (_T_1474) begin
      _T_1448 <= io_in_a_bits_size;
    end
    if (_T_1474) begin
      _T_1449 <= io_in_a_bits_source;
    end
    if (_T_1474) begin
      _T_1450 <= io_in_a_bits_address;
    end
    if (reset) begin
      _T_1483 <= 10'h0;
    end else if (_T_1475) begin
      if (_T_1486) begin
        if (io_in_d_bits_opcode[0]) begin
          _T_1483 <= _T_1479[11:2];
        end else begin
          _T_1483 <= 10'h0;
        end
      end else begin
        _T_1483 <= _T_1485;
      end
    end
    if (_T_1527) begin
      _T_1494 <= io_in_d_bits_opcode;
    end
    if (_T_1527) begin
      _T_1495 <= io_in_d_bits_param;
    end
    if (_T_1527) begin
      _T_1496 <= io_in_d_bits_size;
    end
    if (_T_1527) begin
      _T_1497 <= io_in_d_bits_source;
    end
    if (_T_1527) begin
      _T_1498 <= io_in_d_bits_sink;
    end
    if (_T_1527) begin
      _T_1499 <= io_in_d_bits_denied;
    end
    if (reset) begin
      _T_1537 <= 10'h0;
    end else if (_T_1528) begin
      if (_T_1540) begin
        _T_1537 <= 10'h0;
      end else begin
        _T_1537 <= _T_1539;
      end
    end
    if (_T_1576) begin
      _T_1548 <= io_in_b_bits_opcode;
    end
    if (_T_1576) begin
      _T_1549 <= io_in_b_bits_param;
    end
    if (_T_1576) begin
      _T_1550 <= io_in_b_bits_size;
    end
    if (_T_1576) begin
      _T_1551 <= io_in_b_bits_source;
    end
    if (_T_1576) begin
      _T_1552 <= io_in_b_bits_address;
    end
    if (reset) begin
      _T_1585 <= 10'h0;
    end else if (_T_1577) begin
      if (_T_1588) begin
        if (io_in_c_bits_opcode[0]) begin
          _T_1585 <= _T_1107[11:2];
        end else begin
          _T_1585 <= 10'h0;
        end
      end else begin
        _T_1585 <= _T_1587;
      end
    end
    if (_T_1624) begin
      _T_1596 <= io_in_c_bits_opcode;
    end
    if (_T_1624) begin
      _T_1597 <= io_in_c_bits_param;
    end
    if (_T_1624) begin
      _T_1598 <= io_in_c_bits_size;
    end
    if (_T_1624) begin
      _T_1599 <= io_in_c_bits_source;
    end
    if (_T_1624) begin
      _T_1600 <= io_in_c_bits_address;
    end
    if (reset) begin
      inflight <= 2'h0;
    end else begin
      inflight <= _T_1773;
    end
    if (reset) begin
      inflight_opcodes <= 8'h0;
    end else begin
      inflight_opcodes <= _T_1776;
    end
    if (reset) begin
      inflight_sizes <= 16'h0;
    end else begin
      inflight_sizes <= _T_1779;
    end
    if (reset) begin
      _T_1634 <= 10'h0;
    end else if (_T_1426) begin
      if (a_first) begin
        if (_T_1433) begin
          _T_1634 <= _T_11[11:2];
        end else begin
          _T_1634 <= 10'h0;
        end
      end else begin
        _T_1634 <= _T_1636;
      end
    end
    if (reset) begin
      _T_1652 <= 10'h0;
    end else if (_T_1475) begin
      if (d_first) begin
        if (io_in_d_bits_opcode[0]) begin
          _T_1652 <= _T_1479[11:2];
        end else begin
          _T_1652 <= 10'h0;
        end
      end else begin
        _T_1652 <= _T_1654;
      end
    end
    if (reset) begin
      _T_1780 <= 32'h0;
    end else if (_T_1794) begin
      _T_1780 <= 32'h0;
    end else begin
      _T_1780 <= _T_1791;
    end
    if (reset) begin
      _T_1795 <= 4'h0;
    end else begin
      _T_1795 <= _T_1843;
    end
    if (reset) begin
      _T_1804 <= 10'h0;
    end else if (_T_1475) begin
      if (_T_1807) begin
        if (io_in_d_bits_opcode[0]) begin
          _T_1804 <= _T_1479[11:2];
        end else begin
          _T_1804 <= 10'h0;
        end
      end else begin
        _T_1804 <= _T_1806;
      end
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_85 & _T_119) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel carries AcquireBlock type unsupported by manager (connected at HellaCache.scala:254:21)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@170087.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_85 & _T_119) begin
          $fatal; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@170088.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_85 & _T_130) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel carries AcquireBlock from a client which does not support Probe (connected at HellaCache.scala:254:21)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@170106.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_85 & _T_130) begin
          $fatal; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@170107.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_85 & _T_133) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel AcquireBlock carries invalid source ID (connected at HellaCache.scala:254:21)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@170113.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_85 & _T_133) begin
          $fatal; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@170114.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_85 & _T_137) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel AcquireBlock smaller than a beat (connected at HellaCache.scala:254:21)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@170121.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_85 & _T_137) begin
          $fatal; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@170122.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_85 & _T_140) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel AcquireBlock address not aligned to size (connected at HellaCache.scala:254:21)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@170128.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_85 & _T_140) begin
          $fatal; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@170129.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_85 & _T_144) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel AcquireBlock carries invalid grow param (connected at HellaCache.scala:254:21)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@170136.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_85 & _T_144) begin
          $fatal; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@170137.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_85 & _T_149) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel AcquireBlock contains invalid mask (connected at HellaCache.scala:254:21)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@170145.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_85 & _T_149) begin
          $fatal; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@170146.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_99 & _T_119) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel carries AcquirePerm type unsupported by manager (connected at HellaCache.scala:254:21)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@170212.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_99 & _T_119) begin
          $fatal; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@170213.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_99 & _T_130) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel carries AcquirePerm from a client which does not support Probe (connected at HellaCache.scala:254:21)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@170231.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_99 & _T_130) begin
          $fatal; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@170232.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_99 & _T_133) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel AcquirePerm carries invalid source ID (connected at HellaCache.scala:254:21)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@170238.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_99 & _T_133) begin
          $fatal; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@170239.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_99 & _T_137) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel AcquirePerm smaller than a beat (connected at HellaCache.scala:254:21)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@170246.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_99 & _T_137) begin
          $fatal; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@170247.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_99 & _T_140) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel AcquirePerm address not aligned to size (connected at HellaCache.scala:254:21)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@170253.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_99 & _T_140) begin
          $fatal; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@170254.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_99 & _T_144) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel AcquirePerm carries invalid grow param (connected at HellaCache.scala:254:21)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@170261.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_99 & _T_144) begin
          $fatal; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@170262.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_99 & _T_235) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel AcquirePerm requests NtoB (connected at HellaCache.scala:254:21)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@170269.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_99 & _T_235) begin
          $fatal; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@170270.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_99 & _T_149) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel AcquirePerm contains invalid mask (connected at HellaCache.scala:254:21)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@170278.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_99 & _T_149) begin
          $fatal; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@170279.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_115 & _T_300) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel carries Get type unsupported by manager (connected at HellaCache.scala:254:21)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@170348.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_115 & _T_300) begin
          $fatal; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@170349.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_115 & _T_133) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel Get carries invalid source ID (connected at HellaCache.scala:254:21)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@170355.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_115 & _T_133) begin
          $fatal; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@170356.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_115 & _T_140) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel Get address not aligned to size (connected at HellaCache.scala:254:21)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@170362.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_115 & _T_140) begin
          $fatal; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@170363.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_115 & _T_310) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel Get carries invalid param (connected at HellaCache.scala:254:21)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@170370.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_115 & _T_310) begin
          $fatal; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@170371.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_115 & _T_314) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel Get contains invalid mask (connected at HellaCache.scala:254:21)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@170378.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_115 & _T_314) begin
          $fatal; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@170379.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_125 & _T_381) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel carries PutFull type unsupported by manager (connected at HellaCache.scala:254:21)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@170455.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_125 & _T_381) begin
          $fatal; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@170456.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_125 & _T_133) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel PutFull carries invalid source ID (connected at HellaCache.scala:254:21)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@170462.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_125 & _T_133) begin
          $fatal; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@170463.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_125 & _T_140) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel PutFull address not aligned to size (connected at HellaCache.scala:254:21)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@170469.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_125 & _T_140) begin
          $fatal; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@170470.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_125 & _T_310) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel PutFull carries invalid param (connected at HellaCache.scala:254:21)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@170477.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_125 & _T_310) begin
          $fatal; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@170478.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_125 & _T_314) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel PutFull contains invalid mask (connected at HellaCache.scala:254:21)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@170485.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_125 & _T_314) begin
          $fatal; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@170486.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_135 & _T_381) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel carries PutPartial type unsupported by manager (connected at HellaCache.scala:254:21)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@170554.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_135 & _T_381) begin
          $fatal; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@170555.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_135 & _T_133) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel PutPartial carries invalid source ID (connected at HellaCache.scala:254:21)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@170561.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_135 & _T_133) begin
          $fatal; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@170562.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_135 & _T_140) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel PutPartial address not aligned to size (connected at HellaCache.scala:254:21)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@170568.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_135 & _T_140) begin
          $fatal; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@170569.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_135 & _T_310) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel PutPartial carries invalid param (connected at HellaCache.scala:254:21)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@170576.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_135 & _T_310) begin
          $fatal; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@170577.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_135 & _T_474) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel PutPartial contains invalid mask (connected at HellaCache.scala:254:21)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@170586.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_135 & _T_474) begin
          $fatal; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@170587.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_145 & _T_527) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel carries Arithmetic type unsupported by manager (connected at HellaCache.scala:254:21)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@170645.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_145 & _T_527) begin
          $fatal; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@170646.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_145 & _T_133) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel Arithmetic carries invalid source ID (connected at HellaCache.scala:254:21)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@170652.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_145 & _T_133) begin
          $fatal; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@170653.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_145 & _T_140) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel Arithmetic address not aligned to size (connected at HellaCache.scala:254:21)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@170659.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_145 & _T_140) begin
          $fatal; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@170660.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_145 & _T_537) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel Arithmetic carries invalid opcode param (connected at HellaCache.scala:254:21)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@170667.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_145 & _T_537) begin
          $fatal; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@170668.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_145 & _T_314) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel Arithmetic contains invalid mask (connected at HellaCache.scala:254:21)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@170675.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_145 & _T_314) begin
          $fatal; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@170676.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_155 & _T_527) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel carries Logical type unsupported by manager (connected at HellaCache.scala:254:21)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@170734.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_155 & _T_527) begin
          $fatal; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@170735.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_155 & _T_133) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel Logical carries invalid source ID (connected at HellaCache.scala:254:21)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@170741.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_155 & _T_133) begin
          $fatal; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@170742.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_155 & _T_140) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel Logical address not aligned to size (connected at HellaCache.scala:254:21)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@170748.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_155 & _T_140) begin
          $fatal; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@170749.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_155 & _T_604) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel Logical carries invalid opcode param (connected at HellaCache.scala:254:21)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@170756.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_155 & _T_604) begin
          $fatal; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@170757.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_155 & _T_314) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel Logical contains invalid mask (connected at HellaCache.scala:254:21)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@170764.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_155 & _T_314) begin
          $fatal; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@170765.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_165 & _T_661) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel carries Hint type unsupported by manager (connected at HellaCache.scala:254:21)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@170823.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_165 & _T_661) begin
          $fatal; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@170824.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_165 & _T_133) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel Hint carries invalid source ID (connected at HellaCache.scala:254:21)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@170830.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_165 & _T_133) begin
          $fatal; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@170831.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_165 & _T_140) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel Hint address not aligned to size (connected at HellaCache.scala:254:21)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@170837.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_165 & _T_140) begin
          $fatal; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@170838.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_165 & _T_671) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel Hint carries invalid opcode param (connected at HellaCache.scala:254:21)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@170845.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_165 & _T_671) begin
          $fatal; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@170846.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_165 & _T_314) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel Hint contains invalid mask (connected at HellaCache.scala:254:21)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@170853.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_165 & _T_314) begin
          $fatal; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@170854.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_d_valid & _T_683) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel has invalid opcode (connected at HellaCache.scala:254:21)\n    at Monitor.scala:51 assert(cond, message)\n"); // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@170872.8]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_d_valid & _T_683) begin
          $fatal; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@170873.8]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_175 & _T_692) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel ReleaseAck carries invalid source ID (connected at HellaCache.scala:254:21)\n    at Monitor.scala:51 assert(cond, message)\n"); // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@170889.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_175 & _T_692) begin
          $fatal; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@170890.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_175 & _T_696) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel ReleaseAck smaller than a beat (connected at HellaCache.scala:254:21)\n    at Monitor.scala:51 assert(cond, message)\n"); // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@170897.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_175 & _T_696) begin
          $fatal; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@170898.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_175 & _T_700) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel ReleaseeAck carries invalid param (connected at HellaCache.scala:254:21)\n    at Monitor.scala:51 assert(cond, message)\n"); // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@170905.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_175 & _T_700) begin
          $fatal; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@170906.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_175 & _T_704) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel ReleaseAck is corrupt (connected at HellaCache.scala:254:21)\n    at Monitor.scala:51 assert(cond, message)\n"); // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@170913.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_175 & _T_704) begin
          $fatal; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@170914.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_175 & _T_708) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel ReleaseAck is denied (connected at HellaCache.scala:254:21)\n    at Monitor.scala:51 assert(cond, message)\n"); // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@170921.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_175 & _T_708) begin
          $fatal; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@170922.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_185 & _T_692) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel Grant carries invalid source ID (connected at HellaCache.scala:254:21)\n    at Monitor.scala:51 assert(cond, message)\n"); // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@170931.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_185 & _T_692) begin
          $fatal; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@170932.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_185 & _T_696) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel Grant smaller than a beat (connected at HellaCache.scala:254:21)\n    at Monitor.scala:51 assert(cond, message)\n"); // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@170946.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_185 & _T_696) begin
          $fatal; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@170947.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_185 & _T_723) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel Grant carries invalid cap param (connected at HellaCache.scala:254:21)\n    at Monitor.scala:51 assert(cond, message)\n"); // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@170954.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_185 & _T_723) begin
          $fatal; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@170955.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_185 & _T_727) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel Grant carries toN param (connected at HellaCache.scala:254:21)\n    at Monitor.scala:51 assert(cond, message)\n"); // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@170962.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_185 & _T_727) begin
          $fatal; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@170963.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_185 & _T_704) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel Grant is corrupt (connected at HellaCache.scala:254:21)\n    at Monitor.scala:51 assert(cond, message)\n"); // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@170970.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_185 & _T_704) begin
          $fatal; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@170971.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_195 & _T_692) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel GrantData carries invalid source ID (connected at HellaCache.scala:254:21)\n    at Monitor.scala:51 assert(cond, message)\n"); // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@170989.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_195 & _T_692) begin
          $fatal; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@170990.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_195 & _T_696) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel GrantData smaller than a beat (connected at HellaCache.scala:254:21)\n    at Monitor.scala:51 assert(cond, message)\n"); // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@171004.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_195 & _T_696) begin
          $fatal; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@171005.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_195 & _T_723) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel GrantData carries invalid cap param (connected at HellaCache.scala:254:21)\n    at Monitor.scala:51 assert(cond, message)\n"); // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@171012.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_195 & _T_723) begin
          $fatal; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@171013.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_195 & _T_727) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel GrantData carries toN param (connected at HellaCache.scala:254:21)\n    at Monitor.scala:51 assert(cond, message)\n"); // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@171020.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_195 & _T_727) begin
          $fatal; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@171021.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_195 & _T_760) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel GrantData is denied but not corrupt (connected at HellaCache.scala:254:21)\n    at Monitor.scala:51 assert(cond, message)\n"); // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@171029.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_195 & _T_760) begin
          $fatal; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@171030.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_205 & _T_692) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel AccessAck carries invalid source ID (connected at HellaCache.scala:254:21)\n    at Monitor.scala:51 assert(cond, message)\n"); // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@171048.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_205 & _T_692) begin
          $fatal; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@171049.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_205 & _T_700) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel AccessAck carries invalid param (connected at HellaCache.scala:254:21)\n    at Monitor.scala:51 assert(cond, message)\n"); // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@171056.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_205 & _T_700) begin
          $fatal; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@171057.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_205 & _T_704) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel AccessAck is corrupt (connected at HellaCache.scala:254:21)\n    at Monitor.scala:51 assert(cond, message)\n"); // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@171064.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_205 & _T_704) begin
          $fatal; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@171065.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_211 & _T_692) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel AccessAckData carries invalid source ID (connected at HellaCache.scala:254:21)\n    at Monitor.scala:51 assert(cond, message)\n"); // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@171083.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_211 & _T_692) begin
          $fatal; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@171084.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_211 & _T_700) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel AccessAckData carries invalid param (connected at HellaCache.scala:254:21)\n    at Monitor.scala:51 assert(cond, message)\n"); // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@171091.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_211 & _T_700) begin
          $fatal; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@171092.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_211 & _T_760) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel AccessAckData is denied but not corrupt (connected at HellaCache.scala:254:21)\n    at Monitor.scala:51 assert(cond, message)\n"); // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@171100.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_211 & _T_760) begin
          $fatal; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@171101.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_217 & _T_692) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel HintAck carries invalid source ID (connected at HellaCache.scala:254:21)\n    at Monitor.scala:51 assert(cond, message)\n"); // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@171119.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_217 & _T_692) begin
          $fatal; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@171120.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_217 & _T_700) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel HintAck carries invalid param (connected at HellaCache.scala:254:21)\n    at Monitor.scala:51 assert(cond, message)\n"); // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@171127.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_217 & _T_700) begin
          $fatal; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@171128.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_217 & _T_704) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel HintAck is corrupt (connected at HellaCache.scala:254:21)\n    at Monitor.scala:51 assert(cond, message)\n"); // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@171135.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_217 & _T_704) begin
          $fatal; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@171136.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_b_valid & _T_821) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel has invalid opcode (connected at HellaCache.scala:254:21)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@171155.8]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_b_valid & _T_821) begin
          $fatal; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@171156.8]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_223 & _T_942) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel carries Probe type unsupported by client (connected at HellaCache.scala:254:21)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@171301.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_223 & _T_942) begin
          $fatal; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@171302.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_223 & _T_945) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel Probe carries unmanaged address (connected at HellaCache.scala:254:21)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@171308.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_223 & _T_945) begin
          $fatal; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@171309.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_223 & _T_951) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel Probe address not aligned to size (connected at HellaCache.scala:254:21)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@171322.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_223 & _T_951) begin
          $fatal; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@171323.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_223 & _T_955) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel Probe carries invalid cap param (connected at HellaCache.scala:254:21)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@171330.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_223 & _T_955) begin
          $fatal; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@171331.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_223 & _T_959) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel Probe contains invalid mask (connected at HellaCache.scala:254:21)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@171338.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_223 & _T_959) begin
          $fatal; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@171339.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_223 & _T_963) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel Probe is corrupt (connected at HellaCache.scala:254:21)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@171346.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_223 & _T_963) begin
          $fatal; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@171347.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_235 & _T_967) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel carries Get type unsupported by client (connected at HellaCache.scala:254:21)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@171356.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_235 & _T_967) begin
          $fatal; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@171357.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_235 & _T_945) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel Get carries unmanaged address (connected at HellaCache.scala:254:21)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@171363.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_235 & _T_945) begin
          $fatal; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@171364.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_235 & _T_951) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel Get address not aligned to size (connected at HellaCache.scala:254:21)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@171377.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_235 & _T_951) begin
          $fatal; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@171378.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_235 & _T_980) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel Get carries invalid param (connected at HellaCache.scala:254:21)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@171385.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_235 & _T_980) begin
          $fatal; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@171386.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_235 & _T_959) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel Get contains invalid mask (connected at HellaCache.scala:254:21)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@171393.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_235 & _T_959) begin
          $fatal; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@171394.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_235 & _T_963) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel Get is corrupt (connected at HellaCache.scala:254:21)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@171401.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_235 & _T_963) begin
          $fatal; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@171402.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_247 & _T_967) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel carries PutFull type unsupported by client (connected at HellaCache.scala:254:21)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@171411.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_247 & _T_967) begin
          $fatal; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@171412.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_247 & _T_945) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel PutFull carries unmanaged address (connected at HellaCache.scala:254:21)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@171418.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_247 & _T_945) begin
          $fatal; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@171419.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_247 & _T_951) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel PutFull address not aligned to size (connected at HellaCache.scala:254:21)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@171432.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_247 & _T_951) begin
          $fatal; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@171433.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_247 & _T_980) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel PutFull carries invalid param (connected at HellaCache.scala:254:21)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@171440.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_247 & _T_980) begin
          $fatal; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@171441.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_247 & _T_959) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel PutFull contains invalid mask (connected at HellaCache.scala:254:21)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@171448.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_247 & _T_959) begin
          $fatal; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@171449.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_257 & _T_967) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel carries PutPartial type unsupported by client (connected at HellaCache.scala:254:21)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@171458.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_257 & _T_967) begin
          $fatal; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@171459.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_257 & _T_945) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel PutPartial carries unmanaged address (connected at HellaCache.scala:254:21)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@171465.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_257 & _T_945) begin
          $fatal; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@171466.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_257 & _T_951) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel PutPartial address not aligned to size (connected at HellaCache.scala:254:21)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@171479.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_257 & _T_951) begin
          $fatal; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@171480.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_257 & _T_980) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel PutPartial carries invalid param (connected at HellaCache.scala:254:21)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@171487.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_257 & _T_980) begin
          $fatal; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@171488.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_257 & _T_1032) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel PutPartial contains invalid mask (connected at HellaCache.scala:254:21)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@171497.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_257 & _T_1032) begin
          $fatal; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@171498.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_267 & _T_967) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel carries Arithmetic type unsupported by client (connected at HellaCache.scala:254:21)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@171507.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_267 & _T_967) begin
          $fatal; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@171508.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_267 & _T_945) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel Arithmetic carries unmanaged address (connected at HellaCache.scala:254:21)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@171514.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_267 & _T_945) begin
          $fatal; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@171515.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_267 & _T_951) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel Arithmetic address not aligned to size (connected at HellaCache.scala:254:21)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@171528.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_267 & _T_951) begin
          $fatal; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@171529.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_267 & _T_959) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel Arithmetic contains invalid mask (connected at HellaCache.scala:254:21)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@171544.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_267 & _T_959) begin
          $fatal; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@171545.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_275 & _T_967) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel carries Logical type unsupported by client (connected at HellaCache.scala:254:21)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@171554.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_275 & _T_967) begin
          $fatal; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@171555.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_275 & _T_945) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel Logical carries unmanaged address (connected at HellaCache.scala:254:21)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@171561.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_275 & _T_945) begin
          $fatal; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@171562.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_275 & _T_951) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel Logical address not aligned to size (connected at HellaCache.scala:254:21)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@171575.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_275 & _T_951) begin
          $fatal; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@171576.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_275 & _T_959) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel Logical contains invalid mask (connected at HellaCache.scala:254:21)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@171591.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_275 & _T_959) begin
          $fatal; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@171592.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_283 & _T_967) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel carries Hint type unsupported by client (connected at HellaCache.scala:254:21)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@171601.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_283 & _T_967) begin
          $fatal; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@171602.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_283 & _T_945) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel Hint carries unmanaged address (connected at HellaCache.scala:254:21)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@171608.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_283 & _T_945) begin
          $fatal; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@171609.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_283 & _T_951) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel Hint address not aligned to size (connected at HellaCache.scala:254:21)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@171622.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_283 & _T_951) begin
          $fatal; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@171623.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_283 & _T_959) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel Hint contains invalid mask (connected at HellaCache.scala:254:21)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@171630.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_283 & _T_959) begin
          $fatal; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@171631.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_283 & _T_963) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel Hint is corrupt (connected at HellaCache.scala:254:21)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@171638.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_283 & _T_963) begin
          $fatal; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@171639.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_293 & _T_1175) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel ProbeAck carries unmanaged address (connected at HellaCache.scala:254:21)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@171745.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_293 & _T_1175) begin
          $fatal; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@171746.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_293 & _T_1178) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel ProbeAck carries invalid source ID (connected at HellaCache.scala:254:21)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@171752.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_293 & _T_1178) begin
          $fatal; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@171753.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_293 & _T_1182) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel ProbeAck smaller than a beat (connected at HellaCache.scala:254:21)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@171760.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_293 & _T_1182) begin
          $fatal; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@171761.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_293 & _T_1185) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel ProbeAck address not aligned to size (connected at HellaCache.scala:254:21)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@171767.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_293 & _T_1185) begin
          $fatal; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@171768.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_293 & _T_1189) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel ProbeAck carries invalid report param (connected at HellaCache.scala:254:21)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@171775.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_293 & _T_1189) begin
          $fatal; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@171776.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_303 & _T_1175) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel ProbeAckData carries unmanaged address (connected at HellaCache.scala:254:21)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@171793.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_303 & _T_1175) begin
          $fatal; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@171794.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_303 & _T_1178) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel ProbeAckData carries invalid source ID (connected at HellaCache.scala:254:21)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@171800.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_303 & _T_1178) begin
          $fatal; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@171801.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_303 & _T_1182) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel ProbeAckData smaller than a beat (connected at HellaCache.scala:254:21)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@171808.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_303 & _T_1182) begin
          $fatal; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@171809.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_303 & _T_1185) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel ProbeAckData address not aligned to size (connected at HellaCache.scala:254:21)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@171815.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_303 & _T_1185) begin
          $fatal; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@171816.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_303 & _T_1189) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel ProbeAckData carries invalid report param (connected at HellaCache.scala:254:21)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@171823.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_303 & _T_1189) begin
          $fatal; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@171824.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_313 & _T_1264) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel carries Release type unsupported by manager (connected at HellaCache.scala:254:21)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@171882.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_313 & _T_1264) begin
          $fatal; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@171883.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_313 & _T_1275) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel carries Release from a client which does not support Probe (connected at HellaCache.scala:254:21)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@171901.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_313 & _T_1275) begin
          $fatal; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@171902.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_313 & _T_1178) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel Release carries invalid source ID (connected at HellaCache.scala:254:21)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@171908.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_313 & _T_1178) begin
          $fatal; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@171909.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_313 & _T_1182) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel Release smaller than a beat (connected at HellaCache.scala:254:21)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@171916.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_313 & _T_1182) begin
          $fatal; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@171917.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_313 & _T_1185) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel Release address not aligned to size (connected at HellaCache.scala:254:21)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@171923.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_313 & _T_1185) begin
          $fatal; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@171924.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_313 & _T_1289) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel Release carries invalid shrink param (connected at HellaCache.scala:254:21)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@171931.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_313 & _T_1289) begin
          $fatal; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@171932.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_325 & _T_1264) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel carries ReleaseData type unsupported by manager (connected at HellaCache.scala:254:21)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@171998.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_325 & _T_1264) begin
          $fatal; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@171999.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_325 & _T_1275) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel carries Release from a client which does not support Probe (connected at HellaCache.scala:254:21)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@172017.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_325 & _T_1275) begin
          $fatal; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@172018.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_325 & _T_1178) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel ReleaseData carries invalid source ID (connected at HellaCache.scala:254:21)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@172024.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_325 & _T_1178) begin
          $fatal; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@172025.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_325 & _T_1182) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel ReleaseData smaller than a beat (connected at HellaCache.scala:254:21)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@172032.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_325 & _T_1182) begin
          $fatal; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@172033.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_325 & _T_1185) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel ReleaseData address not aligned to size (connected at HellaCache.scala:254:21)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@172039.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_325 & _T_1185) begin
          $fatal; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@172040.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_325 & _T_1289) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel ReleaseData carries invalid shrink param (connected at HellaCache.scala:254:21)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@172047.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_325 & _T_1289) begin
          $fatal; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@172048.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_337 & _T_1175) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel AccessAck carries unmanaged address (connected at HellaCache.scala:254:21)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@172057.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_337 & _T_1175) begin
          $fatal; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@172058.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_337 & _T_1178) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel AccessAck carries invalid source ID (connected at HellaCache.scala:254:21)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@172064.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_337 & _T_1178) begin
          $fatal; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@172065.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_337 & _T_1185) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel AccessAck address not aligned to size (connected at HellaCache.scala:254:21)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@172071.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_337 & _T_1185) begin
          $fatal; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@172072.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_337 & _T_1385) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel AccessAck carries invalid param (connected at HellaCache.scala:254:21)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@172079.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_337 & _T_1385) begin
          $fatal; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@172080.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_345 & _T_1175) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel AccessAckData carries unmanaged address (connected at HellaCache.scala:254:21)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@172097.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_345 & _T_1175) begin
          $fatal; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@172098.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_345 & _T_1178) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel AccessAckData carries invalid source ID (connected at HellaCache.scala:254:21)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@172104.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_345 & _T_1178) begin
          $fatal; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@172105.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_345 & _T_1185) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel AccessAckData address not aligned to size (connected at HellaCache.scala:254:21)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@172111.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_345 & _T_1185) begin
          $fatal; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@172112.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_345 & _T_1385) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel AccessAckData carries invalid param (connected at HellaCache.scala:254:21)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@172119.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_345 & _T_1385) begin
          $fatal; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@172120.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_353 & _T_1175) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel HintAck carries unmanaged address (connected at HellaCache.scala:254:21)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@172129.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_353 & _T_1175) begin
          $fatal; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@172130.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_353 & _T_1178) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel HintAck carries invalid source ID (connected at HellaCache.scala:254:21)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@172136.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_353 & _T_1178) begin
          $fatal; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@172137.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_353 & _T_1185) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel HintAck address not aligned to size (connected at HellaCache.scala:254:21)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@172143.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_353 & _T_1185) begin
          $fatal; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@172144.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_353 & _T_1385) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel HintAck carries invalid param (connected at HellaCache.scala:254:21)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@172151.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_353 & _T_1385) begin
          $fatal; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@172152.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1452 & _T_1456) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel opcode changed within multibeat operation (connected at HellaCache.scala:254:21)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@172210.8]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_1452 & _T_1456) begin
          $fatal; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@172211.8]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1452 & _T_1460) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel param changed within multibeat operation (connected at HellaCache.scala:254:21)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@172218.8]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_1452 & _T_1460) begin
          $fatal; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@172219.8]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1452 & _T_1464) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel size changed within multibeat operation (connected at HellaCache.scala:254:21)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@172226.8]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_1452 & _T_1464) begin
          $fatal; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@172227.8]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1452 & _T_1468) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel source changed within multibeat operation (connected at HellaCache.scala:254:21)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@172234.8]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_1452 & _T_1468) begin
          $fatal; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@172235.8]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1452 & _T_1472) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel address changed with multibeat operation (connected at HellaCache.scala:254:21)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@172242.8]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_1452 & _T_1472) begin
          $fatal; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@172243.8]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1501 & _T_1505) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel opcode changed within multibeat operation (connected at HellaCache.scala:254:21)\n    at Monitor.scala:51 assert(cond, message)\n"); // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@172291.8]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_1501 & _T_1505) begin
          $fatal; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@172292.8]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1501 & _T_1509) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel param changed within multibeat operation (connected at HellaCache.scala:254:21)\n    at Monitor.scala:51 assert(cond, message)\n"); // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@172299.8]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_1501 & _T_1509) begin
          $fatal; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@172300.8]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1501 & _T_1513) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel size changed within multibeat operation (connected at HellaCache.scala:254:21)\n    at Monitor.scala:51 assert(cond, message)\n"); // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@172307.8]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_1501 & _T_1513) begin
          $fatal; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@172308.8]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1501 & _T_1517) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel source changed within multibeat operation (connected at HellaCache.scala:254:21)\n    at Monitor.scala:51 assert(cond, message)\n"); // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@172315.8]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_1501 & _T_1517) begin
          $fatal; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@172316.8]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1501 & _T_1521) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel sink changed with multibeat operation (connected at HellaCache.scala:254:21)\n    at Monitor.scala:51 assert(cond, message)\n"); // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@172323.8]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_1501 & _T_1521) begin
          $fatal; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@172324.8]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1501 & _T_1525) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel denied changed with multibeat operation (connected at HellaCache.scala:254:21)\n    at Monitor.scala:51 assert(cond, message)\n"); // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@172331.8]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_1501 & _T_1525) begin
          $fatal; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@172332.8]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1554 & _T_1558) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel opcode changed within multibeat operation (connected at HellaCache.scala:254:21)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@172381.8]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_1554 & _T_1558) begin
          $fatal; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@172382.8]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1554 & _T_1562) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel param changed within multibeat operation (connected at HellaCache.scala:254:21)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@172389.8]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_1554 & _T_1562) begin
          $fatal; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@172390.8]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1554 & _T_1566) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel size changed within multibeat operation (connected at HellaCache.scala:254:21)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@172397.8]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_1554 & _T_1566) begin
          $fatal; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@172398.8]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1554 & _T_1570) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel source changed within multibeat operation (connected at HellaCache.scala:254:21)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@172405.8]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_1554 & _T_1570) begin
          $fatal; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@172406.8]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1554 & _T_1574) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel addresss changed with multibeat operation (connected at HellaCache.scala:254:21)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@172413.8]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_1554 & _T_1574) begin
          $fatal; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@172414.8]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1602 & _T_1606) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel opcode changed within multibeat operation (connected at HellaCache.scala:254:21)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@172461.8]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_1602 & _T_1606) begin
          $fatal; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@172462.8]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1602 & _T_1610) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel param changed within multibeat operation (connected at HellaCache.scala:254:21)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@172469.8]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_1602 & _T_1610) begin
          $fatal; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@172470.8]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1602 & _T_1614) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel size changed within multibeat operation (connected at HellaCache.scala:254:21)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@172477.8]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_1602 & _T_1614) begin
          $fatal; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@172478.8]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1602 & _T_1618) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel source changed within multibeat operation (connected at HellaCache.scala:254:21)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@172485.8]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_1602 & _T_1618) begin
          $fatal; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@172486.8]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1602 & _T_1622) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel address changed with multibeat operation (connected at HellaCache.scala:254:21)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@172493.8]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_1602 & _T_1622) begin
          $fatal; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@172494.8]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1681 & _T_1697) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel re-used a source ID (connected at HellaCache.scala:254:21)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@172629.8]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_1681 & _T_1697) begin
          $fatal; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@172630.8]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1720 & _T_1731) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel acknowledged for nothing inflight (connected at HellaCache.scala:254:21)\n    at Monitor.scala:51 assert(cond, message)\n"); // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@172680.8]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_1720 & _T_1731) begin
          $fatal; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@172681.8]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1720 & _T_1744) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel contains improper opcode response (connected at HellaCache.scala:254:21)\n    at Monitor.scala:51 assert(cond, message)\n"); // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@172697.8]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_1720 & _T_1744) begin
          $fatal; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@172698.8]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1720 & _T_1751) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel contains improper response size (connected at HellaCache.scala:254:21)\n    at Monitor.scala:51 assert(cond, message)\n"); // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@172708.8]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_1720 & _T_1751) begin
          $fatal; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@172709.8]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1758 & _T_1763) begin
          $fwrite(32'h80000002,"Assertion failed: ready check\n    at Monitor.scala:51 assert(cond, message)\n"); // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@172726.8]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_1758 & _T_1763) begin
          $fatal; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@172727.8]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1770) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' and 'D' concurrent, despite minlatency 3 (connected at HellaCache.scala:254:21)\n    at Monitor.scala:51 assert(cond, message)\n"); // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@172738.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_1770) begin
          $fatal; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@172739.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1789) begin
          $fwrite(32'h80000002,"Assertion failed: TileLink timeout expired (connected at HellaCache.scala:254:21)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@172766.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_1789) begin
          $fatal; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@172767.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1822 & _T_1829) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel re-used a sink ID (connected at HellaCache.scala:254:21)\n    at Monitor.scala:51 assert(cond, message)\n"); // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@172820.8]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_1822 & _T_1829) begin
          $fatal; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@172821.8]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1831 & _T_1840) begin
          $fwrite(32'h80000002,"Assertion failed: 'E' channel acknowledged for nothing inflight (connected at HellaCache.scala:254:21)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@172839.8]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_1831 & _T_1840) begin
          $fatal; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@172840.8]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
  end
endmodule
