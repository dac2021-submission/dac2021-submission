module TLMonitor_7( // @[:freechips.rocketchip.system.DefaultRV32Config.fir@19303.2]
  input         clock, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@19304.4]
  input         reset, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@19305.4]
  input         io_in_a_ready, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@19306.4]
  input         io_in_a_valid, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@19306.4]
  input  [2:0]  io_in_a_bits_opcode, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@19306.4]
  input  [2:0]  io_in_a_bits_param, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@19306.4]
  input  [3:0]  io_in_a_bits_size, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@19306.4]
  input  [1:0]  io_in_a_bits_source, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@19306.4]
  input  [31:0] io_in_a_bits_address, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@19306.4]
  input  [3:0]  io_in_a_bits_mask, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@19306.4]
  input         io_in_a_bits_corrupt, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@19306.4]
  input         io_in_b_ready, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@19306.4]
  input         io_in_b_valid, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@19306.4]
  input  [1:0]  io_in_b_bits_param, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@19306.4]
  input  [31:0] io_in_b_bits_address, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@19306.4]
  input         io_in_c_ready, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@19306.4]
  input         io_in_c_valid, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@19306.4]
  input  [2:0]  io_in_c_bits_opcode, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@19306.4]
  input  [2:0]  io_in_c_bits_param, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@19306.4]
  input  [3:0]  io_in_c_bits_size, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@19306.4]
  input  [1:0]  io_in_c_bits_source, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@19306.4]
  input  [31:0] io_in_c_bits_address, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@19306.4]
  input         io_in_c_bits_corrupt, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@19306.4]
  input         io_in_d_ready, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@19306.4]
  input         io_in_d_valid, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@19306.4]
  input  [2:0]  io_in_d_bits_opcode, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@19306.4]
  input  [1:0]  io_in_d_bits_param, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@19306.4]
  input  [3:0]  io_in_d_bits_size, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@19306.4]
  input  [1:0]  io_in_d_bits_source, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@19306.4]
  input  [1:0]  io_in_d_bits_sink, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@19306.4]
  input         io_in_d_bits_denied, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@19306.4]
  input         io_in_d_bits_corrupt, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@19306.4]
  input         io_in_e_valid, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@19306.4]
  input  [1:0]  io_in_e_bits_sink // @[:freechips.rocketchip.system.DefaultRV32Config.fir@19306.4]
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
`endif // RANDOMIZE_REG_INIT
  wire [31:0] plusarg_reader_out; // @[PlusArg.scala 80:11:freechips.rocketchip.system.DefaultRV32Config.fir@22169.4]
  wire  _T_4; // @[Parameters.scala 47:9:freechips.rocketchip.system.DefaultRV32Config.fir@19317.6]
  wire  _T_5; // @[Parameters.scala 47:9:freechips.rocketchip.system.DefaultRV32Config.fir@19318.6]
  wire  _T_6; // @[Parameters.scala 47:9:freechips.rocketchip.system.DefaultRV32Config.fir@19319.6]
  wire  _T_8; // @[Parameters.scala 924:46:freechips.rocketchip.system.DefaultRV32Config.fir@19325.6]
  wire  _T_9; // @[Parameters.scala 924:46:freechips.rocketchip.system.DefaultRV32Config.fir@19326.6]
  wire [26:0] _T_11; // @[package.scala 207:77:freechips.rocketchip.system.DefaultRV32Config.fir@19328.6]
  wire [11:0] _T_13; // @[package.scala 207:46:freechips.rocketchip.system.DefaultRV32Config.fir@19330.6]
  wire [31:0] _GEN_71; // @[Edges.scala 22:16:freechips.rocketchip.system.DefaultRV32Config.fir@19331.6]
  wire [31:0] _T_14; // @[Edges.scala 22:16:freechips.rocketchip.system.DefaultRV32Config.fir@19331.6]
  wire  _T_15; // @[Edges.scala 22:24:freechips.rocketchip.system.DefaultRV32Config.fir@19332.6]
  wire [1:0] _T_18; // @[OneHot.scala 65:12:freechips.rocketchip.system.DefaultRV32Config.fir@19335.6]
  wire [1:0] _T_20; // @[Misc.scala 201:81:freechips.rocketchip.system.DefaultRV32Config.fir@19337.6]
  wire  _T_21; // @[Misc.scala 205:21:freechips.rocketchip.system.DefaultRV32Config.fir@19338.6]
  wire  _T_24; // @[Misc.scala 210:20:freechips.rocketchip.system.DefaultRV32Config.fir@19341.6]
  wire  _T_26; // @[Misc.scala 214:38:freechips.rocketchip.system.DefaultRV32Config.fir@19343.6]
  wire  _T_27; // @[Misc.scala 214:29:freechips.rocketchip.system.DefaultRV32Config.fir@19344.6]
  wire  _T_29; // @[Misc.scala 214:38:freechips.rocketchip.system.DefaultRV32Config.fir@19346.6]
  wire  _T_30; // @[Misc.scala 214:29:freechips.rocketchip.system.DefaultRV32Config.fir@19347.6]
  wire  _T_33; // @[Misc.scala 210:20:freechips.rocketchip.system.DefaultRV32Config.fir@19350.6]
  wire  _T_34; // @[Misc.scala 213:27:freechips.rocketchip.system.DefaultRV32Config.fir@19351.6]
  wire  _T_35; // @[Misc.scala 214:38:freechips.rocketchip.system.DefaultRV32Config.fir@19352.6]
  wire  _T_36; // @[Misc.scala 214:29:freechips.rocketchip.system.DefaultRV32Config.fir@19353.6]
  wire  _T_37; // @[Misc.scala 213:27:freechips.rocketchip.system.DefaultRV32Config.fir@19354.6]
  wire  _T_38; // @[Misc.scala 214:38:freechips.rocketchip.system.DefaultRV32Config.fir@19355.6]
  wire  _T_39; // @[Misc.scala 214:29:freechips.rocketchip.system.DefaultRV32Config.fir@19356.6]
  wire  _T_40; // @[Misc.scala 213:27:freechips.rocketchip.system.DefaultRV32Config.fir@19357.6]
  wire  _T_41; // @[Misc.scala 214:38:freechips.rocketchip.system.DefaultRV32Config.fir@19358.6]
  wire  _T_42; // @[Misc.scala 214:29:freechips.rocketchip.system.DefaultRV32Config.fir@19359.6]
  wire  _T_43; // @[Misc.scala 213:27:freechips.rocketchip.system.DefaultRV32Config.fir@19360.6]
  wire  _T_44; // @[Misc.scala 214:38:freechips.rocketchip.system.DefaultRV32Config.fir@19361.6]
  wire  _T_45; // @[Misc.scala 214:29:freechips.rocketchip.system.DefaultRV32Config.fir@19362.6]
  wire [3:0] _T_48; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@19365.6]
  wire [32:0] _T_52; // @[Parameters.scala 137:49:freechips.rocketchip.system.DefaultRV32Config.fir@19369.6]
  wire  _T_78; // @[Monitor.scala 79:25:freechips.rocketchip.system.DefaultRV32Config.fir@19399.6]
  wire [32:0] _T_83; // @[Parameters.scala 137:52:freechips.rocketchip.system.DefaultRV32Config.fir@19405.8]
  wire  _T_84; // @[Parameters.scala 137:67:freechips.rocketchip.system.DefaultRV32Config.fir@19406.8]
  wire [31:0] _T_85; // @[Parameters.scala 137:31:freechips.rocketchip.system.DefaultRV32Config.fir@19407.8]
  wire [32:0] _T_86; // @[Parameters.scala 137:49:freechips.rocketchip.system.DefaultRV32Config.fir@19408.8]
  wire [32:0] _T_88; // @[Parameters.scala 137:52:freechips.rocketchip.system.DefaultRV32Config.fir@19410.8]
  wire  _T_89; // @[Parameters.scala 137:67:freechips.rocketchip.system.DefaultRV32Config.fir@19411.8]
  wire [31:0] _T_90; // @[Parameters.scala 137:31:freechips.rocketchip.system.DefaultRV32Config.fir@19412.8]
  wire [32:0] _T_91; // @[Parameters.scala 137:49:freechips.rocketchip.system.DefaultRV32Config.fir@19413.8]
  wire [32:0] _T_93; // @[Parameters.scala 137:52:freechips.rocketchip.system.DefaultRV32Config.fir@19415.8]
  wire  _T_94; // @[Parameters.scala 137:67:freechips.rocketchip.system.DefaultRV32Config.fir@19416.8]
  wire [31:0] _T_95; // @[Parameters.scala 137:31:freechips.rocketchip.system.DefaultRV32Config.fir@19417.8]
  wire [32:0] _T_96; // @[Parameters.scala 137:49:freechips.rocketchip.system.DefaultRV32Config.fir@19418.8]
  wire [32:0] _T_98; // @[Parameters.scala 137:52:freechips.rocketchip.system.DefaultRV32Config.fir@19420.8]
  wire  _T_99; // @[Parameters.scala 137:67:freechips.rocketchip.system.DefaultRV32Config.fir@19421.8]
  wire [31:0] _T_100; // @[Parameters.scala 137:31:freechips.rocketchip.system.DefaultRV32Config.fir@19422.8]
  wire [32:0] _T_101; // @[Parameters.scala 137:49:freechips.rocketchip.system.DefaultRV32Config.fir@19423.8]
  wire [32:0] _T_103; // @[Parameters.scala 137:52:freechips.rocketchip.system.DefaultRV32Config.fir@19425.8]
  wire  _T_104; // @[Parameters.scala 137:67:freechips.rocketchip.system.DefaultRV32Config.fir@19426.8]
  wire [31:0] _T_105; // @[Parameters.scala 137:31:freechips.rocketchip.system.DefaultRV32Config.fir@19427.8]
  wire [32:0] _T_106; // @[Parameters.scala 137:49:freechips.rocketchip.system.DefaultRV32Config.fir@19428.8]
  wire [32:0] _T_108; // @[Parameters.scala 137:52:freechips.rocketchip.system.DefaultRV32Config.fir@19430.8]
  wire  _T_109; // @[Parameters.scala 137:67:freechips.rocketchip.system.DefaultRV32Config.fir@19431.8]
  wire  _T_110; // @[Parameters.scala 552:42:freechips.rocketchip.system.DefaultRV32Config.fir@19432.8]
  wire  _T_117; // @[Parameters.scala 93:42:freechips.rocketchip.system.DefaultRV32Config.fir@19439.8]
  wire [31:0] _T_120; // @[Parameters.scala 137:31:freechips.rocketchip.system.DefaultRV32Config.fir@19442.8]
  wire [32:0] _T_121; // @[Parameters.scala 137:49:freechips.rocketchip.system.DefaultRV32Config.fir@19443.8]
  wire [32:0] _T_123; // @[Parameters.scala 137:52:freechips.rocketchip.system.DefaultRV32Config.fir@19445.8]
  wire  _T_124; // @[Parameters.scala 137:67:freechips.rocketchip.system.DefaultRV32Config.fir@19446.8]
  wire  _T_125; // @[Parameters.scala 551:56:freechips.rocketchip.system.DefaultRV32Config.fir@19447.8]
  wire  _T_129; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@19451.8]
  wire  _T_130; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@19452.8]
  wire  _T_135; // @[Parameters.scala 92:48:freechips.rocketchip.system.DefaultRV32Config.fir@19465.8]
  wire  _T_136; // @[Mux.scala 27:72:freechips.rocketchip.system.DefaultRV32Config.fir@19466.8]
  wire  _T_143; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@19474.8]
  wire  _T_144; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@19475.8]
  wire  _T_146; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@19481.8]
  wire  _T_147; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@19482.8]
  wire  _T_150; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@19489.8]
  wire  _T_151; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@19490.8]
  wire  _T_153; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@19496.8]
  wire  _T_154; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@19497.8]
  wire  _T_155; // @[Bundles.scala 110:27:freechips.rocketchip.system.DefaultRV32Config.fir@19502.8]
  wire  _T_157; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@19504.8]
  wire  _T_158; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@19505.8]
  wire [3:0] _T_159; // @[Monitor.scala 86:18:freechips.rocketchip.system.DefaultRV32Config.fir@19510.8]
  wire  _T_160; // @[Monitor.scala 86:31:freechips.rocketchip.system.DefaultRV32Config.fir@19511.8]
  wire  _T_162; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@19513.8]
  wire  _T_163; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@19514.8]
  wire  _T_164; // @[Monitor.scala 87:18:freechips.rocketchip.system.DefaultRV32Config.fir@19519.8]
  wire  _T_166; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@19521.8]
  wire  _T_167; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@19522.8]
  wire  _T_168; // @[Monitor.scala 90:25:freechips.rocketchip.system.DefaultRV32Config.fir@19528.6]
  wire  _T_249; // @[Monitor.scala 97:31:freechips.rocketchip.system.DefaultRV32Config.fir@19639.8]
  wire  _T_251; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@19641.8]
  wire  _T_252; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@19642.8]
  wire  _T_262; // @[Monitor.scala 102:25:freechips.rocketchip.system.DefaultRV32Config.fir@19665.6]
  wire  _T_264; // @[Parameters.scala 93:42:freechips.rocketchip.system.DefaultRV32Config.fir@19668.8]
  wire  _T_272; // @[Parameters.scala 551:56:freechips.rocketchip.system.DefaultRV32Config.fir@19676.8]
  wire  _T_307; // @[Parameters.scala 552:42:freechips.rocketchip.system.DefaultRV32Config.fir@19711.8]
  wire  _T_308; // @[Parameters.scala 552:42:freechips.rocketchip.system.DefaultRV32Config.fir@19712.8]
  wire  _T_309; // @[Parameters.scala 552:42:freechips.rocketchip.system.DefaultRV32Config.fir@19713.8]
  wire  _T_310; // @[Parameters.scala 552:42:freechips.rocketchip.system.DefaultRV32Config.fir@19714.8]
  wire  _T_311; // @[Parameters.scala 552:42:freechips.rocketchip.system.DefaultRV32Config.fir@19715.8]
  wire  _T_312; // @[Parameters.scala 551:56:freechips.rocketchip.system.DefaultRV32Config.fir@19716.8]
  wire  _T_314; // @[Parameters.scala 553:30:freechips.rocketchip.system.DefaultRV32Config.fir@19718.8]
  wire  _T_316; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@19720.8]
  wire  _T_317; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@19721.8]
  wire  _T_324; // @[Monitor.scala 106:31:freechips.rocketchip.system.DefaultRV32Config.fir@19740.8]
  wire  _T_326; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@19742.8]
  wire  _T_327; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@19743.8]
  wire  _T_328; // @[Monitor.scala 107:30:freechips.rocketchip.system.DefaultRV32Config.fir@19748.8]
  wire  _T_330; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@19750.8]
  wire  _T_331; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@19751.8]
  wire  _T_336; // @[Monitor.scala 111:25:freechips.rocketchip.system.DefaultRV32Config.fir@19765.6]
  wire  _T_371; // @[Parameters.scala 552:42:freechips.rocketchip.system.DefaultRV32Config.fir@19801.8]
  wire  _T_372; // @[Parameters.scala 552:42:freechips.rocketchip.system.DefaultRV32Config.fir@19802.8]
  wire  _T_373; // @[Parameters.scala 552:42:freechips.rocketchip.system.DefaultRV32Config.fir@19803.8]
  wire  _T_374; // @[Parameters.scala 551:56:freechips.rocketchip.system.DefaultRV32Config.fir@19804.8]
  wire  _T_383; // @[Parameters.scala 93:42:freechips.rocketchip.system.DefaultRV32Config.fir@19813.8]
  wire  _T_391; // @[Parameters.scala 551:56:freechips.rocketchip.system.DefaultRV32Config.fir@19821.8]
  wire  _T_393; // @[Parameters.scala 553:30:freechips.rocketchip.system.DefaultRV32Config.fir@19823.8]
  wire  _T_395; // @[Parameters.scala 553:30:freechips.rocketchip.system.DefaultRV32Config.fir@19825.8]
  wire  _T_397; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@19827.8]
  wire  _T_398; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@19828.8]
  wire  _T_413; // @[Monitor.scala 119:25:freechips.rocketchip.system.DefaultRV32Config.fir@19864.6]
  wire [3:0] _T_486; // @[Monitor.scala 124:33:freechips.rocketchip.system.DefaultRV32Config.fir@19954.8]
  wire [3:0] _T_487; // @[Monitor.scala 124:31:freechips.rocketchip.system.DefaultRV32Config.fir@19955.8]
  wire  _T_488; // @[Monitor.scala 124:40:freechips.rocketchip.system.DefaultRV32Config.fir@19956.8]
  wire  _T_490; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@19958.8]
  wire  _T_491; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@19959.8]
  wire  _T_492; // @[Monitor.scala 127:25:freechips.rocketchip.system.DefaultRV32Config.fir@19965.6]
  wire  _T_494; // @[Parameters.scala 93:42:freechips.rocketchip.system.DefaultRV32Config.fir@19968.8]
  wire  _T_518; // @[Parameters.scala 552:42:freechips.rocketchip.system.DefaultRV32Config.fir@19992.8]
  wire  _T_519; // @[Parameters.scala 552:42:freechips.rocketchip.system.DefaultRV32Config.fir@19993.8]
  wire  _T_520; // @[Parameters.scala 551:56:freechips.rocketchip.system.DefaultRV32Config.fir@19994.8]
  wire  _T_543; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@20017.8]
  wire  _T_544; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@20018.8]
  wire  _T_551; // @[Bundles.scala 140:33:freechips.rocketchip.system.DefaultRV32Config.fir@20037.8]
  wire  _T_553; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@20039.8]
  wire  _T_554; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@20040.8]
  wire  _T_559; // @[Monitor.scala 135:25:freechips.rocketchip.system.DefaultRV32Config.fir@20054.6]
  wire  _T_618; // @[Bundles.scala 147:30:freechips.rocketchip.system.DefaultRV32Config.fir@20126.8]
  wire  _T_620; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@20128.8]
  wire  _T_621; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@20129.8]
  wire  _T_626; // @[Monitor.scala 143:25:freechips.rocketchip.system.DefaultRV32Config.fir@20143.6]
  wire  _T_677; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@20195.8]
  wire  _T_678; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@20196.8]
  wire  _T_685; // @[Bundles.scala 160:28:freechips.rocketchip.system.DefaultRV32Config.fir@20215.8]
  wire  _T_687; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@20217.8]
  wire  _T_688; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@20218.8]
  wire  _T_697; // @[Bundles.scala 44:24:freechips.rocketchip.system.DefaultRV32Config.fir@20242.6]
  wire  _T_699; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@20244.6]
  wire  _T_700; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@20245.6]
  wire  _T_701; // @[Parameters.scala 47:9:freechips.rocketchip.system.DefaultRV32Config.fir@20250.6]
  wire  _T_702; // @[Parameters.scala 47:9:freechips.rocketchip.system.DefaultRV32Config.fir@20251.6]
  wire  _T_703; // @[Parameters.scala 47:9:freechips.rocketchip.system.DefaultRV32Config.fir@20252.6]
  wire  _T_705; // @[Parameters.scala 924:46:freechips.rocketchip.system.DefaultRV32Config.fir@20258.6]
  wire  _T_706; // @[Parameters.scala 924:46:freechips.rocketchip.system.DefaultRV32Config.fir@20259.6]
  wire  _T_708; // @[Monitor.scala 307:25:freechips.rocketchip.system.DefaultRV32Config.fir@20261.6]
  wire  _T_710; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@20264.8]
  wire  _T_711; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@20265.8]
  wire  _T_712; // @[Monitor.scala 309:27:freechips.rocketchip.system.DefaultRV32Config.fir@20270.8]
  wire  _T_714; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@20272.8]
  wire  _T_715; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@20273.8]
  wire  _T_716; // @[Monitor.scala 310:28:freechips.rocketchip.system.DefaultRV32Config.fir@20278.8]
  wire  _T_718; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@20280.8]
  wire  _T_719; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@20281.8]
  wire  _T_720; // @[Monitor.scala 311:15:freechips.rocketchip.system.DefaultRV32Config.fir@20286.8]
  wire  _T_722; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@20288.8]
  wire  _T_723; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@20289.8]
  wire  _T_724; // @[Monitor.scala 312:15:freechips.rocketchip.system.DefaultRV32Config.fir@20294.8]
  wire  _T_726; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@20296.8]
  wire  _T_727; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@20297.8]
  wire  _T_728; // @[Monitor.scala 315:25:freechips.rocketchip.system.DefaultRV32Config.fir@20303.6]
  wire  _T_739; // @[Bundles.scala 104:26:freechips.rocketchip.system.DefaultRV32Config.fir@20327.8]
  wire  _T_741; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@20329.8]
  wire  _T_742; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@20330.8]
  wire  _T_743; // @[Monitor.scala 320:28:freechips.rocketchip.system.DefaultRV32Config.fir@20335.8]
  wire  _T_745; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@20337.8]
  wire  _T_746; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@20338.8]
  wire  _T_756; // @[Monitor.scala 325:25:freechips.rocketchip.system.DefaultRV32Config.fir@20361.6]
  wire  _T_776; // @[Monitor.scala 331:30:freechips.rocketchip.system.DefaultRV32Config.fir@20402.8]
  wire  _T_778; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@20404.8]
  wire  _T_779; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@20405.8]
  wire  _T_785; // @[Monitor.scala 335:25:freechips.rocketchip.system.DefaultRV32Config.fir@20420.6]
  wire  _T_802; // @[Monitor.scala 343:25:freechips.rocketchip.system.DefaultRV32Config.fir@20455.6]
  wire  _T_820; // @[Monitor.scala 351:25:freechips.rocketchip.system.DefaultRV32Config.fir@20491.6]
  wire [32:0] _T_844; // @[Parameters.scala 137:49:freechips.rocketchip.system.DefaultRV32Config.fir@20539.6]
  wire [31:0] _T_870; // @[Parameters.scala 137:31:freechips.rocketchip.system.DefaultRV32Config.fir@20569.6]
  wire [32:0] _T_871; // @[Parameters.scala 137:49:freechips.rocketchip.system.DefaultRV32Config.fir@20570.6]
  wire [32:0] _T_873; // @[Parameters.scala 137:52:freechips.rocketchip.system.DefaultRV32Config.fir@20572.6]
  wire  _T_874; // @[Parameters.scala 137:67:freechips.rocketchip.system.DefaultRV32Config.fir@20573.6]
  wire [31:0] _T_875; // @[Parameters.scala 137:31:freechips.rocketchip.system.DefaultRV32Config.fir@20574.6]
  wire [32:0] _T_876; // @[Parameters.scala 137:49:freechips.rocketchip.system.DefaultRV32Config.fir@20575.6]
  wire [32:0] _T_878; // @[Parameters.scala 137:52:freechips.rocketchip.system.DefaultRV32Config.fir@20577.6]
  wire  _T_879; // @[Parameters.scala 137:67:freechips.rocketchip.system.DefaultRV32Config.fir@20578.6]
  wire [31:0] _T_880; // @[Parameters.scala 137:31:freechips.rocketchip.system.DefaultRV32Config.fir@20579.6]
  wire [32:0] _T_881; // @[Parameters.scala 137:49:freechips.rocketchip.system.DefaultRV32Config.fir@20580.6]
  wire [32:0] _T_883; // @[Parameters.scala 137:52:freechips.rocketchip.system.DefaultRV32Config.fir@20582.6]
  wire  _T_884; // @[Parameters.scala 137:67:freechips.rocketchip.system.DefaultRV32Config.fir@20583.6]
  wire [32:0] _T_888; // @[Parameters.scala 137:52:freechips.rocketchip.system.DefaultRV32Config.fir@20587.6]
  wire  _T_889; // @[Parameters.scala 137:67:freechips.rocketchip.system.DefaultRV32Config.fir@20588.6]
  wire [31:0] _T_890; // @[Parameters.scala 137:31:freechips.rocketchip.system.DefaultRV32Config.fir@20589.6]
  wire [32:0] _T_891; // @[Parameters.scala 137:49:freechips.rocketchip.system.DefaultRV32Config.fir@20590.6]
  wire [32:0] _T_893; // @[Parameters.scala 137:52:freechips.rocketchip.system.DefaultRV32Config.fir@20592.6]
  wire  _T_894; // @[Parameters.scala 137:67:freechips.rocketchip.system.DefaultRV32Config.fir@20593.6]
  wire [31:0] _T_895; // @[Parameters.scala 137:31:freechips.rocketchip.system.DefaultRV32Config.fir@20594.6]
  wire [32:0] _T_896; // @[Parameters.scala 137:49:freechips.rocketchip.system.DefaultRV32Config.fir@20595.6]
  wire [32:0] _T_898; // @[Parameters.scala 137:52:freechips.rocketchip.system.DefaultRV32Config.fir@20597.6]
  wire  _T_899; // @[Parameters.scala 137:67:freechips.rocketchip.system.DefaultRV32Config.fir@20598.6]
  wire [31:0] _T_900; // @[Parameters.scala 137:31:freechips.rocketchip.system.DefaultRV32Config.fir@20599.6]
  wire [32:0] _T_901; // @[Parameters.scala 137:49:freechips.rocketchip.system.DefaultRV32Config.fir@20600.6]
  wire [32:0] _T_903; // @[Parameters.scala 137:52:freechips.rocketchip.system.DefaultRV32Config.fir@20602.6]
  wire  _T_904; // @[Parameters.scala 137:67:freechips.rocketchip.system.DefaultRV32Config.fir@20603.6]
  wire  _T_906; // @[Parameters.scala 535:64:freechips.rocketchip.system.DefaultRV32Config.fir@20613.6]
  wire  _T_907; // @[Parameters.scala 535:64:freechips.rocketchip.system.DefaultRV32Config.fir@20614.6]
  wire  _T_908; // @[Parameters.scala 535:64:freechips.rocketchip.system.DefaultRV32Config.fir@20615.6]
  wire  _T_909; // @[Parameters.scala 535:64:freechips.rocketchip.system.DefaultRV32Config.fir@20616.6]
  wire  _T_910; // @[Parameters.scala 535:64:freechips.rocketchip.system.DefaultRV32Config.fir@20617.6]
  wire  _T_911; // @[Parameters.scala 535:64:freechips.rocketchip.system.DefaultRV32Config.fir@20618.6]
  wire [31:0] _T_916; // @[Edges.scala 22:16:freechips.rocketchip.system.DefaultRV32Config.fir@20623.6]
  wire  _T_917; // @[Edges.scala 22:24:freechips.rocketchip.system.DefaultRV32Config.fir@20624.6]
  wire  _T_978; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@20700.8]
  wire  _T_979; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@20701.8]
  wire  _T_984; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@20714.8]
  wire  _T_985; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@20715.8]
  wire  _T_986; // @[Bundles.scala 104:26:freechips.rocketchip.system.DefaultRV32Config.fir@20720.8]
  wire  _T_988; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@20722.8]
  wire  _T_989; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@20723.8]
  wire  _T_1134; // @[Parameters.scala 47:9:freechips.rocketchip.system.DefaultRV32Config.fir@21047.6]
  wire  _T_1135; // @[Parameters.scala 47:9:freechips.rocketchip.system.DefaultRV32Config.fir@21048.6]
  wire  _T_1136; // @[Parameters.scala 47:9:freechips.rocketchip.system.DefaultRV32Config.fir@21049.6]
  wire  _T_1138; // @[Parameters.scala 924:46:freechips.rocketchip.system.DefaultRV32Config.fir@21055.6]
  wire  _T_1139; // @[Parameters.scala 924:46:freechips.rocketchip.system.DefaultRV32Config.fir@21056.6]
  wire [26:0] _T_1141; // @[package.scala 207:77:freechips.rocketchip.system.DefaultRV32Config.fir@21058.6]
  wire [11:0] _T_1143; // @[package.scala 207:46:freechips.rocketchip.system.DefaultRV32Config.fir@21060.6]
  wire [31:0] _GEN_72; // @[Edges.scala 22:16:freechips.rocketchip.system.DefaultRV32Config.fir@21061.6]
  wire [31:0] _T_1144; // @[Edges.scala 22:16:freechips.rocketchip.system.DefaultRV32Config.fir@21061.6]
  wire  _T_1145; // @[Edges.scala 22:24:freechips.rocketchip.system.DefaultRV32Config.fir@21062.6]
  wire [31:0] _T_1146; // @[Parameters.scala 137:31:freechips.rocketchip.system.DefaultRV32Config.fir@21063.6]
  wire [32:0] _T_1147; // @[Parameters.scala 137:49:freechips.rocketchip.system.DefaultRV32Config.fir@21064.6]
  wire [32:0] _T_1149; // @[Parameters.scala 137:52:freechips.rocketchip.system.DefaultRV32Config.fir@21066.6]
  wire  _T_1150; // @[Parameters.scala 137:67:freechips.rocketchip.system.DefaultRV32Config.fir@21067.6]
  wire [31:0] _T_1151; // @[Parameters.scala 137:31:freechips.rocketchip.system.DefaultRV32Config.fir@21068.6]
  wire [32:0] _T_1152; // @[Parameters.scala 137:49:freechips.rocketchip.system.DefaultRV32Config.fir@21069.6]
  wire [32:0] _T_1154; // @[Parameters.scala 137:52:freechips.rocketchip.system.DefaultRV32Config.fir@21071.6]
  wire  _T_1155; // @[Parameters.scala 137:67:freechips.rocketchip.system.DefaultRV32Config.fir@21072.6]
  wire [31:0] _T_1156; // @[Parameters.scala 137:31:freechips.rocketchip.system.DefaultRV32Config.fir@21073.6]
  wire [32:0] _T_1157; // @[Parameters.scala 137:49:freechips.rocketchip.system.DefaultRV32Config.fir@21074.6]
  wire [32:0] _T_1159; // @[Parameters.scala 137:52:freechips.rocketchip.system.DefaultRV32Config.fir@21076.6]
  wire  _T_1160; // @[Parameters.scala 137:67:freechips.rocketchip.system.DefaultRV32Config.fir@21077.6]
  wire [32:0] _T_1162; // @[Parameters.scala 137:49:freechips.rocketchip.system.DefaultRV32Config.fir@21079.6]
  wire [32:0] _T_1164; // @[Parameters.scala 137:52:freechips.rocketchip.system.DefaultRV32Config.fir@21081.6]
  wire  _T_1165; // @[Parameters.scala 137:67:freechips.rocketchip.system.DefaultRV32Config.fir@21082.6]
  wire [31:0] _T_1166; // @[Parameters.scala 137:31:freechips.rocketchip.system.DefaultRV32Config.fir@21083.6]
  wire [32:0] _T_1167; // @[Parameters.scala 137:49:freechips.rocketchip.system.DefaultRV32Config.fir@21084.6]
  wire [32:0] _T_1169; // @[Parameters.scala 137:52:freechips.rocketchip.system.DefaultRV32Config.fir@21086.6]
  wire  _T_1170; // @[Parameters.scala 137:67:freechips.rocketchip.system.DefaultRV32Config.fir@21087.6]
  wire [31:0] _T_1171; // @[Parameters.scala 137:31:freechips.rocketchip.system.DefaultRV32Config.fir@21088.6]
  wire [32:0] _T_1172; // @[Parameters.scala 137:49:freechips.rocketchip.system.DefaultRV32Config.fir@21089.6]
  wire [32:0] _T_1174; // @[Parameters.scala 137:52:freechips.rocketchip.system.DefaultRV32Config.fir@21091.6]
  wire  _T_1175; // @[Parameters.scala 137:67:freechips.rocketchip.system.DefaultRV32Config.fir@21092.6]
  wire [31:0] _T_1176; // @[Parameters.scala 137:31:freechips.rocketchip.system.DefaultRV32Config.fir@21093.6]
  wire [32:0] _T_1177; // @[Parameters.scala 137:49:freechips.rocketchip.system.DefaultRV32Config.fir@21094.6]
  wire [32:0] _T_1179; // @[Parameters.scala 137:52:freechips.rocketchip.system.DefaultRV32Config.fir@21096.6]
  wire  _T_1180; // @[Parameters.scala 137:67:freechips.rocketchip.system.DefaultRV32Config.fir@21097.6]
  wire  _T_1182; // @[Parameters.scala 535:64:freechips.rocketchip.system.DefaultRV32Config.fir@21107.6]
  wire  _T_1183; // @[Parameters.scala 535:64:freechips.rocketchip.system.DefaultRV32Config.fir@21108.6]
  wire  _T_1184; // @[Parameters.scala 535:64:freechips.rocketchip.system.DefaultRV32Config.fir@21109.6]
  wire  _T_1185; // @[Parameters.scala 535:64:freechips.rocketchip.system.DefaultRV32Config.fir@21110.6]
  wire  _T_1186; // @[Parameters.scala 535:64:freechips.rocketchip.system.DefaultRV32Config.fir@21111.6]
  wire  _T_1187; // @[Parameters.scala 535:64:freechips.rocketchip.system.DefaultRV32Config.fir@21112.6]
  wire  _T_1217; // @[Monitor.scala 239:25:freechips.rocketchip.system.DefaultRV32Config.fir@21146.6]
  wire  _T_1219; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@21149.8]
  wire  _T_1220; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@21150.8]
  wire  _T_1222; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@21156.8]
  wire  _T_1223; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@21157.8]
  wire  _T_1224; // @[Monitor.scala 242:30:freechips.rocketchip.system.DefaultRV32Config.fir@21162.8]
  wire  _T_1226; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@21164.8]
  wire  _T_1227; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@21165.8]
  wire  _T_1229; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@21171.8]
  wire  _T_1230; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@21172.8]
  wire  _T_1231; // @[Bundles.scala 122:29:freechips.rocketchip.system.DefaultRV32Config.fir@21177.8]
  wire  _T_1233; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@21179.8]
  wire  _T_1234; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@21180.8]
  wire  _T_1235; // @[Monitor.scala 245:18:freechips.rocketchip.system.DefaultRV32Config.fir@21185.8]
  wire  _T_1237; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@21187.8]
  wire  _T_1238; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@21188.8]
  wire  _T_1239; // @[Monitor.scala 248:25:freechips.rocketchip.system.DefaultRV32Config.fir@21194.6]
  wire  _T_1257; // @[Monitor.scala 256:25:freechips.rocketchip.system.DefaultRV32Config.fir@21234.6]
  wire  _T_1296; // @[Parameters.scala 93:42:freechips.rocketchip.system.DefaultRV32Config.fir@21274.8]
  wire  _T_1304; // @[Parameters.scala 551:56:freechips.rocketchip.system.DefaultRV32Config.fir@21282.8]
  wire  _T_1308; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@21286.8]
  wire  _T_1309; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@21287.8]
  wire  _T_1314; // @[Parameters.scala 92:48:freechips.rocketchip.system.DefaultRV32Config.fir@21300.8]
  wire  _T_1315; // @[Mux.scala 27:72:freechips.rocketchip.system.DefaultRV32Config.fir@21301.8]
  wire  _T_1322; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@21309.8]
  wire  _T_1323; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@21310.8]
  wire  _T_1334; // @[Bundles.scala 116:29:freechips.rocketchip.system.DefaultRV32Config.fir@21337.8]
  wire  _T_1336; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@21339.8]
  wire  _T_1337; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@21340.8]
  wire  _T_1342; // @[Monitor.scala 266:25:freechips.rocketchip.system.DefaultRV32Config.fir@21354.6]
  wire  _T_1423; // @[Monitor.scala 275:25:freechips.rocketchip.system.DefaultRV32Config.fir@21466.6]
  wire  _T_1433; // @[Monitor.scala 279:31:freechips.rocketchip.system.DefaultRV32Config.fir@21489.8]
  wire  _T_1435; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@21491.8]
  wire  _T_1436; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@21492.8]
  wire  _T_1441; // @[Monitor.scala 283:25:freechips.rocketchip.system.DefaultRV32Config.fir@21506.6]
  wire  _T_1455; // @[Monitor.scala 290:25:freechips.rocketchip.system.DefaultRV32Config.fir@21538.6]
  wire  _T_1477; // @[Decoupled.scala 40:37:freechips.rocketchip.system.DefaultRV32Config.fir@21589.4]
  wire  _T_1484; // @[Edges.scala 93:28:freechips.rocketchip.system.DefaultRV32Config.fir@21596.4]
  reg [9:0] _T_1486; // @[Edges.scala 230:27:freechips.rocketchip.system.DefaultRV32Config.fir@21598.4]
  wire [9:0] _T_1488; // @[Edges.scala 231:28:freechips.rocketchip.system.DefaultRV32Config.fir@21600.4]
  wire  _T_1489; // @[Edges.scala 232:25:freechips.rocketchip.system.DefaultRV32Config.fir@21601.4]
  reg [2:0] _T_1497; // @[Monitor.scala 381:22:freechips.rocketchip.system.DefaultRV32Config.fir@21612.4]
  reg [2:0] _T_1498; // @[Monitor.scala 382:22:freechips.rocketchip.system.DefaultRV32Config.fir@21613.4]
  reg [3:0] _T_1499; // @[Monitor.scala 383:22:freechips.rocketchip.system.DefaultRV32Config.fir@21614.4]
  reg [1:0] _T_1500; // @[Monitor.scala 384:22:freechips.rocketchip.system.DefaultRV32Config.fir@21615.4]
  reg [31:0] _T_1501; // @[Monitor.scala 385:22:freechips.rocketchip.system.DefaultRV32Config.fir@21616.4]
  wire  _T_1502; // @[Monitor.scala 386:22:freechips.rocketchip.system.DefaultRV32Config.fir@21617.4]
  wire  _T_1503; // @[Monitor.scala 386:19:freechips.rocketchip.system.DefaultRV32Config.fir@21618.4]
  wire  _T_1504; // @[Monitor.scala 387:32:freechips.rocketchip.system.DefaultRV32Config.fir@21620.6]
  wire  _T_1506; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@21622.6]
  wire  _T_1507; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@21623.6]
  wire  _T_1508; // @[Monitor.scala 388:32:freechips.rocketchip.system.DefaultRV32Config.fir@21628.6]
  wire  _T_1510; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@21630.6]
  wire  _T_1511; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@21631.6]
  wire  _T_1512; // @[Monitor.scala 389:32:freechips.rocketchip.system.DefaultRV32Config.fir@21636.6]
  wire  _T_1514; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@21638.6]
  wire  _T_1515; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@21639.6]
  wire  _T_1516; // @[Monitor.scala 390:32:freechips.rocketchip.system.DefaultRV32Config.fir@21644.6]
  wire  _T_1518; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@21646.6]
  wire  _T_1519; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@21647.6]
  wire  _T_1520; // @[Monitor.scala 391:32:freechips.rocketchip.system.DefaultRV32Config.fir@21652.6]
  wire  _T_1522; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@21654.6]
  wire  _T_1523; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@21655.6]
  wire  _T_1525; // @[Monitor.scala 393:20:freechips.rocketchip.system.DefaultRV32Config.fir@21662.4]
  wire  _T_1526; // @[Decoupled.scala 40:37:freechips.rocketchip.system.DefaultRV32Config.fir@21670.4]
  wire [26:0] _T_1528; // @[package.scala 207:77:freechips.rocketchip.system.DefaultRV32Config.fir@21672.4]
  wire [11:0] _T_1530; // @[package.scala 207:46:freechips.rocketchip.system.DefaultRV32Config.fir@21674.4]
  reg [9:0] _T_1534; // @[Edges.scala 230:27:freechips.rocketchip.system.DefaultRV32Config.fir@21678.4]
  wire [9:0] _T_1536; // @[Edges.scala 231:28:freechips.rocketchip.system.DefaultRV32Config.fir@21680.4]
  wire  _T_1537; // @[Edges.scala 232:25:freechips.rocketchip.system.DefaultRV32Config.fir@21681.4]
  reg [2:0] _T_1545; // @[Monitor.scala 532:22:freechips.rocketchip.system.DefaultRV32Config.fir@21692.4]
  reg [1:0] _T_1546; // @[Monitor.scala 533:22:freechips.rocketchip.system.DefaultRV32Config.fir@21693.4]
  reg [3:0] _T_1547; // @[Monitor.scala 534:22:freechips.rocketchip.system.DefaultRV32Config.fir@21694.4]
  reg [1:0] _T_1548; // @[Monitor.scala 535:22:freechips.rocketchip.system.DefaultRV32Config.fir@21695.4]
  reg [1:0] _T_1549; // @[Monitor.scala 536:22:freechips.rocketchip.system.DefaultRV32Config.fir@21696.4]
  reg  _T_1550; // @[Monitor.scala 537:22:freechips.rocketchip.system.DefaultRV32Config.fir@21697.4]
  wire  _T_1551; // @[Monitor.scala 538:22:freechips.rocketchip.system.DefaultRV32Config.fir@21698.4]
  wire  _T_1552; // @[Monitor.scala 538:19:freechips.rocketchip.system.DefaultRV32Config.fir@21699.4]
  wire  _T_1553; // @[Monitor.scala 539:29:freechips.rocketchip.system.DefaultRV32Config.fir@21701.6]
  wire  _T_1555; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@21703.6]
  wire  _T_1556; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@21704.6]
  wire  _T_1557; // @[Monitor.scala 540:29:freechips.rocketchip.system.DefaultRV32Config.fir@21709.6]
  wire  _T_1559; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@21711.6]
  wire  _T_1560; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@21712.6]
  wire  _T_1561; // @[Monitor.scala 541:29:freechips.rocketchip.system.DefaultRV32Config.fir@21717.6]
  wire  _T_1563; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@21719.6]
  wire  _T_1564; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@21720.6]
  wire  _T_1565; // @[Monitor.scala 542:29:freechips.rocketchip.system.DefaultRV32Config.fir@21725.6]
  wire  _T_1567; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@21727.6]
  wire  _T_1568; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@21728.6]
  wire  _T_1569; // @[Monitor.scala 543:29:freechips.rocketchip.system.DefaultRV32Config.fir@21733.6]
  wire  _T_1571; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@21735.6]
  wire  _T_1572; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@21736.6]
  wire  _T_1573; // @[Monitor.scala 544:29:freechips.rocketchip.system.DefaultRV32Config.fir@21741.6]
  wire  _T_1575; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@21743.6]
  wire  _T_1576; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@21744.6]
  wire  _T_1578; // @[Monitor.scala 546:20:freechips.rocketchip.system.DefaultRV32Config.fir@21751.4]
  wire  _T_1579; // @[Decoupled.scala 40:37:freechips.rocketchip.system.DefaultRV32Config.fir@21760.4]
  reg [9:0] _T_1588; // @[Edges.scala 230:27:freechips.rocketchip.system.DefaultRV32Config.fir@21769.4]
  wire [9:0] _T_1590; // @[Edges.scala 231:28:freechips.rocketchip.system.DefaultRV32Config.fir@21771.4]
  wire  _T_1591; // @[Edges.scala 232:25:freechips.rocketchip.system.DefaultRV32Config.fir@21772.4]
  reg [1:0] _T_1600; // @[Monitor.scala 405:22:freechips.rocketchip.system.DefaultRV32Config.fir@21784.4]
  reg [31:0] _T_1603; // @[Monitor.scala 408:22:freechips.rocketchip.system.DefaultRV32Config.fir@21787.4]
  wire  _T_1604; // @[Monitor.scala 409:22:freechips.rocketchip.system.DefaultRV32Config.fir@21788.4]
  wire  _T_1605; // @[Monitor.scala 409:19:freechips.rocketchip.system.DefaultRV32Config.fir@21789.4]
  wire  _T_1610; // @[Monitor.scala 411:32:freechips.rocketchip.system.DefaultRV32Config.fir@21799.6]
  wire  _T_1612; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@21801.6]
  wire  _T_1613; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@21802.6]
  wire  _T_1622; // @[Monitor.scala 414:32:freechips.rocketchip.system.DefaultRV32Config.fir@21823.6]
  wire  _T_1624; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@21825.6]
  wire  _T_1625; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@21826.6]
  wire  _T_1627; // @[Monitor.scala 416:20:freechips.rocketchip.system.DefaultRV32Config.fir@21833.4]
  wire  _T_1628; // @[Decoupled.scala 40:37:freechips.rocketchip.system.DefaultRV32Config.fir@21841.4]
  reg [9:0] _T_1636; // @[Edges.scala 230:27:freechips.rocketchip.system.DefaultRV32Config.fir@21849.4]
  wire [9:0] _T_1638; // @[Edges.scala 231:28:freechips.rocketchip.system.DefaultRV32Config.fir@21851.4]
  wire  _T_1639; // @[Edges.scala 232:25:freechips.rocketchip.system.DefaultRV32Config.fir@21852.4]
  reg [2:0] _T_1647; // @[Monitor.scala 509:22:freechips.rocketchip.system.DefaultRV32Config.fir@21863.4]
  reg [2:0] _T_1648; // @[Monitor.scala 510:22:freechips.rocketchip.system.DefaultRV32Config.fir@21864.4]
  reg [3:0] _T_1649; // @[Monitor.scala 511:22:freechips.rocketchip.system.DefaultRV32Config.fir@21865.4]
  reg [1:0] _T_1650; // @[Monitor.scala 512:22:freechips.rocketchip.system.DefaultRV32Config.fir@21866.4]
  reg [31:0] _T_1651; // @[Monitor.scala 513:22:freechips.rocketchip.system.DefaultRV32Config.fir@21867.4]
  wire  _T_1652; // @[Monitor.scala 514:22:freechips.rocketchip.system.DefaultRV32Config.fir@21868.4]
  wire  _T_1653; // @[Monitor.scala 514:19:freechips.rocketchip.system.DefaultRV32Config.fir@21869.4]
  wire  _T_1654; // @[Monitor.scala 515:32:freechips.rocketchip.system.DefaultRV32Config.fir@21871.6]
  wire  _T_1656; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@21873.6]
  wire  _T_1657; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@21874.6]
  wire  _T_1658; // @[Monitor.scala 516:32:freechips.rocketchip.system.DefaultRV32Config.fir@21879.6]
  wire  _T_1660; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@21881.6]
  wire  _T_1661; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@21882.6]
  wire  _T_1662; // @[Monitor.scala 517:32:freechips.rocketchip.system.DefaultRV32Config.fir@21887.6]
  wire  _T_1664; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@21889.6]
  wire  _T_1665; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@21890.6]
  wire  _T_1666; // @[Monitor.scala 518:32:freechips.rocketchip.system.DefaultRV32Config.fir@21895.6]
  wire  _T_1668; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@21897.6]
  wire  _T_1669; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@21898.6]
  wire  _T_1670; // @[Monitor.scala 519:32:freechips.rocketchip.system.DefaultRV32Config.fir@21903.6]
  wire  _T_1672; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@21905.6]
  wire  _T_1673; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@21906.6]
  wire  _T_1675; // @[Monitor.scala 521:20:freechips.rocketchip.system.DefaultRV32Config.fir@21913.4]
  reg [2:0] inflight; // @[Monitor.scala 608:27:freechips.rocketchip.system.DefaultRV32Config.fir@21921.4]
  reg [11:0] inflight_opcodes; // @[Monitor.scala 610:35:freechips.rocketchip.system.DefaultRV32Config.fir@21922.4]
  reg [23:0] inflight_sizes; // @[Monitor.scala 612:33:freechips.rocketchip.system.DefaultRV32Config.fir@21923.4]
  reg [9:0] _T_1685; // @[Edges.scala 230:27:freechips.rocketchip.system.DefaultRV32Config.fir@21933.4]
  wire [9:0] _T_1687; // @[Edges.scala 231:28:freechips.rocketchip.system.DefaultRV32Config.fir@21935.4]
  wire  a_first; // @[Edges.scala 232:25:freechips.rocketchip.system.DefaultRV32Config.fir@21936.4]
  reg [9:0] _T_1703; // @[Edges.scala 230:27:freechips.rocketchip.system.DefaultRV32Config.fir@21955.4]
  wire [9:0] _T_1705; // @[Edges.scala 231:28:freechips.rocketchip.system.DefaultRV32Config.fir@21957.4]
  wire  d_first; // @[Edges.scala 232:25:freechips.rocketchip.system.DefaultRV32Config.fir@21958.4]
  wire [3:0] _GEN_73; // @[Monitor.scala 629:69:freechips.rocketchip.system.DefaultRV32Config.fir@21977.4]
  wire [4:0] _T_1713; // @[Monitor.scala 629:69:freechips.rocketchip.system.DefaultRV32Config.fir@21977.4]
  wire [11:0] _T_1714; // @[Monitor.scala 629:44:freechips.rocketchip.system.DefaultRV32Config.fir@21978.4]
  wire [15:0] _T_1718; // @[Monitor.scala 606:57:freechips.rocketchip.system.DefaultRV32Config.fir@21982.4]
  wire [15:0] _GEN_74; // @[Monitor.scala 629:97:freechips.rocketchip.system.DefaultRV32Config.fir@21983.4]
  wire [15:0] _T_1719; // @[Monitor.scala 629:97:freechips.rocketchip.system.DefaultRV32Config.fir@21983.4]
  wire [15:0] _T_1720; // @[Monitor.scala 629:152:freechips.rocketchip.system.DefaultRV32Config.fir@21984.4]
  wire [4:0] _T_1721; // @[Monitor.scala 633:65:freechips.rocketchip.system.DefaultRV32Config.fir@21988.4]
  wire [23:0] _T_1722; // @[Monitor.scala 633:40:freechips.rocketchip.system.DefaultRV32Config.fir@21989.4]
  wire [15:0] _T_1726; // @[Monitor.scala 606:57:freechips.rocketchip.system.DefaultRV32Config.fir@21993.4]
  wire [23:0] _GEN_76; // @[Monitor.scala 633:91:freechips.rocketchip.system.DefaultRV32Config.fir@21994.4]
  wire [23:0] _T_1727; // @[Monitor.scala 633:91:freechips.rocketchip.system.DefaultRV32Config.fir@21994.4]
  wire [23:0] _T_1728; // @[Monitor.scala 633:144:freechips.rocketchip.system.DefaultRV32Config.fir@21995.4]
  wire  _T_1732; // @[Monitor.scala 643:27:freechips.rocketchip.system.DefaultRV32Config.fir@22020.4]
  wire [3:0] _T_1734; // @[OneHot.scala 58:35:freechips.rocketchip.system.DefaultRV32Config.fir@22023.6]
  wire [3:0] _T_1735; // @[Monitor.scala 645:53:freechips.rocketchip.system.DefaultRV32Config.fir@22025.6]
  wire [3:0] _T_1736; // @[Monitor.scala 645:61:freechips.rocketchip.system.DefaultRV32Config.fir@22026.6]
  wire [4:0] _T_1737; // @[Monitor.scala 646:49:freechips.rocketchip.system.DefaultRV32Config.fir@22028.6]
  wire [4:0] _T_1738; // @[Monitor.scala 646:57:freechips.rocketchip.system.DefaultRV32Config.fir@22029.6]
  wire [3:0] _GEN_78; // @[Monitor.scala 647:72:freechips.rocketchip.system.DefaultRV32Config.fir@22031.6]
  wire [4:0] _T_1739; // @[Monitor.scala 647:72:freechips.rocketchip.system.DefaultRV32Config.fir@22031.6]
  wire [3:0] a_opcodes_set_interm; // @[Monitor.scala 643:72:freechips.rocketchip.system.DefaultRV32Config.fir@22022.4]
  wire [34:0] _GEN_79; // @[Monitor.scala 647:47:freechips.rocketchip.system.DefaultRV32Config.fir@22032.6]
  wire [34:0] _T_1740; // @[Monitor.scala 647:47:freechips.rocketchip.system.DefaultRV32Config.fir@22032.6]
  wire [4:0] _T_1741; // @[Monitor.scala 648:68:freechips.rocketchip.system.DefaultRV32Config.fir@22034.6]
  wire [4:0] a_sizes_set_interm; // @[Monitor.scala 643:72:freechips.rocketchip.system.DefaultRV32Config.fir@22022.4]
  wire [35:0] _GEN_80; // @[Monitor.scala 648:43:freechips.rocketchip.system.DefaultRV32Config.fir@22035.6]
  wire [35:0] _T_1742; // @[Monitor.scala 648:43:freechips.rocketchip.system.DefaultRV32Config.fir@22035.6]
  wire [2:0] _T_1743; // @[Monitor.scala 649:26:freechips.rocketchip.system.DefaultRV32Config.fir@22037.6]
  wire  _T_1745; // @[Monitor.scala 649:17:freechips.rocketchip.system.DefaultRV32Config.fir@22039.6]
  wire  _T_1747; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@22041.6]
  wire  _T_1748; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@22042.6]
  wire [3:0] _GEN_27; // @[Monitor.scala 643:72:freechips.rocketchip.system.DefaultRV32Config.fir@22022.4]
  wire [34:0] _GEN_30; // @[Monitor.scala 643:72:freechips.rocketchip.system.DefaultRV32Config.fir@22022.4]
  wire [35:0] _GEN_31; // @[Monitor.scala 643:72:freechips.rocketchip.system.DefaultRV32Config.fir@22022.4]
  wire  _T_1751; // @[Monitor.scala 660:27:freechips.rocketchip.system.DefaultRV32Config.fir@22056.4]
  wire  _T_1753; // @[Monitor.scala 660:75:freechips.rocketchip.system.DefaultRV32Config.fir@22058.4]
  wire  _T_1754; // @[Monitor.scala 660:72:freechips.rocketchip.system.DefaultRV32Config.fir@22059.4]
  wire [3:0] _T_1755; // @[OneHot.scala 58:35:freechips.rocketchip.system.DefaultRV32Config.fir@22061.6]
  wire [46:0] _GEN_82; // @[Monitor.scala 662:76:freechips.rocketchip.system.DefaultRV32Config.fir@22068.6]
  wire [46:0] _T_1761; // @[Monitor.scala 662:76:freechips.rocketchip.system.DefaultRV32Config.fir@22068.6]
  wire [46:0] _GEN_83; // @[Monitor.scala 663:72:freechips.rocketchip.system.DefaultRV32Config.fir@22075.6]
  wire [46:0] _T_1767; // @[Monitor.scala 663:72:freechips.rocketchip.system.DefaultRV32Config.fir@22075.6]
  wire [3:0] _GEN_32; // @[Monitor.scala 660:91:freechips.rocketchip.system.DefaultRV32Config.fir@22060.4]
  wire [46:0] _GEN_33; // @[Monitor.scala 660:91:freechips.rocketchip.system.DefaultRV32Config.fir@22060.4]
  wire [46:0] _GEN_34; // @[Monitor.scala 660:91:freechips.rocketchip.system.DefaultRV32Config.fir@22060.4]
  wire  _T_1768; // @[Monitor.scala 665:26:freechips.rocketchip.system.DefaultRV32Config.fir@22078.4]
  wire  _T_1771; // @[Monitor.scala 665:71:freechips.rocketchip.system.DefaultRV32Config.fir@22081.4]
  wire [2:0] _T_1772; // @[Monitor.scala 666:25:freechips.rocketchip.system.DefaultRV32Config.fir@22083.6]
  wire  _T_1774; // @[Monitor.scala 666:93:freechips.rocketchip.system.DefaultRV32Config.fir@22085.6]
  wire  _T_1775; // @[Monitor.scala 666:68:freechips.rocketchip.system.DefaultRV32Config.fir@22086.6]
  wire  _T_1776; // @[Monitor.scala 666:142:freechips.rocketchip.system.DefaultRV32Config.fir@22087.6]
  wire  _T_1777; // @[Monitor.scala 666:119:freechips.rocketchip.system.DefaultRV32Config.fir@22088.6]
  wire  _T_1778; // @[Monitor.scala 666:166:freechips.rocketchip.system.DefaultRV32Config.fir@22089.6]
  wire  _T_1779; // @[Monitor.scala 666:49:freechips.rocketchip.system.DefaultRV32Config.fir@22090.6]
  wire  _T_1781; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@22092.6]
  wire  _T_1782; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@22093.6]
  wire [3:0] a_opcode_lookup; // @[:freechips.rocketchip.system.DefaultRV32Config.fir@21975.4 :freechips.rocketchip.system.DefaultRV32Config.fir@21976.4 Monitor.scala 629:21:freechips.rocketchip.system.DefaultRV32Config.fir@21985.4]
  wire [2:0] _GEN_37; // @[Monitor.scala 667:37:freechips.rocketchip.system.DefaultRV32Config.fir@22099.6]
  wire [2:0] _GEN_38; // @[Monitor.scala 667:37:freechips.rocketchip.system.DefaultRV32Config.fir@22099.6]
  wire [2:0] _GEN_39; // @[Monitor.scala 667:37:freechips.rocketchip.system.DefaultRV32Config.fir@22099.6]
  wire [2:0] _GEN_40; // @[Monitor.scala 667:37:freechips.rocketchip.system.DefaultRV32Config.fir@22099.6]
  wire [2:0] _GEN_41; // @[Monitor.scala 667:37:freechips.rocketchip.system.DefaultRV32Config.fir@22099.6]
  wire [2:0] _GEN_42; // @[Monitor.scala 667:37:freechips.rocketchip.system.DefaultRV32Config.fir@22099.6]
  wire  _T_1784; // @[Monitor.scala 667:37:freechips.rocketchip.system.DefaultRV32Config.fir@22099.6]
  wire [2:0] _GEN_49; // @[Monitor.scala 667:96:freechips.rocketchip.system.DefaultRV32Config.fir@22101.6]
  wire [2:0] _GEN_50; // @[Monitor.scala 667:96:freechips.rocketchip.system.DefaultRV32Config.fir@22101.6]
  wire  _T_1786; // @[Monitor.scala 667:96:freechips.rocketchip.system.DefaultRV32Config.fir@22101.6]
  wire  _T_1787; // @[Monitor.scala 667:71:freechips.rocketchip.system.DefaultRV32Config.fir@22102.6]
  wire [2:0] _GEN_53; // @[Monitor.scala 668:60:freechips.rocketchip.system.DefaultRV32Config.fir@22103.6]
  wire [2:0] _GEN_54; // @[Monitor.scala 668:60:freechips.rocketchip.system.DefaultRV32Config.fir@22103.6]
  wire [2:0] _GEN_55; // @[Monitor.scala 668:60:freechips.rocketchip.system.DefaultRV32Config.fir@22103.6]
  wire [2:0] _GEN_56; // @[Monitor.scala 668:60:freechips.rocketchip.system.DefaultRV32Config.fir@22103.6]
  wire [2:0] _GEN_57; // @[Monitor.scala 668:60:freechips.rocketchip.system.DefaultRV32Config.fir@22103.6]
  wire [2:0] _GEN_58; // @[Monitor.scala 668:60:freechips.rocketchip.system.DefaultRV32Config.fir@22103.6]
  wire  _T_1788; // @[Monitor.scala 668:60:freechips.rocketchip.system.DefaultRV32Config.fir@22103.6]
  wire [2:0] _GEN_65; // @[Monitor.scala 668:124:freechips.rocketchip.system.DefaultRV32Config.fir@22104.6]
  wire [2:0] _GEN_66; // @[Monitor.scala 668:124:freechips.rocketchip.system.DefaultRV32Config.fir@22104.6]
  wire  _T_1789; // @[Monitor.scala 668:124:freechips.rocketchip.system.DefaultRV32Config.fir@22104.6]
  wire  _T_1790; // @[Monitor.scala 668:99:freechips.rocketchip.system.DefaultRV32Config.fir@22105.6]
  wire  _T_1791; // @[Monitor.scala 668:34:freechips.rocketchip.system.DefaultRV32Config.fir@22106.6]
  wire  _T_1792; // @[Monitor.scala 668:15:freechips.rocketchip.system.DefaultRV32Config.fir@22107.6]
  wire  _T_1794; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@22109.6]
  wire  _T_1795; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@22110.6]
  wire [7:0] a_size_lookup; // @[:freechips.rocketchip.system.DefaultRV32Config.fir@21986.4 :freechips.rocketchip.system.DefaultRV32Config.fir@21987.4 Monitor.scala 633:19:freechips.rocketchip.system.DefaultRV32Config.fir@21996.4]
  wire [7:0] _GEN_84; // @[Monitor.scala 670:34:freechips.rocketchip.system.DefaultRV32Config.fir@22115.6]
  wire  _T_1796; // @[Monitor.scala 670:34:freechips.rocketchip.system.DefaultRV32Config.fir@22115.6]
  wire  _T_1798; // @[Monitor.scala 670:72:freechips.rocketchip.system.DefaultRV32Config.fir@22117.6]
  wire  _T_1799; // @[Monitor.scala 670:53:freechips.rocketchip.system.DefaultRV32Config.fir@22118.6]
  wire  _T_1801; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@22120.6]
  wire  _T_1802; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@22121.6]
  wire  _T_1804; // @[Monitor.scala 672:36:freechips.rocketchip.system.DefaultRV32Config.fir@22128.4]
  wire  _T_1805; // @[Monitor.scala 672:47:freechips.rocketchip.system.DefaultRV32Config.fir@22129.4]
  wire  _T_1807; // @[Monitor.scala 672:65:freechips.rocketchip.system.DefaultRV32Config.fir@22131.4]
  wire  _T_1809; // @[Monitor.scala 672:116:freechips.rocketchip.system.DefaultRV32Config.fir@22133.4]
  wire  _T_1810; // @[Monitor.scala 673:15:freechips.rocketchip.system.DefaultRV32Config.fir@22135.6]
  wire  _T_1811; // @[Monitor.scala 673:32:freechips.rocketchip.system.DefaultRV32Config.fir@22136.6]
  wire  _T_1813; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@22138.6]
  wire  _T_1814; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@22139.6]
  wire [2:0] a_set; // @[:freechips.rocketchip.system.DefaultRV32Config.fir@21969.4 :freechips.rocketchip.system.DefaultRV32Config.fir@21970.4 Monitor.scala 644:13:freechips.rocketchip.system.DefaultRV32Config.fir@22024.6]
  wire [2:0] d_clr; // @[:freechips.rocketchip.system.DefaultRV32Config.fir@22048.4 :freechips.rocketchip.system.DefaultRV32Config.fir@22049.4 Monitor.scala 661:13:freechips.rocketchip.system.DefaultRV32Config.fir@22062.6]
  wire  _T_1815; // @[Monitor.scala 677:20:freechips.rocketchip.system.DefaultRV32Config.fir@22145.4]
  wire  _T_1816; // @[Monitor.scala 677:40:freechips.rocketchip.system.DefaultRV32Config.fir@22146.4]
  wire  _T_1817; // @[Monitor.scala 677:33:freechips.rocketchip.system.DefaultRV32Config.fir@22147.4]
  wire  _T_1818; // @[Monitor.scala 677:30:freechips.rocketchip.system.DefaultRV32Config.fir@22148.4]
  wire  _T_1820; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@22150.4]
  wire  _T_1821; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@22151.4]
  wire [2:0] _T_1822; // @[Monitor.scala 680:27:freechips.rocketchip.system.DefaultRV32Config.fir@22156.4]
  wire [2:0] _T_1823; // @[Monitor.scala 680:38:freechips.rocketchip.system.DefaultRV32Config.fir@22157.4]
  wire [2:0] _T_1824; // @[Monitor.scala 680:36:freechips.rocketchip.system.DefaultRV32Config.fir@22158.4]
  wire [11:0] a_opcodes_set; // @[:freechips.rocketchip.system.DefaultRV32Config.fir@21971.4 :freechips.rocketchip.system.DefaultRV32Config.fir@21972.4 Monitor.scala 647:21:freechips.rocketchip.system.DefaultRV32Config.fir@22033.6]
  wire [11:0] _T_1825; // @[Monitor.scala 681:43:freechips.rocketchip.system.DefaultRV32Config.fir@22160.4]
  wire [11:0] d_opcodes_clr; // @[:freechips.rocketchip.system.DefaultRV32Config.fir@22050.4 :freechips.rocketchip.system.DefaultRV32Config.fir@22051.4 Monitor.scala 662:21:freechips.rocketchip.system.DefaultRV32Config.fir@22069.6]
  wire [11:0] _T_1826; // @[Monitor.scala 681:62:freechips.rocketchip.system.DefaultRV32Config.fir@22161.4]
  wire [11:0] _T_1827; // @[Monitor.scala 681:60:freechips.rocketchip.system.DefaultRV32Config.fir@22162.4]
  wire [23:0] a_sizes_set; // @[:freechips.rocketchip.system.DefaultRV32Config.fir@21973.4 :freechips.rocketchip.system.DefaultRV32Config.fir@21974.4 Monitor.scala 648:19:freechips.rocketchip.system.DefaultRV32Config.fir@22036.6]
  wire [23:0] _T_1828; // @[Monitor.scala 682:39:freechips.rocketchip.system.DefaultRV32Config.fir@22164.4]
  wire [23:0] d_sizes_clr; // @[:freechips.rocketchip.system.DefaultRV32Config.fir@22052.4 :freechips.rocketchip.system.DefaultRV32Config.fir@22053.4 Monitor.scala 663:19:freechips.rocketchip.system.DefaultRV32Config.fir@22076.6]
  wire [23:0] _T_1829; // @[Monitor.scala 682:56:freechips.rocketchip.system.DefaultRV32Config.fir@22165.4]
  wire [23:0] _T_1830; // @[Monitor.scala 682:54:freechips.rocketchip.system.DefaultRV32Config.fir@22166.4]
  reg [31:0] _T_1831; // @[Monitor.scala 684:27:freechips.rocketchip.system.DefaultRV32Config.fir@22168.4]
  wire  _T_1832; // @[Monitor.scala 687:26:freechips.rocketchip.system.DefaultRV32Config.fir@22171.4]
  wire  _T_1833; // @[Monitor.scala 687:16:freechips.rocketchip.system.DefaultRV32Config.fir@22172.4]
  wire  _T_1834; // @[Monitor.scala 687:39:freechips.rocketchip.system.DefaultRV32Config.fir@22173.4]
  wire  _T_1835; // @[Monitor.scala 687:30:freechips.rocketchip.system.DefaultRV32Config.fir@22174.4]
  wire  _T_1836; // @[Monitor.scala 687:59:freechips.rocketchip.system.DefaultRV32Config.fir@22175.4]
  wire  _T_1837; // @[Monitor.scala 687:47:freechips.rocketchip.system.DefaultRV32Config.fir@22176.4]
  wire  _T_1839; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@22178.4]
  wire  _T_1840; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@22179.4]
  wire [31:0] _T_1842; // @[Monitor.scala 689:26:freechips.rocketchip.system.DefaultRV32Config.fir@22185.4]
  wire  _T_1845; // @[Monitor.scala 690:27:freechips.rocketchip.system.DefaultRV32Config.fir@22189.4]
  reg [3:0] _T_1846; // @[Monitor.scala 694:27:freechips.rocketchip.system.DefaultRV32Config.fir@22193.4]
  reg [9:0] _T_1855; // @[Edges.scala 230:27:freechips.rocketchip.system.DefaultRV32Config.fir@22202.4]
  wire [9:0] _T_1857; // @[Edges.scala 231:28:freechips.rocketchip.system.DefaultRV32Config.fir@22204.4]
  wire  _T_1858; // @[Edges.scala 232:25:freechips.rocketchip.system.DefaultRV32Config.fir@22205.4]
  wire  _T_1868; // @[Monitor.scala 700:27:freechips.rocketchip.system.DefaultRV32Config.fir@22219.4]
  wire  _T_1871; // @[Edges.scala 72:43:freechips.rocketchip.system.DefaultRV32Config.fir@22222.4]
  wire  _T_1872; // @[Edges.scala 72:40:freechips.rocketchip.system.DefaultRV32Config.fir@22223.4]
  wire  _T_1873; // @[Monitor.scala 700:38:freechips.rocketchip.system.DefaultRV32Config.fir@22224.4]
  wire [3:0] _T_1874; // @[OneHot.scala 58:35:freechips.rocketchip.system.DefaultRV32Config.fir@22226.6]
  wire [3:0] _T_1875; // @[Monitor.scala 702:23:freechips.rocketchip.system.DefaultRV32Config.fir@22228.6]
  wire  _T_1877; // @[Monitor.scala 702:14:freechips.rocketchip.system.DefaultRV32Config.fir@22230.6]
  wire  _T_1879; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@22232.6]
  wire  _T_1880; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@22233.6]
  wire [3:0] _GEN_69; // @[Monitor.scala 700:72:freechips.rocketchip.system.DefaultRV32Config.fir@22225.4]
  wire [3:0] _T_1885; // @[OneHot.scala 58:35:freechips.rocketchip.system.DefaultRV32Config.fir@22245.6]
  wire [3:0] _T_1886; // @[Monitor.scala 708:24:freechips.rocketchip.system.DefaultRV32Config.fir@22247.6]
  wire [3:0] _T_1887; // @[Monitor.scala 708:35:freechips.rocketchip.system.DefaultRV32Config.fir@22248.6]
  wire  _T_1890; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@22251.6]
  wire  _T_1891; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@22252.6]
  wire [3:0] _GEN_70; // @[Monitor.scala 706:73:freechips.rocketchip.system.DefaultRV32Config.fir@22244.4]
  wire [3:0] _T_1892; // @[Monitor.scala 713:27:freechips.rocketchip.system.DefaultRV32Config.fir@22258.4]
  wire [3:0] _T_1893; // @[Monitor.scala 713:38:freechips.rocketchip.system.DefaultRV32Config.fir@22259.4]
  wire [3:0] _T_1894; // @[Monitor.scala 713:36:freechips.rocketchip.system.DefaultRV32Config.fir@22260.4]
  wire  _GEN_85; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@19454.10]
  wire  _GEN_101; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@19583.10]
  wire  _GEN_119; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@19723.10]
  wire  _GEN_131; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@19830.10]
  wire  _GEN_141; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@19929.10]
  wire  _GEN_151; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@20020.10]
  wire  _GEN_161; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@20109.10]
  wire  _GEN_171; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@20198.10]
  wire  _GEN_183; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@20267.10]
  wire  _GEN_193; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@20309.10]
  wire  _GEN_203; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@20367.10]
  wire  _GEN_213; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@20426.10]
  wire  _GEN_219; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@20461.10]
  wire  _GEN_225; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@20497.10]
  wire  _GEN_231; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@21152.10]
  wire  _GEN_243; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@21200.10]
  wire  _GEN_253; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@21289.10]
  wire  _GEN_267; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@21409.10]
  wire  _GEN_279; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@21472.10]
  wire  _GEN_289; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@21512.10]
  wire  _GEN_297; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@21544.10]
  plusarg_reader #(.FORMAT("tilelink_timeout=%d"), .DEFAULT(0), .WIDTH(32)) plusarg_reader ( // @[PlusArg.scala 80:11:freechips.rocketchip.system.DefaultRV32Config.fir@22169.4]
    .out(plusarg_reader_out)
  );
  assign _T_4 = io_in_a_bits_source == 2'h0; // @[Parameters.scala 47:9:freechips.rocketchip.system.DefaultRV32Config.fir@19317.6]
  assign _T_5 = io_in_a_bits_source == 2'h1; // @[Parameters.scala 47:9:freechips.rocketchip.system.DefaultRV32Config.fir@19318.6]
  assign _T_6 = io_in_a_bits_source == 2'h2; // @[Parameters.scala 47:9:freechips.rocketchip.system.DefaultRV32Config.fir@19319.6]
  assign _T_8 = _T_4 | _T_5; // @[Parameters.scala 924:46:freechips.rocketchip.system.DefaultRV32Config.fir@19325.6]
  assign _T_9 = _T_8 | _T_6; // @[Parameters.scala 924:46:freechips.rocketchip.system.DefaultRV32Config.fir@19326.6]
  assign _T_11 = 27'hfff << io_in_a_bits_size; // @[package.scala 207:77:freechips.rocketchip.system.DefaultRV32Config.fir@19328.6]
  assign _T_13 = ~_T_11[11:0]; // @[package.scala 207:46:freechips.rocketchip.system.DefaultRV32Config.fir@19330.6]
  assign _GEN_71 = {{20'd0}, _T_13}; // @[Edges.scala 22:16:freechips.rocketchip.system.DefaultRV32Config.fir@19331.6]
  assign _T_14 = io_in_a_bits_address & _GEN_71; // @[Edges.scala 22:16:freechips.rocketchip.system.DefaultRV32Config.fir@19331.6]
  assign _T_15 = _T_14 == 32'h0; // @[Edges.scala 22:24:freechips.rocketchip.system.DefaultRV32Config.fir@19332.6]
  assign _T_18 = 2'h1 << io_in_a_bits_size[0]; // @[OneHot.scala 65:12:freechips.rocketchip.system.DefaultRV32Config.fir@19335.6]
  assign _T_20 = _T_18 | 2'h1; // @[Misc.scala 201:81:freechips.rocketchip.system.DefaultRV32Config.fir@19337.6]
  assign _T_21 = io_in_a_bits_size >= 4'h2; // @[Misc.scala 205:21:freechips.rocketchip.system.DefaultRV32Config.fir@19338.6]
  assign _T_24 = ~io_in_a_bits_address[1]; // @[Misc.scala 210:20:freechips.rocketchip.system.DefaultRV32Config.fir@19341.6]
  assign _T_26 = _T_20[1] & _T_24; // @[Misc.scala 214:38:freechips.rocketchip.system.DefaultRV32Config.fir@19343.6]
  assign _T_27 = _T_21 | _T_26; // @[Misc.scala 214:29:freechips.rocketchip.system.DefaultRV32Config.fir@19344.6]
  assign _T_29 = _T_20[1] & io_in_a_bits_address[1]; // @[Misc.scala 214:38:freechips.rocketchip.system.DefaultRV32Config.fir@19346.6]
  assign _T_30 = _T_21 | _T_29; // @[Misc.scala 214:29:freechips.rocketchip.system.DefaultRV32Config.fir@19347.6]
  assign _T_33 = ~io_in_a_bits_address[0]; // @[Misc.scala 210:20:freechips.rocketchip.system.DefaultRV32Config.fir@19350.6]
  assign _T_34 = _T_24 & _T_33; // @[Misc.scala 213:27:freechips.rocketchip.system.DefaultRV32Config.fir@19351.6]
  assign _T_35 = _T_20[0] & _T_34; // @[Misc.scala 214:38:freechips.rocketchip.system.DefaultRV32Config.fir@19352.6]
  assign _T_36 = _T_27 | _T_35; // @[Misc.scala 214:29:freechips.rocketchip.system.DefaultRV32Config.fir@19353.6]
  assign _T_37 = _T_24 & io_in_a_bits_address[0]; // @[Misc.scala 213:27:freechips.rocketchip.system.DefaultRV32Config.fir@19354.6]
  assign _T_38 = _T_20[0] & _T_37; // @[Misc.scala 214:38:freechips.rocketchip.system.DefaultRV32Config.fir@19355.6]
  assign _T_39 = _T_27 | _T_38; // @[Misc.scala 214:29:freechips.rocketchip.system.DefaultRV32Config.fir@19356.6]
  assign _T_40 = io_in_a_bits_address[1] & _T_33; // @[Misc.scala 213:27:freechips.rocketchip.system.DefaultRV32Config.fir@19357.6]
  assign _T_41 = _T_20[0] & _T_40; // @[Misc.scala 214:38:freechips.rocketchip.system.DefaultRV32Config.fir@19358.6]
  assign _T_42 = _T_30 | _T_41; // @[Misc.scala 214:29:freechips.rocketchip.system.DefaultRV32Config.fir@19359.6]
  assign _T_43 = io_in_a_bits_address[1] & io_in_a_bits_address[0]; // @[Misc.scala 213:27:freechips.rocketchip.system.DefaultRV32Config.fir@19360.6]
  assign _T_44 = _T_20[0] & _T_43; // @[Misc.scala 214:38:freechips.rocketchip.system.DefaultRV32Config.fir@19361.6]
  assign _T_45 = _T_30 | _T_44; // @[Misc.scala 214:29:freechips.rocketchip.system.DefaultRV32Config.fir@19362.6]
  assign _T_48 = {_T_45,_T_42,_T_39,_T_36}; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@19365.6]
  assign _T_52 = {1'b0,$signed(io_in_a_bits_address)}; // @[Parameters.scala 137:49:freechips.rocketchip.system.DefaultRV32Config.fir@19369.6]
  assign _T_78 = io_in_a_bits_opcode == 3'h6; // @[Monitor.scala 79:25:freechips.rocketchip.system.DefaultRV32Config.fir@19399.6]
  assign _T_83 = $signed(_T_52) & -33'sh1000; // @[Parameters.scala 137:52:freechips.rocketchip.system.DefaultRV32Config.fir@19405.8]
  assign _T_84 = $signed(_T_83) == 33'sh0; // @[Parameters.scala 137:67:freechips.rocketchip.system.DefaultRV32Config.fir@19406.8]
  assign _T_85 = io_in_a_bits_address ^ 32'h3000; // @[Parameters.scala 137:31:freechips.rocketchip.system.DefaultRV32Config.fir@19407.8]
  assign _T_86 = {1'b0,$signed(_T_85)}; // @[Parameters.scala 137:49:freechips.rocketchip.system.DefaultRV32Config.fir@19408.8]
  assign _T_88 = $signed(_T_86) & -33'sh1000; // @[Parameters.scala 137:52:freechips.rocketchip.system.DefaultRV32Config.fir@19410.8]
  assign _T_89 = $signed(_T_88) == 33'sh0; // @[Parameters.scala 137:67:freechips.rocketchip.system.DefaultRV32Config.fir@19411.8]
  assign _T_90 = io_in_a_bits_address ^ 32'h10000; // @[Parameters.scala 137:31:freechips.rocketchip.system.DefaultRV32Config.fir@19412.8]
  assign _T_91 = {1'b0,$signed(_T_90)}; // @[Parameters.scala 137:49:freechips.rocketchip.system.DefaultRV32Config.fir@19413.8]
  assign _T_93 = $signed(_T_91) & -33'sh10000; // @[Parameters.scala 137:52:freechips.rocketchip.system.DefaultRV32Config.fir@19415.8]
  assign _T_94 = $signed(_T_93) == 33'sh0; // @[Parameters.scala 137:67:freechips.rocketchip.system.DefaultRV32Config.fir@19416.8]
  assign _T_95 = io_in_a_bits_address ^ 32'h2000000; // @[Parameters.scala 137:31:freechips.rocketchip.system.DefaultRV32Config.fir@19417.8]
  assign _T_96 = {1'b0,$signed(_T_95)}; // @[Parameters.scala 137:49:freechips.rocketchip.system.DefaultRV32Config.fir@19418.8]
  assign _T_98 = $signed(_T_96) & -33'sh10000; // @[Parameters.scala 137:52:freechips.rocketchip.system.DefaultRV32Config.fir@19420.8]
  assign _T_99 = $signed(_T_98) == 33'sh0; // @[Parameters.scala 137:67:freechips.rocketchip.system.DefaultRV32Config.fir@19421.8]
  assign _T_100 = io_in_a_bits_address ^ 32'hc000000; // @[Parameters.scala 137:31:freechips.rocketchip.system.DefaultRV32Config.fir@19422.8]
  assign _T_101 = {1'b0,$signed(_T_100)}; // @[Parameters.scala 137:49:freechips.rocketchip.system.DefaultRV32Config.fir@19423.8]
  assign _T_103 = $signed(_T_101) & -33'sh4000000; // @[Parameters.scala 137:52:freechips.rocketchip.system.DefaultRV32Config.fir@19425.8]
  assign _T_104 = $signed(_T_103) == 33'sh0; // @[Parameters.scala 137:67:freechips.rocketchip.system.DefaultRV32Config.fir@19426.8]
  assign _T_105 = io_in_a_bits_address ^ 32'h60000000; // @[Parameters.scala 137:31:freechips.rocketchip.system.DefaultRV32Config.fir@19427.8]
  assign _T_106 = {1'b0,$signed(_T_105)}; // @[Parameters.scala 137:49:freechips.rocketchip.system.DefaultRV32Config.fir@19428.8]
  assign _T_108 = $signed(_T_106) & -33'sh20000000; // @[Parameters.scala 137:52:freechips.rocketchip.system.DefaultRV32Config.fir@19430.8]
  assign _T_109 = $signed(_T_108) == 33'sh0; // @[Parameters.scala 137:67:freechips.rocketchip.system.DefaultRV32Config.fir@19431.8]
  assign _T_110 = _T_84 | _T_89; // @[Parameters.scala 552:42:freechips.rocketchip.system.DefaultRV32Config.fir@19432.8]
  assign _T_117 = io_in_a_bits_size <= 4'h6; // @[Parameters.scala 93:42:freechips.rocketchip.system.DefaultRV32Config.fir@19439.8]
  assign _T_120 = io_in_a_bits_address ^ 32'h80000000; // @[Parameters.scala 137:31:freechips.rocketchip.system.DefaultRV32Config.fir@19442.8]
  assign _T_121 = {1'b0,$signed(_T_120)}; // @[Parameters.scala 137:49:freechips.rocketchip.system.DefaultRV32Config.fir@19443.8]
  assign _T_123 = $signed(_T_121) & -33'sh10000000; // @[Parameters.scala 137:52:freechips.rocketchip.system.DefaultRV32Config.fir@19445.8]
  assign _T_124 = $signed(_T_123) == 33'sh0; // @[Parameters.scala 137:67:freechips.rocketchip.system.DefaultRV32Config.fir@19446.8]
  assign _T_125 = _T_117 & _T_124; // @[Parameters.scala 551:56:freechips.rocketchip.system.DefaultRV32Config.fir@19447.8]
  assign _T_129 = _T_125 | reset; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@19451.8]
  assign _T_130 = ~_T_129; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@19452.8]
  assign _T_135 = 4'h6 == io_in_a_bits_size; // @[Parameters.scala 92:48:freechips.rocketchip.system.DefaultRV32Config.fir@19465.8]
  assign _T_136 = _T_4 & _T_135; // @[Mux.scala 27:72:freechips.rocketchip.system.DefaultRV32Config.fir@19466.8]
  assign _T_143 = _T_136 | reset; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@19474.8]
  assign _T_144 = ~_T_143; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@19475.8]
  assign _T_146 = _T_9 | reset; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@19481.8]
  assign _T_147 = ~_T_146; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@19482.8]
  assign _T_150 = _T_21 | reset; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@19489.8]
  assign _T_151 = ~_T_150; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@19490.8]
  assign _T_153 = _T_15 | reset; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@19496.8]
  assign _T_154 = ~_T_153; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@19497.8]
  assign _T_155 = io_in_a_bits_param <= 3'h2; // @[Bundles.scala 110:27:freechips.rocketchip.system.DefaultRV32Config.fir@19502.8]
  assign _T_157 = _T_155 | reset; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@19504.8]
  assign _T_158 = ~_T_157; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@19505.8]
  assign _T_159 = ~io_in_a_bits_mask; // @[Monitor.scala 86:18:freechips.rocketchip.system.DefaultRV32Config.fir@19510.8]
  assign _T_160 = _T_159 == 4'h0; // @[Monitor.scala 86:31:freechips.rocketchip.system.DefaultRV32Config.fir@19511.8]
  assign _T_162 = _T_160 | reset; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@19513.8]
  assign _T_163 = ~_T_162; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@19514.8]
  assign _T_164 = ~io_in_a_bits_corrupt; // @[Monitor.scala 87:18:freechips.rocketchip.system.DefaultRV32Config.fir@19519.8]
  assign _T_166 = _T_164 | reset; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@19521.8]
  assign _T_167 = ~_T_166; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@19522.8]
  assign _T_168 = io_in_a_bits_opcode == 3'h7; // @[Monitor.scala 90:25:freechips.rocketchip.system.DefaultRV32Config.fir@19528.6]
  assign _T_249 = io_in_a_bits_param != 3'h0; // @[Monitor.scala 97:31:freechips.rocketchip.system.DefaultRV32Config.fir@19639.8]
  assign _T_251 = _T_249 | reset; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@19641.8]
  assign _T_252 = ~_T_251; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@19642.8]
  assign _T_262 = io_in_a_bits_opcode == 3'h4; // @[Monitor.scala 102:25:freechips.rocketchip.system.DefaultRV32Config.fir@19665.6]
  assign _T_264 = io_in_a_bits_size <= 4'hc; // @[Parameters.scala 93:42:freechips.rocketchip.system.DefaultRV32Config.fir@19668.8]
  assign _T_272 = _T_264 & _T_89; // @[Parameters.scala 551:56:freechips.rocketchip.system.DefaultRV32Config.fir@19676.8]
  assign _T_307 = _T_84 | _T_94; // @[Parameters.scala 552:42:freechips.rocketchip.system.DefaultRV32Config.fir@19711.8]
  assign _T_308 = _T_307 | _T_99; // @[Parameters.scala 552:42:freechips.rocketchip.system.DefaultRV32Config.fir@19712.8]
  assign _T_309 = _T_308 | _T_104; // @[Parameters.scala 552:42:freechips.rocketchip.system.DefaultRV32Config.fir@19713.8]
  assign _T_310 = _T_309 | _T_109; // @[Parameters.scala 552:42:freechips.rocketchip.system.DefaultRV32Config.fir@19714.8]
  assign _T_311 = _T_310 | _T_124; // @[Parameters.scala 552:42:freechips.rocketchip.system.DefaultRV32Config.fir@19715.8]
  assign _T_312 = _T_117 & _T_311; // @[Parameters.scala 551:56:freechips.rocketchip.system.DefaultRV32Config.fir@19716.8]
  assign _T_314 = _T_272 | _T_312; // @[Parameters.scala 553:30:freechips.rocketchip.system.DefaultRV32Config.fir@19718.8]
  assign _T_316 = _T_314 | reset; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@19720.8]
  assign _T_317 = ~_T_316; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@19721.8]
  assign _T_324 = io_in_a_bits_param == 3'h0; // @[Monitor.scala 106:31:freechips.rocketchip.system.DefaultRV32Config.fir@19740.8]
  assign _T_326 = _T_324 | reset; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@19742.8]
  assign _T_327 = ~_T_326; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@19743.8]
  assign _T_328 = io_in_a_bits_mask == _T_48; // @[Monitor.scala 107:30:freechips.rocketchip.system.DefaultRV32Config.fir@19748.8]
  assign _T_330 = _T_328 | reset; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@19750.8]
  assign _T_331 = ~_T_330; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@19751.8]
  assign _T_336 = io_in_a_bits_opcode == 3'h0; // @[Monitor.scala 111:25:freechips.rocketchip.system.DefaultRV32Config.fir@19765.6]
  assign _T_371 = _T_84 | _T_99; // @[Parameters.scala 552:42:freechips.rocketchip.system.DefaultRV32Config.fir@19801.8]
  assign _T_372 = _T_371 | _T_104; // @[Parameters.scala 552:42:freechips.rocketchip.system.DefaultRV32Config.fir@19802.8]
  assign _T_373 = _T_372 | _T_124; // @[Parameters.scala 552:42:freechips.rocketchip.system.DefaultRV32Config.fir@19803.8]
  assign _T_374 = _T_117 & _T_373; // @[Parameters.scala 551:56:freechips.rocketchip.system.DefaultRV32Config.fir@19804.8]
  assign _T_383 = io_in_a_bits_size <= 4'h8; // @[Parameters.scala 93:42:freechips.rocketchip.system.DefaultRV32Config.fir@19813.8]
  assign _T_391 = _T_383 & _T_109; // @[Parameters.scala 551:56:freechips.rocketchip.system.DefaultRV32Config.fir@19821.8]
  assign _T_393 = _T_272 | _T_374; // @[Parameters.scala 553:30:freechips.rocketchip.system.DefaultRV32Config.fir@19823.8]
  assign _T_395 = _T_393 | _T_391; // @[Parameters.scala 553:30:freechips.rocketchip.system.DefaultRV32Config.fir@19825.8]
  assign _T_397 = _T_395 | reset; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@19827.8]
  assign _T_398 = ~_T_397; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@19828.8]
  assign _T_413 = io_in_a_bits_opcode == 3'h1; // @[Monitor.scala 119:25:freechips.rocketchip.system.DefaultRV32Config.fir@19864.6]
  assign _T_486 = ~_T_48; // @[Monitor.scala 124:33:freechips.rocketchip.system.DefaultRV32Config.fir@19954.8]
  assign _T_487 = io_in_a_bits_mask & _T_486; // @[Monitor.scala 124:31:freechips.rocketchip.system.DefaultRV32Config.fir@19955.8]
  assign _T_488 = _T_487 == 4'h0; // @[Monitor.scala 124:40:freechips.rocketchip.system.DefaultRV32Config.fir@19956.8]
  assign _T_490 = _T_488 | reset; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@19958.8]
  assign _T_491 = ~_T_490; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@19959.8]
  assign _T_492 = io_in_a_bits_opcode == 3'h2; // @[Monitor.scala 127:25:freechips.rocketchip.system.DefaultRV32Config.fir@19965.6]
  assign _T_494 = io_in_a_bits_size <= 4'h2; // @[Parameters.scala 93:42:freechips.rocketchip.system.DefaultRV32Config.fir@19968.8]
  assign _T_518 = _T_110 | _T_99; // @[Parameters.scala 552:42:freechips.rocketchip.system.DefaultRV32Config.fir@19992.8]
  assign _T_519 = _T_518 | _T_104; // @[Parameters.scala 552:42:freechips.rocketchip.system.DefaultRV32Config.fir@19993.8]
  assign _T_520 = _T_494 & _T_519; // @[Parameters.scala 551:56:freechips.rocketchip.system.DefaultRV32Config.fir@19994.8]
  assign _T_543 = _T_520 | reset; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@20017.8]
  assign _T_544 = ~_T_543; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@20018.8]
  assign _T_551 = io_in_a_bits_param <= 3'h4; // @[Bundles.scala 140:33:freechips.rocketchip.system.DefaultRV32Config.fir@20037.8]
  assign _T_553 = _T_551 | reset; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@20039.8]
  assign _T_554 = ~_T_553; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@20040.8]
  assign _T_559 = io_in_a_bits_opcode == 3'h3; // @[Monitor.scala 135:25:freechips.rocketchip.system.DefaultRV32Config.fir@20054.6]
  assign _T_618 = io_in_a_bits_param <= 3'h3; // @[Bundles.scala 147:30:freechips.rocketchip.system.DefaultRV32Config.fir@20126.8]
  assign _T_620 = _T_618 | reset; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@20128.8]
  assign _T_621 = ~_T_620; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@20129.8]
  assign _T_626 = io_in_a_bits_opcode == 3'h5; // @[Monitor.scala 143:25:freechips.rocketchip.system.DefaultRV32Config.fir@20143.6]
  assign _T_677 = _T_272 | reset; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@20195.8]
  assign _T_678 = ~_T_677; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@20196.8]
  assign _T_685 = io_in_a_bits_param <= 3'h1; // @[Bundles.scala 160:28:freechips.rocketchip.system.DefaultRV32Config.fir@20215.8]
  assign _T_687 = _T_685 | reset; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@20217.8]
  assign _T_688 = ~_T_687; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@20218.8]
  assign _T_697 = io_in_d_bits_opcode <= 3'h6; // @[Bundles.scala 44:24:freechips.rocketchip.system.DefaultRV32Config.fir@20242.6]
  assign _T_699 = _T_697 | reset; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@20244.6]
  assign _T_700 = ~_T_699; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@20245.6]
  assign _T_701 = io_in_d_bits_source == 2'h0; // @[Parameters.scala 47:9:freechips.rocketchip.system.DefaultRV32Config.fir@20250.6]
  assign _T_702 = io_in_d_bits_source == 2'h1; // @[Parameters.scala 47:9:freechips.rocketchip.system.DefaultRV32Config.fir@20251.6]
  assign _T_703 = io_in_d_bits_source == 2'h2; // @[Parameters.scala 47:9:freechips.rocketchip.system.DefaultRV32Config.fir@20252.6]
  assign _T_705 = _T_701 | _T_702; // @[Parameters.scala 924:46:freechips.rocketchip.system.DefaultRV32Config.fir@20258.6]
  assign _T_706 = _T_705 | _T_703; // @[Parameters.scala 924:46:freechips.rocketchip.system.DefaultRV32Config.fir@20259.6]
  assign _T_708 = io_in_d_bits_opcode == 3'h6; // @[Monitor.scala 307:25:freechips.rocketchip.system.DefaultRV32Config.fir@20261.6]
  assign _T_710 = _T_706 | reset; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@20264.8]
  assign _T_711 = ~_T_710; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@20265.8]
  assign _T_712 = io_in_d_bits_size >= 4'h2; // @[Monitor.scala 309:27:freechips.rocketchip.system.DefaultRV32Config.fir@20270.8]
  assign _T_714 = _T_712 | reset; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@20272.8]
  assign _T_715 = ~_T_714; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@20273.8]
  assign _T_716 = io_in_d_bits_param == 2'h0; // @[Monitor.scala 310:28:freechips.rocketchip.system.DefaultRV32Config.fir@20278.8]
  assign _T_718 = _T_716 | reset; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@20280.8]
  assign _T_719 = ~_T_718; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@20281.8]
  assign _T_720 = ~io_in_d_bits_corrupt; // @[Monitor.scala 311:15:freechips.rocketchip.system.DefaultRV32Config.fir@20286.8]
  assign _T_722 = _T_720 | reset; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@20288.8]
  assign _T_723 = ~_T_722; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@20289.8]
  assign _T_724 = ~io_in_d_bits_denied; // @[Monitor.scala 312:15:freechips.rocketchip.system.DefaultRV32Config.fir@20294.8]
  assign _T_726 = _T_724 | reset; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@20296.8]
  assign _T_727 = ~_T_726; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@20297.8]
  assign _T_728 = io_in_d_bits_opcode == 3'h4; // @[Monitor.scala 315:25:freechips.rocketchip.system.DefaultRV32Config.fir@20303.6]
  assign _T_739 = io_in_d_bits_param <= 2'h2; // @[Bundles.scala 104:26:freechips.rocketchip.system.DefaultRV32Config.fir@20327.8]
  assign _T_741 = _T_739 | reset; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@20329.8]
  assign _T_742 = ~_T_741; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@20330.8]
  assign _T_743 = io_in_d_bits_param != 2'h2; // @[Monitor.scala 320:28:freechips.rocketchip.system.DefaultRV32Config.fir@20335.8]
  assign _T_745 = _T_743 | reset; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@20337.8]
  assign _T_746 = ~_T_745; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@20338.8]
  assign _T_756 = io_in_d_bits_opcode == 3'h5; // @[Monitor.scala 325:25:freechips.rocketchip.system.DefaultRV32Config.fir@20361.6]
  assign _T_776 = _T_724 | io_in_d_bits_corrupt; // @[Monitor.scala 331:30:freechips.rocketchip.system.DefaultRV32Config.fir@20402.8]
  assign _T_778 = _T_776 | reset; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@20404.8]
  assign _T_779 = ~_T_778; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@20405.8]
  assign _T_785 = io_in_d_bits_opcode == 3'h0; // @[Monitor.scala 335:25:freechips.rocketchip.system.DefaultRV32Config.fir@20420.6]
  assign _T_802 = io_in_d_bits_opcode == 3'h1; // @[Monitor.scala 343:25:freechips.rocketchip.system.DefaultRV32Config.fir@20455.6]
  assign _T_820 = io_in_d_bits_opcode == 3'h2; // @[Monitor.scala 351:25:freechips.rocketchip.system.DefaultRV32Config.fir@20491.6]
  assign _T_844 = {1'b0,$signed(io_in_b_bits_address)}; // @[Parameters.scala 137:49:freechips.rocketchip.system.DefaultRV32Config.fir@20539.6]
  assign _T_870 = io_in_b_bits_address ^ 32'h3000; // @[Parameters.scala 137:31:freechips.rocketchip.system.DefaultRV32Config.fir@20569.6]
  assign _T_871 = {1'b0,$signed(_T_870)}; // @[Parameters.scala 137:49:freechips.rocketchip.system.DefaultRV32Config.fir@20570.6]
  assign _T_873 = $signed(_T_871) & -33'sh1000; // @[Parameters.scala 137:52:freechips.rocketchip.system.DefaultRV32Config.fir@20572.6]
  assign _T_874 = $signed(_T_873) == 33'sh0; // @[Parameters.scala 137:67:freechips.rocketchip.system.DefaultRV32Config.fir@20573.6]
  assign _T_875 = io_in_b_bits_address ^ 32'hc000000; // @[Parameters.scala 137:31:freechips.rocketchip.system.DefaultRV32Config.fir@20574.6]
  assign _T_876 = {1'b0,$signed(_T_875)}; // @[Parameters.scala 137:49:freechips.rocketchip.system.DefaultRV32Config.fir@20575.6]
  assign _T_878 = $signed(_T_876) & -33'sh4000000; // @[Parameters.scala 137:52:freechips.rocketchip.system.DefaultRV32Config.fir@20577.6]
  assign _T_879 = $signed(_T_878) == 33'sh0; // @[Parameters.scala 137:67:freechips.rocketchip.system.DefaultRV32Config.fir@20578.6]
  assign _T_880 = io_in_b_bits_address ^ 32'h2000000; // @[Parameters.scala 137:31:freechips.rocketchip.system.DefaultRV32Config.fir@20579.6]
  assign _T_881 = {1'b0,$signed(_T_880)}; // @[Parameters.scala 137:49:freechips.rocketchip.system.DefaultRV32Config.fir@20580.6]
  assign _T_883 = $signed(_T_881) & -33'sh10000; // @[Parameters.scala 137:52:freechips.rocketchip.system.DefaultRV32Config.fir@20582.6]
  assign _T_884 = $signed(_T_883) == 33'sh0; // @[Parameters.scala 137:67:freechips.rocketchip.system.DefaultRV32Config.fir@20583.6]
  assign _T_888 = $signed(_T_844) & -33'sh1000; // @[Parameters.scala 137:52:freechips.rocketchip.system.DefaultRV32Config.fir@20587.6]
  assign _T_889 = $signed(_T_888) == 33'sh0; // @[Parameters.scala 137:67:freechips.rocketchip.system.DefaultRV32Config.fir@20588.6]
  assign _T_890 = io_in_b_bits_address ^ 32'h10000; // @[Parameters.scala 137:31:freechips.rocketchip.system.DefaultRV32Config.fir@20589.6]
  assign _T_891 = {1'b0,$signed(_T_890)}; // @[Parameters.scala 137:49:freechips.rocketchip.system.DefaultRV32Config.fir@20590.6]
  assign _T_893 = $signed(_T_891) & -33'sh10000; // @[Parameters.scala 137:52:freechips.rocketchip.system.DefaultRV32Config.fir@20592.6]
  assign _T_894 = $signed(_T_893) == 33'sh0; // @[Parameters.scala 137:67:freechips.rocketchip.system.DefaultRV32Config.fir@20593.6]
  assign _T_895 = io_in_b_bits_address ^ 32'h80000000; // @[Parameters.scala 137:31:freechips.rocketchip.system.DefaultRV32Config.fir@20594.6]
  assign _T_896 = {1'b0,$signed(_T_895)}; // @[Parameters.scala 137:49:freechips.rocketchip.system.DefaultRV32Config.fir@20595.6]
  assign _T_898 = $signed(_T_896) & -33'sh10000000; // @[Parameters.scala 137:52:freechips.rocketchip.system.DefaultRV32Config.fir@20597.6]
  assign _T_899 = $signed(_T_898) == 33'sh0; // @[Parameters.scala 137:67:freechips.rocketchip.system.DefaultRV32Config.fir@20598.6]
  assign _T_900 = io_in_b_bits_address ^ 32'h60000000; // @[Parameters.scala 137:31:freechips.rocketchip.system.DefaultRV32Config.fir@20599.6]
  assign _T_901 = {1'b0,$signed(_T_900)}; // @[Parameters.scala 137:49:freechips.rocketchip.system.DefaultRV32Config.fir@20600.6]
  assign _T_903 = $signed(_T_901) & -33'sh20000000; // @[Parameters.scala 137:52:freechips.rocketchip.system.DefaultRV32Config.fir@20602.6]
  assign _T_904 = $signed(_T_903) == 33'sh0; // @[Parameters.scala 137:67:freechips.rocketchip.system.DefaultRV32Config.fir@20603.6]
  assign _T_906 = _T_874 | _T_879; // @[Parameters.scala 535:64:freechips.rocketchip.system.DefaultRV32Config.fir@20613.6]
  assign _T_907 = _T_906 | _T_884; // @[Parameters.scala 535:64:freechips.rocketchip.system.DefaultRV32Config.fir@20614.6]
  assign _T_908 = _T_907 | _T_889; // @[Parameters.scala 535:64:freechips.rocketchip.system.DefaultRV32Config.fir@20615.6]
  assign _T_909 = _T_908 | _T_894; // @[Parameters.scala 535:64:freechips.rocketchip.system.DefaultRV32Config.fir@20616.6]
  assign _T_910 = _T_909 | _T_899; // @[Parameters.scala 535:64:freechips.rocketchip.system.DefaultRV32Config.fir@20617.6]
  assign _T_911 = _T_910 | _T_904; // @[Parameters.scala 535:64:freechips.rocketchip.system.DefaultRV32Config.fir@20618.6]
  assign _T_916 = io_in_b_bits_address & 32'h3f; // @[Edges.scala 22:16:freechips.rocketchip.system.DefaultRV32Config.fir@20623.6]
  assign _T_917 = _T_916 == 32'h0; // @[Edges.scala 22:24:freechips.rocketchip.system.DefaultRV32Config.fir@20624.6]
  assign _T_978 = _T_911 | reset; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@20700.8]
  assign _T_979 = ~_T_978; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@20701.8]
  assign _T_984 = _T_917 | reset; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@20714.8]
  assign _T_985 = ~_T_984; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@20715.8]
  assign _T_986 = io_in_b_bits_param <= 2'h2; // @[Bundles.scala 104:26:freechips.rocketchip.system.DefaultRV32Config.fir@20720.8]
  assign _T_988 = _T_986 | reset; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@20722.8]
  assign _T_989 = ~_T_988; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@20723.8]
  assign _T_1134 = io_in_c_bits_source == 2'h0; // @[Parameters.scala 47:9:freechips.rocketchip.system.DefaultRV32Config.fir@21047.6]
  assign _T_1135 = io_in_c_bits_source == 2'h1; // @[Parameters.scala 47:9:freechips.rocketchip.system.DefaultRV32Config.fir@21048.6]
  assign _T_1136 = io_in_c_bits_source == 2'h2; // @[Parameters.scala 47:9:freechips.rocketchip.system.DefaultRV32Config.fir@21049.6]
  assign _T_1138 = _T_1134 | _T_1135; // @[Parameters.scala 924:46:freechips.rocketchip.system.DefaultRV32Config.fir@21055.6]
  assign _T_1139 = _T_1138 | _T_1136; // @[Parameters.scala 924:46:freechips.rocketchip.system.DefaultRV32Config.fir@21056.6]
  assign _T_1141 = 27'hfff << io_in_c_bits_size; // @[package.scala 207:77:freechips.rocketchip.system.DefaultRV32Config.fir@21058.6]
  assign _T_1143 = ~_T_1141[11:0]; // @[package.scala 207:46:freechips.rocketchip.system.DefaultRV32Config.fir@21060.6]
  assign _GEN_72 = {{20'd0}, _T_1143}; // @[Edges.scala 22:16:freechips.rocketchip.system.DefaultRV32Config.fir@21061.6]
  assign _T_1144 = io_in_c_bits_address & _GEN_72; // @[Edges.scala 22:16:freechips.rocketchip.system.DefaultRV32Config.fir@21061.6]
  assign _T_1145 = _T_1144 == 32'h0; // @[Edges.scala 22:24:freechips.rocketchip.system.DefaultRV32Config.fir@21062.6]
  assign _T_1146 = io_in_c_bits_address ^ 32'h3000; // @[Parameters.scala 137:31:freechips.rocketchip.system.DefaultRV32Config.fir@21063.6]
  assign _T_1147 = {1'b0,$signed(_T_1146)}; // @[Parameters.scala 137:49:freechips.rocketchip.system.DefaultRV32Config.fir@21064.6]
  assign _T_1149 = $signed(_T_1147) & -33'sh1000; // @[Parameters.scala 137:52:freechips.rocketchip.system.DefaultRV32Config.fir@21066.6]
  assign _T_1150 = $signed(_T_1149) == 33'sh0; // @[Parameters.scala 137:67:freechips.rocketchip.system.DefaultRV32Config.fir@21067.6]
  assign _T_1151 = io_in_c_bits_address ^ 32'hc000000; // @[Parameters.scala 137:31:freechips.rocketchip.system.DefaultRV32Config.fir@21068.6]
  assign _T_1152 = {1'b0,$signed(_T_1151)}; // @[Parameters.scala 137:49:freechips.rocketchip.system.DefaultRV32Config.fir@21069.6]
  assign _T_1154 = $signed(_T_1152) & -33'sh4000000; // @[Parameters.scala 137:52:freechips.rocketchip.system.DefaultRV32Config.fir@21071.6]
  assign _T_1155 = $signed(_T_1154) == 33'sh0; // @[Parameters.scala 137:67:freechips.rocketchip.system.DefaultRV32Config.fir@21072.6]
  assign _T_1156 = io_in_c_bits_address ^ 32'h2000000; // @[Parameters.scala 137:31:freechips.rocketchip.system.DefaultRV32Config.fir@21073.6]
  assign _T_1157 = {1'b0,$signed(_T_1156)}; // @[Parameters.scala 137:49:freechips.rocketchip.system.DefaultRV32Config.fir@21074.6]
  assign _T_1159 = $signed(_T_1157) & -33'sh10000; // @[Parameters.scala 137:52:freechips.rocketchip.system.DefaultRV32Config.fir@21076.6]
  assign _T_1160 = $signed(_T_1159) == 33'sh0; // @[Parameters.scala 137:67:freechips.rocketchip.system.DefaultRV32Config.fir@21077.6]
  assign _T_1162 = {1'b0,$signed(io_in_c_bits_address)}; // @[Parameters.scala 137:49:freechips.rocketchip.system.DefaultRV32Config.fir@21079.6]
  assign _T_1164 = $signed(_T_1162) & -33'sh1000; // @[Parameters.scala 137:52:freechips.rocketchip.system.DefaultRV32Config.fir@21081.6]
  assign _T_1165 = $signed(_T_1164) == 33'sh0; // @[Parameters.scala 137:67:freechips.rocketchip.system.DefaultRV32Config.fir@21082.6]
  assign _T_1166 = io_in_c_bits_address ^ 32'h10000; // @[Parameters.scala 137:31:freechips.rocketchip.system.DefaultRV32Config.fir@21083.6]
  assign _T_1167 = {1'b0,$signed(_T_1166)}; // @[Parameters.scala 137:49:freechips.rocketchip.system.DefaultRV32Config.fir@21084.6]
  assign _T_1169 = $signed(_T_1167) & -33'sh10000; // @[Parameters.scala 137:52:freechips.rocketchip.system.DefaultRV32Config.fir@21086.6]
  assign _T_1170 = $signed(_T_1169) == 33'sh0; // @[Parameters.scala 137:67:freechips.rocketchip.system.DefaultRV32Config.fir@21087.6]
  assign _T_1171 = io_in_c_bits_address ^ 32'h80000000; // @[Parameters.scala 137:31:freechips.rocketchip.system.DefaultRV32Config.fir@21088.6]
  assign _T_1172 = {1'b0,$signed(_T_1171)}; // @[Parameters.scala 137:49:freechips.rocketchip.system.DefaultRV32Config.fir@21089.6]
  assign _T_1174 = $signed(_T_1172) & -33'sh10000000; // @[Parameters.scala 137:52:freechips.rocketchip.system.DefaultRV32Config.fir@21091.6]
  assign _T_1175 = $signed(_T_1174) == 33'sh0; // @[Parameters.scala 137:67:freechips.rocketchip.system.DefaultRV32Config.fir@21092.6]
  assign _T_1176 = io_in_c_bits_address ^ 32'h60000000; // @[Parameters.scala 137:31:freechips.rocketchip.system.DefaultRV32Config.fir@21093.6]
  assign _T_1177 = {1'b0,$signed(_T_1176)}; // @[Parameters.scala 137:49:freechips.rocketchip.system.DefaultRV32Config.fir@21094.6]
  assign _T_1179 = $signed(_T_1177) & -33'sh20000000; // @[Parameters.scala 137:52:freechips.rocketchip.system.DefaultRV32Config.fir@21096.6]
  assign _T_1180 = $signed(_T_1179) == 33'sh0; // @[Parameters.scala 137:67:freechips.rocketchip.system.DefaultRV32Config.fir@21097.6]
  assign _T_1182 = _T_1150 | _T_1155; // @[Parameters.scala 535:64:freechips.rocketchip.system.DefaultRV32Config.fir@21107.6]
  assign _T_1183 = _T_1182 | _T_1160; // @[Parameters.scala 535:64:freechips.rocketchip.system.DefaultRV32Config.fir@21108.6]
  assign _T_1184 = _T_1183 | _T_1165; // @[Parameters.scala 535:64:freechips.rocketchip.system.DefaultRV32Config.fir@21109.6]
  assign _T_1185 = _T_1184 | _T_1170; // @[Parameters.scala 535:64:freechips.rocketchip.system.DefaultRV32Config.fir@21110.6]
  assign _T_1186 = _T_1185 | _T_1175; // @[Parameters.scala 535:64:freechips.rocketchip.system.DefaultRV32Config.fir@21111.6]
  assign _T_1187 = _T_1186 | _T_1180; // @[Parameters.scala 535:64:freechips.rocketchip.system.DefaultRV32Config.fir@21112.6]
  assign _T_1217 = io_in_c_bits_opcode == 3'h4; // @[Monitor.scala 239:25:freechips.rocketchip.system.DefaultRV32Config.fir@21146.6]
  assign _T_1219 = _T_1187 | reset; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@21149.8]
  assign _T_1220 = ~_T_1219; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@21150.8]
  assign _T_1222 = _T_1139 | reset; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@21156.8]
  assign _T_1223 = ~_T_1222; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@21157.8]
  assign _T_1224 = io_in_c_bits_size >= 4'h2; // @[Monitor.scala 242:30:freechips.rocketchip.system.DefaultRV32Config.fir@21162.8]
  assign _T_1226 = _T_1224 | reset; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@21164.8]
  assign _T_1227 = ~_T_1226; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@21165.8]
  assign _T_1229 = _T_1145 | reset; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@21171.8]
  assign _T_1230 = ~_T_1229; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@21172.8]
  assign _T_1231 = io_in_c_bits_param <= 3'h5; // @[Bundles.scala 122:29:freechips.rocketchip.system.DefaultRV32Config.fir@21177.8]
  assign _T_1233 = _T_1231 | reset; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@21179.8]
  assign _T_1234 = ~_T_1233; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@21180.8]
  assign _T_1235 = ~io_in_c_bits_corrupt; // @[Monitor.scala 245:18:freechips.rocketchip.system.DefaultRV32Config.fir@21185.8]
  assign _T_1237 = _T_1235 | reset; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@21187.8]
  assign _T_1238 = ~_T_1237; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@21188.8]
  assign _T_1239 = io_in_c_bits_opcode == 3'h5; // @[Monitor.scala 248:25:freechips.rocketchip.system.DefaultRV32Config.fir@21194.6]
  assign _T_1257 = io_in_c_bits_opcode == 3'h6; // @[Monitor.scala 256:25:freechips.rocketchip.system.DefaultRV32Config.fir@21234.6]
  assign _T_1296 = io_in_c_bits_size <= 4'h6; // @[Parameters.scala 93:42:freechips.rocketchip.system.DefaultRV32Config.fir@21274.8]
  assign _T_1304 = _T_1296 & _T_1175; // @[Parameters.scala 551:56:freechips.rocketchip.system.DefaultRV32Config.fir@21282.8]
  assign _T_1308 = _T_1304 | reset; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@21286.8]
  assign _T_1309 = ~_T_1308; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@21287.8]
  assign _T_1314 = 4'h6 == io_in_c_bits_size; // @[Parameters.scala 92:48:freechips.rocketchip.system.DefaultRV32Config.fir@21300.8]
  assign _T_1315 = _T_1134 & _T_1314; // @[Mux.scala 27:72:freechips.rocketchip.system.DefaultRV32Config.fir@21301.8]
  assign _T_1322 = _T_1315 | reset; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@21309.8]
  assign _T_1323 = ~_T_1322; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@21310.8]
  assign _T_1334 = io_in_c_bits_param <= 3'h2; // @[Bundles.scala 116:29:freechips.rocketchip.system.DefaultRV32Config.fir@21337.8]
  assign _T_1336 = _T_1334 | reset; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@21339.8]
  assign _T_1337 = ~_T_1336; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@21340.8]
  assign _T_1342 = io_in_c_bits_opcode == 3'h7; // @[Monitor.scala 266:25:freechips.rocketchip.system.DefaultRV32Config.fir@21354.6]
  assign _T_1423 = io_in_c_bits_opcode == 3'h0; // @[Monitor.scala 275:25:freechips.rocketchip.system.DefaultRV32Config.fir@21466.6]
  assign _T_1433 = io_in_c_bits_param == 3'h0; // @[Monitor.scala 279:31:freechips.rocketchip.system.DefaultRV32Config.fir@21489.8]
  assign _T_1435 = _T_1433 | reset; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@21491.8]
  assign _T_1436 = ~_T_1435; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@21492.8]
  assign _T_1441 = io_in_c_bits_opcode == 3'h1; // @[Monitor.scala 283:25:freechips.rocketchip.system.DefaultRV32Config.fir@21506.6]
  assign _T_1455 = io_in_c_bits_opcode == 3'h2; // @[Monitor.scala 290:25:freechips.rocketchip.system.DefaultRV32Config.fir@21538.6]
  assign _T_1477 = io_in_a_ready & io_in_a_valid; // @[Decoupled.scala 40:37:freechips.rocketchip.system.DefaultRV32Config.fir@21589.4]
  assign _T_1484 = ~io_in_a_bits_opcode[2]; // @[Edges.scala 93:28:freechips.rocketchip.system.DefaultRV32Config.fir@21596.4]
  assign _T_1488 = _T_1486 - 10'h1; // @[Edges.scala 231:28:freechips.rocketchip.system.DefaultRV32Config.fir@21600.4]
  assign _T_1489 = _T_1486 == 10'h0; // @[Edges.scala 232:25:freechips.rocketchip.system.DefaultRV32Config.fir@21601.4]
  assign _T_1502 = ~_T_1489; // @[Monitor.scala 386:22:freechips.rocketchip.system.DefaultRV32Config.fir@21617.4]
  assign _T_1503 = io_in_a_valid & _T_1502; // @[Monitor.scala 386:19:freechips.rocketchip.system.DefaultRV32Config.fir@21618.4]
  assign _T_1504 = io_in_a_bits_opcode == _T_1497; // @[Monitor.scala 387:32:freechips.rocketchip.system.DefaultRV32Config.fir@21620.6]
  assign _T_1506 = _T_1504 | reset; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@21622.6]
  assign _T_1507 = ~_T_1506; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@21623.6]
  assign _T_1508 = io_in_a_bits_param == _T_1498; // @[Monitor.scala 388:32:freechips.rocketchip.system.DefaultRV32Config.fir@21628.6]
  assign _T_1510 = _T_1508 | reset; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@21630.6]
  assign _T_1511 = ~_T_1510; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@21631.6]
  assign _T_1512 = io_in_a_bits_size == _T_1499; // @[Monitor.scala 389:32:freechips.rocketchip.system.DefaultRV32Config.fir@21636.6]
  assign _T_1514 = _T_1512 | reset; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@21638.6]
  assign _T_1515 = ~_T_1514; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@21639.6]
  assign _T_1516 = io_in_a_bits_source == _T_1500; // @[Monitor.scala 390:32:freechips.rocketchip.system.DefaultRV32Config.fir@21644.6]
  assign _T_1518 = _T_1516 | reset; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@21646.6]
  assign _T_1519 = ~_T_1518; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@21647.6]
  assign _T_1520 = io_in_a_bits_address == _T_1501; // @[Monitor.scala 391:32:freechips.rocketchip.system.DefaultRV32Config.fir@21652.6]
  assign _T_1522 = _T_1520 | reset; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@21654.6]
  assign _T_1523 = ~_T_1522; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@21655.6]
  assign _T_1525 = _T_1477 & _T_1489; // @[Monitor.scala 393:20:freechips.rocketchip.system.DefaultRV32Config.fir@21662.4]
  assign _T_1526 = io_in_d_ready & io_in_d_valid; // @[Decoupled.scala 40:37:freechips.rocketchip.system.DefaultRV32Config.fir@21670.4]
  assign _T_1528 = 27'hfff << io_in_d_bits_size; // @[package.scala 207:77:freechips.rocketchip.system.DefaultRV32Config.fir@21672.4]
  assign _T_1530 = ~_T_1528[11:0]; // @[package.scala 207:46:freechips.rocketchip.system.DefaultRV32Config.fir@21674.4]
  assign _T_1536 = _T_1534 - 10'h1; // @[Edges.scala 231:28:freechips.rocketchip.system.DefaultRV32Config.fir@21680.4]
  assign _T_1537 = _T_1534 == 10'h0; // @[Edges.scala 232:25:freechips.rocketchip.system.DefaultRV32Config.fir@21681.4]
  assign _T_1551 = ~_T_1537; // @[Monitor.scala 538:22:freechips.rocketchip.system.DefaultRV32Config.fir@21698.4]
  assign _T_1552 = io_in_d_valid & _T_1551; // @[Monitor.scala 538:19:freechips.rocketchip.system.DefaultRV32Config.fir@21699.4]
  assign _T_1553 = io_in_d_bits_opcode == _T_1545; // @[Monitor.scala 539:29:freechips.rocketchip.system.DefaultRV32Config.fir@21701.6]
  assign _T_1555 = _T_1553 | reset; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@21703.6]
  assign _T_1556 = ~_T_1555; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@21704.6]
  assign _T_1557 = io_in_d_bits_param == _T_1546; // @[Monitor.scala 540:29:freechips.rocketchip.system.DefaultRV32Config.fir@21709.6]
  assign _T_1559 = _T_1557 | reset; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@21711.6]
  assign _T_1560 = ~_T_1559; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@21712.6]
  assign _T_1561 = io_in_d_bits_size == _T_1547; // @[Monitor.scala 541:29:freechips.rocketchip.system.DefaultRV32Config.fir@21717.6]
  assign _T_1563 = _T_1561 | reset; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@21719.6]
  assign _T_1564 = ~_T_1563; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@21720.6]
  assign _T_1565 = io_in_d_bits_source == _T_1548; // @[Monitor.scala 542:29:freechips.rocketchip.system.DefaultRV32Config.fir@21725.6]
  assign _T_1567 = _T_1565 | reset; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@21727.6]
  assign _T_1568 = ~_T_1567; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@21728.6]
  assign _T_1569 = io_in_d_bits_sink == _T_1549; // @[Monitor.scala 543:29:freechips.rocketchip.system.DefaultRV32Config.fir@21733.6]
  assign _T_1571 = _T_1569 | reset; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@21735.6]
  assign _T_1572 = ~_T_1571; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@21736.6]
  assign _T_1573 = io_in_d_bits_denied == _T_1550; // @[Monitor.scala 544:29:freechips.rocketchip.system.DefaultRV32Config.fir@21741.6]
  assign _T_1575 = _T_1573 | reset; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@21743.6]
  assign _T_1576 = ~_T_1575; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@21744.6]
  assign _T_1578 = _T_1526 & _T_1537; // @[Monitor.scala 546:20:freechips.rocketchip.system.DefaultRV32Config.fir@21751.4]
  assign _T_1579 = io_in_b_ready & io_in_b_valid; // @[Decoupled.scala 40:37:freechips.rocketchip.system.DefaultRV32Config.fir@21760.4]
  assign _T_1590 = _T_1588 - 10'h1; // @[Edges.scala 231:28:freechips.rocketchip.system.DefaultRV32Config.fir@21771.4]
  assign _T_1591 = _T_1588 == 10'h0; // @[Edges.scala 232:25:freechips.rocketchip.system.DefaultRV32Config.fir@21772.4]
  assign _T_1604 = ~_T_1591; // @[Monitor.scala 409:22:freechips.rocketchip.system.DefaultRV32Config.fir@21788.4]
  assign _T_1605 = io_in_b_valid & _T_1604; // @[Monitor.scala 409:19:freechips.rocketchip.system.DefaultRV32Config.fir@21789.4]
  assign _T_1610 = io_in_b_bits_param == _T_1600; // @[Monitor.scala 411:32:freechips.rocketchip.system.DefaultRV32Config.fir@21799.6]
  assign _T_1612 = _T_1610 | reset; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@21801.6]
  assign _T_1613 = ~_T_1612; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@21802.6]
  assign _T_1622 = io_in_b_bits_address == _T_1603; // @[Monitor.scala 414:32:freechips.rocketchip.system.DefaultRV32Config.fir@21823.6]
  assign _T_1624 = _T_1622 | reset; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@21825.6]
  assign _T_1625 = ~_T_1624; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@21826.6]
  assign _T_1627 = _T_1579 & _T_1591; // @[Monitor.scala 416:20:freechips.rocketchip.system.DefaultRV32Config.fir@21833.4]
  assign _T_1628 = io_in_c_ready & io_in_c_valid; // @[Decoupled.scala 40:37:freechips.rocketchip.system.DefaultRV32Config.fir@21841.4]
  assign _T_1638 = _T_1636 - 10'h1; // @[Edges.scala 231:28:freechips.rocketchip.system.DefaultRV32Config.fir@21851.4]
  assign _T_1639 = _T_1636 == 10'h0; // @[Edges.scala 232:25:freechips.rocketchip.system.DefaultRV32Config.fir@21852.4]
  assign _T_1652 = ~_T_1639; // @[Monitor.scala 514:22:freechips.rocketchip.system.DefaultRV32Config.fir@21868.4]
  assign _T_1653 = io_in_c_valid & _T_1652; // @[Monitor.scala 514:19:freechips.rocketchip.system.DefaultRV32Config.fir@21869.4]
  assign _T_1654 = io_in_c_bits_opcode == _T_1647; // @[Monitor.scala 515:32:freechips.rocketchip.system.DefaultRV32Config.fir@21871.6]
  assign _T_1656 = _T_1654 | reset; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@21873.6]
  assign _T_1657 = ~_T_1656; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@21874.6]
  assign _T_1658 = io_in_c_bits_param == _T_1648; // @[Monitor.scala 516:32:freechips.rocketchip.system.DefaultRV32Config.fir@21879.6]
  assign _T_1660 = _T_1658 | reset; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@21881.6]
  assign _T_1661 = ~_T_1660; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@21882.6]
  assign _T_1662 = io_in_c_bits_size == _T_1649; // @[Monitor.scala 517:32:freechips.rocketchip.system.DefaultRV32Config.fir@21887.6]
  assign _T_1664 = _T_1662 | reset; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@21889.6]
  assign _T_1665 = ~_T_1664; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@21890.6]
  assign _T_1666 = io_in_c_bits_source == _T_1650; // @[Monitor.scala 518:32:freechips.rocketchip.system.DefaultRV32Config.fir@21895.6]
  assign _T_1668 = _T_1666 | reset; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@21897.6]
  assign _T_1669 = ~_T_1668; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@21898.6]
  assign _T_1670 = io_in_c_bits_address == _T_1651; // @[Monitor.scala 519:32:freechips.rocketchip.system.DefaultRV32Config.fir@21903.6]
  assign _T_1672 = _T_1670 | reset; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@21905.6]
  assign _T_1673 = ~_T_1672; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@21906.6]
  assign _T_1675 = _T_1628 & _T_1639; // @[Monitor.scala 521:20:freechips.rocketchip.system.DefaultRV32Config.fir@21913.4]
  assign _T_1687 = _T_1685 - 10'h1; // @[Edges.scala 231:28:freechips.rocketchip.system.DefaultRV32Config.fir@21935.4]
  assign a_first = _T_1685 == 10'h0; // @[Edges.scala 232:25:freechips.rocketchip.system.DefaultRV32Config.fir@21936.4]
  assign _T_1705 = _T_1703 - 10'h1; // @[Edges.scala 231:28:freechips.rocketchip.system.DefaultRV32Config.fir@21957.4]
  assign d_first = _T_1703 == 10'h0; // @[Edges.scala 232:25:freechips.rocketchip.system.DefaultRV32Config.fir@21958.4]
  assign _GEN_73 = {io_in_d_bits_source, 2'h0}; // @[Monitor.scala 629:69:freechips.rocketchip.system.DefaultRV32Config.fir@21977.4]
  assign _T_1713 = {{1'd0}, _GEN_73}; // @[Monitor.scala 629:69:freechips.rocketchip.system.DefaultRV32Config.fir@21977.4]
  assign _T_1714 = inflight_opcodes >> _T_1713; // @[Monitor.scala 629:44:freechips.rocketchip.system.DefaultRV32Config.fir@21978.4]
  assign _T_1718 = 16'h10 - 16'h1; // @[Monitor.scala 606:57:freechips.rocketchip.system.DefaultRV32Config.fir@21982.4]
  assign _GEN_74 = {{4'd0}, _T_1714}; // @[Monitor.scala 629:97:freechips.rocketchip.system.DefaultRV32Config.fir@21983.4]
  assign _T_1719 = _GEN_74 & _T_1718; // @[Monitor.scala 629:97:freechips.rocketchip.system.DefaultRV32Config.fir@21983.4]
  assign _T_1720 = {{1'd0}, _T_1719[15:1]}; // @[Monitor.scala 629:152:freechips.rocketchip.system.DefaultRV32Config.fir@21984.4]
  assign _T_1721 = {io_in_d_bits_source, 3'h0}; // @[Monitor.scala 633:65:freechips.rocketchip.system.DefaultRV32Config.fir@21988.4]
  assign _T_1722 = inflight_sizes >> _T_1721; // @[Monitor.scala 633:40:freechips.rocketchip.system.DefaultRV32Config.fir@21989.4]
  assign _T_1726 = 16'h100 - 16'h1; // @[Monitor.scala 606:57:freechips.rocketchip.system.DefaultRV32Config.fir@21993.4]
  assign _GEN_76 = {{8'd0}, _T_1726}; // @[Monitor.scala 633:91:freechips.rocketchip.system.DefaultRV32Config.fir@21994.4]
  assign _T_1727 = _T_1722 & _GEN_76; // @[Monitor.scala 633:91:freechips.rocketchip.system.DefaultRV32Config.fir@21994.4]
  assign _T_1728 = {{1'd0}, _T_1727[23:1]}; // @[Monitor.scala 633:144:freechips.rocketchip.system.DefaultRV32Config.fir@21995.4]
  assign _T_1732 = _T_1477 & a_first; // @[Monitor.scala 643:27:freechips.rocketchip.system.DefaultRV32Config.fir@22020.4]
  assign _T_1734 = 4'h1 << io_in_a_bits_source; // @[OneHot.scala 58:35:freechips.rocketchip.system.DefaultRV32Config.fir@22023.6]
  assign _T_1735 = {io_in_a_bits_opcode, 1'h0}; // @[Monitor.scala 645:53:freechips.rocketchip.system.DefaultRV32Config.fir@22025.6]
  assign _T_1736 = _T_1735 | 4'h1; // @[Monitor.scala 645:61:freechips.rocketchip.system.DefaultRV32Config.fir@22026.6]
  assign _T_1737 = {io_in_a_bits_size, 1'h0}; // @[Monitor.scala 646:49:freechips.rocketchip.system.DefaultRV32Config.fir@22028.6]
  assign _T_1738 = _T_1737 | 5'h1; // @[Monitor.scala 646:57:freechips.rocketchip.system.DefaultRV32Config.fir@22029.6]
  assign _GEN_78 = {io_in_a_bits_source, 2'h0}; // @[Monitor.scala 647:72:freechips.rocketchip.system.DefaultRV32Config.fir@22031.6]
  assign _T_1739 = {{1'd0}, _GEN_78}; // @[Monitor.scala 647:72:freechips.rocketchip.system.DefaultRV32Config.fir@22031.6]
  assign a_opcodes_set_interm = _T_1732 ? _T_1736 : 4'h0; // @[Monitor.scala 643:72:freechips.rocketchip.system.DefaultRV32Config.fir@22022.4]
  assign _GEN_79 = {{31'd0}, a_opcodes_set_interm}; // @[Monitor.scala 647:47:freechips.rocketchip.system.DefaultRV32Config.fir@22032.6]
  assign _T_1740 = _GEN_79 << _T_1739; // @[Monitor.scala 647:47:freechips.rocketchip.system.DefaultRV32Config.fir@22032.6]
  assign _T_1741 = {io_in_a_bits_source, 3'h0}; // @[Monitor.scala 648:68:freechips.rocketchip.system.DefaultRV32Config.fir@22034.6]
  assign a_sizes_set_interm = _T_1732 ? _T_1738 : 5'h0; // @[Monitor.scala 643:72:freechips.rocketchip.system.DefaultRV32Config.fir@22022.4]
  assign _GEN_80 = {{31'd0}, a_sizes_set_interm}; // @[Monitor.scala 648:43:freechips.rocketchip.system.DefaultRV32Config.fir@22035.6]
  assign _T_1742 = _GEN_80 << _T_1741; // @[Monitor.scala 648:43:freechips.rocketchip.system.DefaultRV32Config.fir@22035.6]
  assign _T_1743 = inflight >> io_in_a_bits_source; // @[Monitor.scala 649:26:freechips.rocketchip.system.DefaultRV32Config.fir@22037.6]
  assign _T_1745 = ~_T_1743[0]; // @[Monitor.scala 649:17:freechips.rocketchip.system.DefaultRV32Config.fir@22039.6]
  assign _T_1747 = _T_1745 | reset; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@22041.6]
  assign _T_1748 = ~_T_1747; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@22042.6]
  assign _GEN_27 = _T_1732 ? _T_1734 : 4'h0; // @[Monitor.scala 643:72:freechips.rocketchip.system.DefaultRV32Config.fir@22022.4]
  assign _GEN_30 = _T_1732 ? _T_1740 : 35'h0; // @[Monitor.scala 643:72:freechips.rocketchip.system.DefaultRV32Config.fir@22022.4]
  assign _GEN_31 = _T_1732 ? _T_1742 : 36'h0; // @[Monitor.scala 643:72:freechips.rocketchip.system.DefaultRV32Config.fir@22022.4]
  assign _T_1751 = _T_1526 & d_first; // @[Monitor.scala 660:27:freechips.rocketchip.system.DefaultRV32Config.fir@22056.4]
  assign _T_1753 = ~_T_708; // @[Monitor.scala 660:75:freechips.rocketchip.system.DefaultRV32Config.fir@22058.4]
  assign _T_1754 = _T_1751 & _T_1753; // @[Monitor.scala 660:72:freechips.rocketchip.system.DefaultRV32Config.fir@22059.4]
  assign _T_1755 = 4'h1 << io_in_d_bits_source; // @[OneHot.scala 58:35:freechips.rocketchip.system.DefaultRV32Config.fir@22061.6]
  assign _GEN_82 = {{31'd0}, _T_1718}; // @[Monitor.scala 662:76:freechips.rocketchip.system.DefaultRV32Config.fir@22068.6]
  assign _T_1761 = _GEN_82 << _T_1713; // @[Monitor.scala 662:76:freechips.rocketchip.system.DefaultRV32Config.fir@22068.6]
  assign _GEN_83 = {{31'd0}, _T_1726}; // @[Monitor.scala 663:72:freechips.rocketchip.system.DefaultRV32Config.fir@22075.6]
  assign _T_1767 = _GEN_83 << _T_1721; // @[Monitor.scala 663:72:freechips.rocketchip.system.DefaultRV32Config.fir@22075.6]
  assign _GEN_32 = _T_1754 ? _T_1755 : 4'h0; // @[Monitor.scala 660:91:freechips.rocketchip.system.DefaultRV32Config.fir@22060.4]
  assign _GEN_33 = _T_1754 ? _T_1761 : 47'h0; // @[Monitor.scala 660:91:freechips.rocketchip.system.DefaultRV32Config.fir@22060.4]
  assign _GEN_34 = _T_1754 ? _T_1767 : 47'h0; // @[Monitor.scala 660:91:freechips.rocketchip.system.DefaultRV32Config.fir@22060.4]
  assign _T_1768 = io_in_d_valid & d_first; // @[Monitor.scala 665:26:freechips.rocketchip.system.DefaultRV32Config.fir@22078.4]
  assign _T_1771 = _T_1768 & _T_1753; // @[Monitor.scala 665:71:freechips.rocketchip.system.DefaultRV32Config.fir@22081.4]
  assign _T_1772 = inflight >> io_in_d_bits_source; // @[Monitor.scala 666:25:freechips.rocketchip.system.DefaultRV32Config.fir@22083.6]
  assign _T_1774 = io_in_a_bits_source == io_in_d_bits_source; // @[Monitor.scala 666:93:freechips.rocketchip.system.DefaultRV32Config.fir@22085.6]
  assign _T_1775 = io_in_a_valid & _T_1774; // @[Monitor.scala 666:68:freechips.rocketchip.system.DefaultRV32Config.fir@22086.6]
  assign _T_1776 = io_in_a_bits_size == io_in_d_bits_size; // @[Monitor.scala 666:142:freechips.rocketchip.system.DefaultRV32Config.fir@22087.6]
  assign _T_1777 = _T_1775 & _T_1776; // @[Monitor.scala 666:119:freechips.rocketchip.system.DefaultRV32Config.fir@22088.6]
  assign _T_1778 = _T_1777 & a_first; // @[Monitor.scala 666:166:freechips.rocketchip.system.DefaultRV32Config.fir@22089.6]
  assign _T_1779 = _T_1772[0] | _T_1778; // @[Monitor.scala 666:49:freechips.rocketchip.system.DefaultRV32Config.fir@22090.6]
  assign _T_1781 = _T_1779 | reset; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@22092.6]
  assign _T_1782 = ~_T_1781; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@22093.6]
  assign a_opcode_lookup = _T_1720[3:0]; // @[:freechips.rocketchip.system.DefaultRV32Config.fir@21975.4 :freechips.rocketchip.system.DefaultRV32Config.fir@21976.4 Monitor.scala 629:21:freechips.rocketchip.system.DefaultRV32Config.fir@21985.4]
  assign _GEN_37 = 3'h2 == a_opcode_lookup[2:0] ? 3'h1 : 3'h0; // @[Monitor.scala 667:37:freechips.rocketchip.system.DefaultRV32Config.fir@22099.6]
  assign _GEN_38 = 3'h3 == a_opcode_lookup[2:0] ? 3'h1 : _GEN_37; // @[Monitor.scala 667:37:freechips.rocketchip.system.DefaultRV32Config.fir@22099.6]
  assign _GEN_39 = 3'h4 == a_opcode_lookup[2:0] ? 3'h1 : _GEN_38; // @[Monitor.scala 667:37:freechips.rocketchip.system.DefaultRV32Config.fir@22099.6]
  assign _GEN_40 = 3'h5 == a_opcode_lookup[2:0] ? 3'h2 : _GEN_39; // @[Monitor.scala 667:37:freechips.rocketchip.system.DefaultRV32Config.fir@22099.6]
  assign _GEN_41 = 3'h6 == a_opcode_lookup[2:0] ? 3'h4 : _GEN_40; // @[Monitor.scala 667:37:freechips.rocketchip.system.DefaultRV32Config.fir@22099.6]
  assign _GEN_42 = 3'h7 == a_opcode_lookup[2:0] ? 3'h4 : _GEN_41; // @[Monitor.scala 667:37:freechips.rocketchip.system.DefaultRV32Config.fir@22099.6]
  assign _T_1784 = io_in_d_bits_opcode == _GEN_42; // @[Monitor.scala 667:37:freechips.rocketchip.system.DefaultRV32Config.fir@22099.6]
  assign _GEN_49 = 3'h6 == a_opcode_lookup[2:0] ? 3'h5 : _GEN_40; // @[Monitor.scala 667:96:freechips.rocketchip.system.DefaultRV32Config.fir@22101.6]
  assign _GEN_50 = 3'h7 == a_opcode_lookup[2:0] ? 3'h4 : _GEN_49; // @[Monitor.scala 667:96:freechips.rocketchip.system.DefaultRV32Config.fir@22101.6]
  assign _T_1786 = io_in_d_bits_opcode == _GEN_50; // @[Monitor.scala 667:96:freechips.rocketchip.system.DefaultRV32Config.fir@22101.6]
  assign _T_1787 = _T_1784 | _T_1786; // @[Monitor.scala 667:71:freechips.rocketchip.system.DefaultRV32Config.fir@22102.6]
  assign _GEN_53 = 3'h2 == io_in_a_bits_opcode ? 3'h1 : 3'h0; // @[Monitor.scala 668:60:freechips.rocketchip.system.DefaultRV32Config.fir@22103.6]
  assign _GEN_54 = 3'h3 == io_in_a_bits_opcode ? 3'h1 : _GEN_53; // @[Monitor.scala 668:60:freechips.rocketchip.system.DefaultRV32Config.fir@22103.6]
  assign _GEN_55 = 3'h4 == io_in_a_bits_opcode ? 3'h1 : _GEN_54; // @[Monitor.scala 668:60:freechips.rocketchip.system.DefaultRV32Config.fir@22103.6]
  assign _GEN_56 = 3'h5 == io_in_a_bits_opcode ? 3'h2 : _GEN_55; // @[Monitor.scala 668:60:freechips.rocketchip.system.DefaultRV32Config.fir@22103.6]
  assign _GEN_57 = 3'h6 == io_in_a_bits_opcode ? 3'h4 : _GEN_56; // @[Monitor.scala 668:60:freechips.rocketchip.system.DefaultRV32Config.fir@22103.6]
  assign _GEN_58 = 3'h7 == io_in_a_bits_opcode ? 3'h4 : _GEN_57; // @[Monitor.scala 668:60:freechips.rocketchip.system.DefaultRV32Config.fir@22103.6]
  assign _T_1788 = io_in_d_bits_opcode == _GEN_58; // @[Monitor.scala 668:60:freechips.rocketchip.system.DefaultRV32Config.fir@22103.6]
  assign _GEN_65 = 3'h6 == io_in_a_bits_opcode ? 3'h5 : _GEN_56; // @[Monitor.scala 668:124:freechips.rocketchip.system.DefaultRV32Config.fir@22104.6]
  assign _GEN_66 = 3'h7 == io_in_a_bits_opcode ? 3'h4 : _GEN_65; // @[Monitor.scala 668:124:freechips.rocketchip.system.DefaultRV32Config.fir@22104.6]
  assign _T_1789 = io_in_d_bits_opcode == _GEN_66; // @[Monitor.scala 668:124:freechips.rocketchip.system.DefaultRV32Config.fir@22104.6]
  assign _T_1790 = _T_1788 | _T_1789; // @[Monitor.scala 668:99:freechips.rocketchip.system.DefaultRV32Config.fir@22105.6]
  assign _T_1791 = io_in_a_valid & _T_1790; // @[Monitor.scala 668:34:freechips.rocketchip.system.DefaultRV32Config.fir@22106.6]
  assign _T_1792 = _T_1787 | _T_1791; // @[Monitor.scala 668:15:freechips.rocketchip.system.DefaultRV32Config.fir@22107.6]
  assign _T_1794 = _T_1792 | reset; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@22109.6]
  assign _T_1795 = ~_T_1794; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@22110.6]
  assign a_size_lookup = _T_1728[7:0]; // @[:freechips.rocketchip.system.DefaultRV32Config.fir@21986.4 :freechips.rocketchip.system.DefaultRV32Config.fir@21987.4 Monitor.scala 633:19:freechips.rocketchip.system.DefaultRV32Config.fir@21996.4]
  assign _GEN_84 = {{4'd0}, io_in_d_bits_size}; // @[Monitor.scala 670:34:freechips.rocketchip.system.DefaultRV32Config.fir@22115.6]
  assign _T_1796 = _GEN_84 == a_size_lookup; // @[Monitor.scala 670:34:freechips.rocketchip.system.DefaultRV32Config.fir@22115.6]
  assign _T_1798 = io_in_a_valid & _T_1776; // @[Monitor.scala 670:72:freechips.rocketchip.system.DefaultRV32Config.fir@22117.6]
  assign _T_1799 = _T_1796 | _T_1798; // @[Monitor.scala 670:53:freechips.rocketchip.system.DefaultRV32Config.fir@22118.6]
  assign _T_1801 = _T_1799 | reset; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@22120.6]
  assign _T_1802 = ~_T_1801; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@22121.6]
  assign _T_1804 = _T_1768 & a_first; // @[Monitor.scala 672:36:freechips.rocketchip.system.DefaultRV32Config.fir@22128.4]
  assign _T_1805 = _T_1804 & io_in_a_valid; // @[Monitor.scala 672:47:freechips.rocketchip.system.DefaultRV32Config.fir@22129.4]
  assign _T_1807 = _T_1805 & _T_1774; // @[Monitor.scala 672:65:freechips.rocketchip.system.DefaultRV32Config.fir@22131.4]
  assign _T_1809 = _T_1807 & _T_1753; // @[Monitor.scala 672:116:freechips.rocketchip.system.DefaultRV32Config.fir@22133.4]
  assign _T_1810 = ~io_in_d_ready; // @[Monitor.scala 673:15:freechips.rocketchip.system.DefaultRV32Config.fir@22135.6]
  assign _T_1811 = _T_1810 | io_in_a_ready; // @[Monitor.scala 673:32:freechips.rocketchip.system.DefaultRV32Config.fir@22136.6]
  assign _T_1813 = _T_1811 | reset; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@22138.6]
  assign _T_1814 = ~_T_1813; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@22139.6]
  assign a_set = _GEN_27[2:0]; // @[:freechips.rocketchip.system.DefaultRV32Config.fir@21969.4 :freechips.rocketchip.system.DefaultRV32Config.fir@21970.4 Monitor.scala 644:13:freechips.rocketchip.system.DefaultRV32Config.fir@22024.6]
  assign d_clr = _GEN_32[2:0]; // @[:freechips.rocketchip.system.DefaultRV32Config.fir@22048.4 :freechips.rocketchip.system.DefaultRV32Config.fir@22049.4 Monitor.scala 661:13:freechips.rocketchip.system.DefaultRV32Config.fir@22062.6]
  assign _T_1815 = a_set != d_clr; // @[Monitor.scala 677:20:freechips.rocketchip.system.DefaultRV32Config.fir@22145.4]
  assign _T_1816 = |a_set; // @[Monitor.scala 677:40:freechips.rocketchip.system.DefaultRV32Config.fir@22146.4]
  assign _T_1817 = ~_T_1816; // @[Monitor.scala 677:33:freechips.rocketchip.system.DefaultRV32Config.fir@22147.4]
  assign _T_1818 = _T_1815 | _T_1817; // @[Monitor.scala 677:30:freechips.rocketchip.system.DefaultRV32Config.fir@22148.4]
  assign _T_1820 = _T_1818 | reset; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@22150.4]
  assign _T_1821 = ~_T_1820; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@22151.4]
  assign _T_1822 = inflight | a_set; // @[Monitor.scala 680:27:freechips.rocketchip.system.DefaultRV32Config.fir@22156.4]
  assign _T_1823 = ~d_clr; // @[Monitor.scala 680:38:freechips.rocketchip.system.DefaultRV32Config.fir@22157.4]
  assign _T_1824 = _T_1822 & _T_1823; // @[Monitor.scala 680:36:freechips.rocketchip.system.DefaultRV32Config.fir@22158.4]
  assign a_opcodes_set = _GEN_30[11:0]; // @[:freechips.rocketchip.system.DefaultRV32Config.fir@21971.4 :freechips.rocketchip.system.DefaultRV32Config.fir@21972.4 Monitor.scala 647:21:freechips.rocketchip.system.DefaultRV32Config.fir@22033.6]
  assign _T_1825 = inflight_opcodes | a_opcodes_set; // @[Monitor.scala 681:43:freechips.rocketchip.system.DefaultRV32Config.fir@22160.4]
  assign d_opcodes_clr = _GEN_33[11:0]; // @[:freechips.rocketchip.system.DefaultRV32Config.fir@22050.4 :freechips.rocketchip.system.DefaultRV32Config.fir@22051.4 Monitor.scala 662:21:freechips.rocketchip.system.DefaultRV32Config.fir@22069.6]
  assign _T_1826 = ~d_opcodes_clr; // @[Monitor.scala 681:62:freechips.rocketchip.system.DefaultRV32Config.fir@22161.4]
  assign _T_1827 = _T_1825 & _T_1826; // @[Monitor.scala 681:60:freechips.rocketchip.system.DefaultRV32Config.fir@22162.4]
  assign a_sizes_set = _GEN_31[23:0]; // @[:freechips.rocketchip.system.DefaultRV32Config.fir@21973.4 :freechips.rocketchip.system.DefaultRV32Config.fir@21974.4 Monitor.scala 648:19:freechips.rocketchip.system.DefaultRV32Config.fir@22036.6]
  assign _T_1828 = inflight_sizes | a_sizes_set; // @[Monitor.scala 682:39:freechips.rocketchip.system.DefaultRV32Config.fir@22164.4]
  assign d_sizes_clr = _GEN_34[23:0]; // @[:freechips.rocketchip.system.DefaultRV32Config.fir@22052.4 :freechips.rocketchip.system.DefaultRV32Config.fir@22053.4 Monitor.scala 663:19:freechips.rocketchip.system.DefaultRV32Config.fir@22076.6]
  assign _T_1829 = ~d_sizes_clr; // @[Monitor.scala 682:56:freechips.rocketchip.system.DefaultRV32Config.fir@22165.4]
  assign _T_1830 = _T_1828 & _T_1829; // @[Monitor.scala 682:54:freechips.rocketchip.system.DefaultRV32Config.fir@22166.4]
  assign _T_1832 = |inflight; // @[Monitor.scala 687:26:freechips.rocketchip.system.DefaultRV32Config.fir@22171.4]
  assign _T_1833 = ~_T_1832; // @[Monitor.scala 687:16:freechips.rocketchip.system.DefaultRV32Config.fir@22172.4]
  assign _T_1834 = plusarg_reader_out == 32'h0; // @[Monitor.scala 687:39:freechips.rocketchip.system.DefaultRV32Config.fir@22173.4]
  assign _T_1835 = _T_1833 | _T_1834; // @[Monitor.scala 687:30:freechips.rocketchip.system.DefaultRV32Config.fir@22174.4]
  assign _T_1836 = _T_1831 < plusarg_reader_out; // @[Monitor.scala 687:59:freechips.rocketchip.system.DefaultRV32Config.fir@22175.4]
  assign _T_1837 = _T_1835 | _T_1836; // @[Monitor.scala 687:47:freechips.rocketchip.system.DefaultRV32Config.fir@22176.4]
  assign _T_1839 = _T_1837 | reset; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@22178.4]
  assign _T_1840 = ~_T_1839; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@22179.4]
  assign _T_1842 = _T_1831 + 32'h1; // @[Monitor.scala 689:26:freechips.rocketchip.system.DefaultRV32Config.fir@22185.4]
  assign _T_1845 = _T_1477 | _T_1526; // @[Monitor.scala 690:27:freechips.rocketchip.system.DefaultRV32Config.fir@22189.4]
  assign _T_1857 = _T_1855 - 10'h1; // @[Edges.scala 231:28:freechips.rocketchip.system.DefaultRV32Config.fir@22204.4]
  assign _T_1858 = _T_1855 == 10'h0; // @[Edges.scala 232:25:freechips.rocketchip.system.DefaultRV32Config.fir@22205.4]
  assign _T_1868 = _T_1526 & _T_1858; // @[Monitor.scala 700:27:freechips.rocketchip.system.DefaultRV32Config.fir@22219.4]
  assign _T_1871 = ~io_in_d_bits_opcode[1]; // @[Edges.scala 72:43:freechips.rocketchip.system.DefaultRV32Config.fir@22222.4]
  assign _T_1872 = io_in_d_bits_opcode[2] & _T_1871; // @[Edges.scala 72:40:freechips.rocketchip.system.DefaultRV32Config.fir@22223.4]
  assign _T_1873 = _T_1868 & _T_1872; // @[Monitor.scala 700:38:freechips.rocketchip.system.DefaultRV32Config.fir@22224.4]
  assign _T_1874 = 4'h1 << io_in_d_bits_sink; // @[OneHot.scala 58:35:freechips.rocketchip.system.DefaultRV32Config.fir@22226.6]
  assign _T_1875 = _T_1846 >> io_in_d_bits_sink; // @[Monitor.scala 702:23:freechips.rocketchip.system.DefaultRV32Config.fir@22228.6]
  assign _T_1877 = ~_T_1875[0]; // @[Monitor.scala 702:14:freechips.rocketchip.system.DefaultRV32Config.fir@22230.6]
  assign _T_1879 = _T_1877 | reset; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@22232.6]
  assign _T_1880 = ~_T_1879; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@22233.6]
  assign _GEN_69 = _T_1873 ? _T_1874 : 4'h0; // @[Monitor.scala 700:72:freechips.rocketchip.system.DefaultRV32Config.fir@22225.4]
  assign _T_1885 = 4'h1 << io_in_e_bits_sink; // @[OneHot.scala 58:35:freechips.rocketchip.system.DefaultRV32Config.fir@22245.6]
  assign _T_1886 = _GEN_69 | _T_1846; // @[Monitor.scala 708:24:freechips.rocketchip.system.DefaultRV32Config.fir@22247.6]
  assign _T_1887 = _T_1886 >> io_in_e_bits_sink; // @[Monitor.scala 708:35:freechips.rocketchip.system.DefaultRV32Config.fir@22248.6]
  assign _T_1890 = _T_1887[0] | reset; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@22251.6]
  assign _T_1891 = ~_T_1890; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@22252.6]
  assign _GEN_70 = io_in_e_valid ? _T_1885 : 4'h0; // @[Monitor.scala 706:73:freechips.rocketchip.system.DefaultRV32Config.fir@22244.4]
  assign _T_1892 = _T_1846 | _GEN_69; // @[Monitor.scala 713:27:freechips.rocketchip.system.DefaultRV32Config.fir@22258.4]
  assign _T_1893 = ~_GEN_70; // @[Monitor.scala 713:38:freechips.rocketchip.system.DefaultRV32Config.fir@22259.4]
  assign _T_1894 = _T_1892 & _T_1893; // @[Monitor.scala 713:36:freechips.rocketchip.system.DefaultRV32Config.fir@22260.4]
  assign _GEN_85 = io_in_a_valid & _T_78; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@19454.10]
  assign _GEN_101 = io_in_a_valid & _T_168; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@19583.10]
  assign _GEN_119 = io_in_a_valid & _T_262; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@19723.10]
  assign _GEN_131 = io_in_a_valid & _T_336; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@19830.10]
  assign _GEN_141 = io_in_a_valid & _T_413; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@19929.10]
  assign _GEN_151 = io_in_a_valid & _T_492; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@20020.10]
  assign _GEN_161 = io_in_a_valid & _T_559; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@20109.10]
  assign _GEN_171 = io_in_a_valid & _T_626; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@20198.10]
  assign _GEN_183 = io_in_d_valid & _T_708; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@20267.10]
  assign _GEN_193 = io_in_d_valid & _T_728; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@20309.10]
  assign _GEN_203 = io_in_d_valid & _T_756; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@20367.10]
  assign _GEN_213 = io_in_d_valid & _T_785; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@20426.10]
  assign _GEN_219 = io_in_d_valid & _T_802; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@20461.10]
  assign _GEN_225 = io_in_d_valid & _T_820; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@20497.10]
  assign _GEN_231 = io_in_c_valid & _T_1217; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@21152.10]
  assign _GEN_243 = io_in_c_valid & _T_1239; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@21200.10]
  assign _GEN_253 = io_in_c_valid & _T_1257; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@21289.10]
  assign _GEN_267 = io_in_c_valid & _T_1342; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@21409.10]
  assign _GEN_279 = io_in_c_valid & _T_1423; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@21472.10]
  assign _GEN_289 = io_in_c_valid & _T_1441; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@21512.10]
  assign _GEN_297 = io_in_c_valid & _T_1455; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@21544.10]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_1486 = _RAND_0[9:0];
  _RAND_1 = {1{`RANDOM}};
  _T_1497 = _RAND_1[2:0];
  _RAND_2 = {1{`RANDOM}};
  _T_1498 = _RAND_2[2:0];
  _RAND_3 = {1{`RANDOM}};
  _T_1499 = _RAND_3[3:0];
  _RAND_4 = {1{`RANDOM}};
  _T_1500 = _RAND_4[1:0];
  _RAND_5 = {1{`RANDOM}};
  _T_1501 = _RAND_5[31:0];
  _RAND_6 = {1{`RANDOM}};
  _T_1534 = _RAND_6[9:0];
  _RAND_7 = {1{`RANDOM}};
  _T_1545 = _RAND_7[2:0];
  _RAND_8 = {1{`RANDOM}};
  _T_1546 = _RAND_8[1:0];
  _RAND_9 = {1{`RANDOM}};
  _T_1547 = _RAND_9[3:0];
  _RAND_10 = {1{`RANDOM}};
  _T_1548 = _RAND_10[1:0];
  _RAND_11 = {1{`RANDOM}};
  _T_1549 = _RAND_11[1:0];
  _RAND_12 = {1{`RANDOM}};
  _T_1550 = _RAND_12[0:0];
  _RAND_13 = {1{`RANDOM}};
  _T_1588 = _RAND_13[9:0];
  _RAND_14 = {1{`RANDOM}};
  _T_1600 = _RAND_14[1:0];
  _RAND_15 = {1{`RANDOM}};
  _T_1603 = _RAND_15[31:0];
  _RAND_16 = {1{`RANDOM}};
  _T_1636 = _RAND_16[9:0];
  _RAND_17 = {1{`RANDOM}};
  _T_1647 = _RAND_17[2:0];
  _RAND_18 = {1{`RANDOM}};
  _T_1648 = _RAND_18[2:0];
  _RAND_19 = {1{`RANDOM}};
  _T_1649 = _RAND_19[3:0];
  _RAND_20 = {1{`RANDOM}};
  _T_1650 = _RAND_20[1:0];
  _RAND_21 = {1{`RANDOM}};
  _T_1651 = _RAND_21[31:0];
  _RAND_22 = {1{`RANDOM}};
  inflight = _RAND_22[2:0];
  _RAND_23 = {1{`RANDOM}};
  inflight_opcodes = _RAND_23[11:0];
  _RAND_24 = {1{`RANDOM}};
  inflight_sizes = _RAND_24[23:0];
  _RAND_25 = {1{`RANDOM}};
  _T_1685 = _RAND_25[9:0];
  _RAND_26 = {1{`RANDOM}};
  _T_1703 = _RAND_26[9:0];
  _RAND_27 = {1{`RANDOM}};
  _T_1831 = _RAND_27[31:0];
  _RAND_28 = {1{`RANDOM}};
  _T_1846 = _RAND_28[3:0];
  _RAND_29 = {1{`RANDOM}};
  _T_1855 = _RAND_29[9:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      _T_1486 <= 10'h0;
    end else if (_T_1477) begin
      if (_T_1489) begin
        if (_T_1484) begin
          _T_1486 <= _T_13[11:2];
        end else begin
          _T_1486 <= 10'h0;
        end
      end else begin
        _T_1486 <= _T_1488;
      end
    end
    if (_T_1525) begin
      _T_1497 <= io_in_a_bits_opcode;
    end
    if (_T_1525) begin
      _T_1498 <= io_in_a_bits_param;
    end
    if (_T_1525) begin
      _T_1499 <= io_in_a_bits_size;
    end
    if (_T_1525) begin
      _T_1500 <= io_in_a_bits_source;
    end
    if (_T_1525) begin
      _T_1501 <= io_in_a_bits_address;
    end
    if (reset) begin
      _T_1534 <= 10'h0;
    end else if (_T_1526) begin
      if (_T_1537) begin
        if (io_in_d_bits_opcode[0]) begin
          _T_1534 <= _T_1530[11:2];
        end else begin
          _T_1534 <= 10'h0;
        end
      end else begin
        _T_1534 <= _T_1536;
      end
    end
    if (_T_1578) begin
      _T_1545 <= io_in_d_bits_opcode;
    end
    if (_T_1578) begin
      _T_1546 <= io_in_d_bits_param;
    end
    if (_T_1578) begin
      _T_1547 <= io_in_d_bits_size;
    end
    if (_T_1578) begin
      _T_1548 <= io_in_d_bits_source;
    end
    if (_T_1578) begin
      _T_1549 <= io_in_d_bits_sink;
    end
    if (_T_1578) begin
      _T_1550 <= io_in_d_bits_denied;
    end
    if (reset) begin
      _T_1588 <= 10'h0;
    end else if (_T_1579) begin
      if (_T_1591) begin
        _T_1588 <= 10'h0;
      end else begin
        _T_1588 <= _T_1590;
      end
    end
    if (_T_1627) begin
      _T_1600 <= io_in_b_bits_param;
    end
    if (_T_1627) begin
      _T_1603 <= io_in_b_bits_address;
    end
    if (reset) begin
      _T_1636 <= 10'h0;
    end else if (_T_1628) begin
      if (_T_1639) begin
        if (io_in_c_bits_opcode[0]) begin
          _T_1636 <= _T_1143[11:2];
        end else begin
          _T_1636 <= 10'h0;
        end
      end else begin
        _T_1636 <= _T_1638;
      end
    end
    if (_T_1675) begin
      _T_1647 <= io_in_c_bits_opcode;
    end
    if (_T_1675) begin
      _T_1648 <= io_in_c_bits_param;
    end
    if (_T_1675) begin
      _T_1649 <= io_in_c_bits_size;
    end
    if (_T_1675) begin
      _T_1650 <= io_in_c_bits_source;
    end
    if (_T_1675) begin
      _T_1651 <= io_in_c_bits_address;
    end
    if (reset) begin
      inflight <= 3'h0;
    end else begin
      inflight <= _T_1824;
    end
    if (reset) begin
      inflight_opcodes <= 12'h0;
    end else begin
      inflight_opcodes <= _T_1827;
    end
    if (reset) begin
      inflight_sizes <= 24'h0;
    end else begin
      inflight_sizes <= _T_1830;
    end
    if (reset) begin
      _T_1685 <= 10'h0;
    end else if (_T_1477) begin
      if (a_first) begin
        if (_T_1484) begin
          _T_1685 <= _T_13[11:2];
        end else begin
          _T_1685 <= 10'h0;
        end
      end else begin
        _T_1685 <= _T_1687;
      end
    end
    if (reset) begin
      _T_1703 <= 10'h0;
    end else if (_T_1526) begin
      if (d_first) begin
        if (io_in_d_bits_opcode[0]) begin
          _T_1703 <= _T_1530[11:2];
        end else begin
          _T_1703 <= 10'h0;
        end
      end else begin
        _T_1703 <= _T_1705;
      end
    end
    if (reset) begin
      _T_1831 <= 32'h0;
    end else if (_T_1845) begin
      _T_1831 <= 32'h0;
    end else begin
      _T_1831 <= _T_1842;
    end
    if (reset) begin
      _T_1846 <= 4'h0;
    end else begin
      _T_1846 <= _T_1894;
    end
    if (reset) begin
      _T_1855 <= 10'h0;
    end else if (_T_1526) begin
      if (_T_1858) begin
        if (io_in_d_bits_opcode[0]) begin
          _T_1855 <= _T_1530[11:2];
        end else begin
          _T_1855 <= 10'h0;
        end
      end else begin
        _T_1855 <= _T_1857;
      end
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_85 & _T_130) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel carries AcquireBlock type unsupported by manager (connected at HasTiles.scala:49:43)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@19454.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_85 & _T_130) begin
          $fatal; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@19455.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_85 & _T_144) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel carries AcquireBlock from a client which does not support Probe (connected at HasTiles.scala:49:43)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@19477.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_85 & _T_144) begin
          $fatal; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@19478.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_85 & _T_147) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel AcquireBlock carries invalid source ID (connected at HasTiles.scala:49:43)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@19484.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_85 & _T_147) begin
          $fatal; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@19485.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_85 & _T_151) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel AcquireBlock smaller than a beat (connected at HasTiles.scala:49:43)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@19492.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_85 & _T_151) begin
          $fatal; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@19493.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_85 & _T_154) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel AcquireBlock address not aligned to size (connected at HasTiles.scala:49:43)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@19499.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_85 & _T_154) begin
          $fatal; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@19500.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_85 & _T_158) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel AcquireBlock carries invalid grow param (connected at HasTiles.scala:49:43)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@19507.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_85 & _T_158) begin
          $fatal; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@19508.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_85 & _T_163) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel AcquireBlock contains invalid mask (connected at HasTiles.scala:49:43)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@19516.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_85 & _T_163) begin
          $fatal; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@19517.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_85 & _T_167) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel AcquireBlock is corrupt (connected at HasTiles.scala:49:43)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@19524.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_85 & _T_167) begin
          $fatal; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@19525.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_101 & _T_130) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel carries AcquirePerm type unsupported by manager (connected at HasTiles.scala:49:43)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@19583.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_101 & _T_130) begin
          $fatal; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@19584.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_101 & _T_144) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel carries AcquirePerm from a client which does not support Probe (connected at HasTiles.scala:49:43)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@19606.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_101 & _T_144) begin
          $fatal; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@19607.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_101 & _T_147) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel AcquirePerm carries invalid source ID (connected at HasTiles.scala:49:43)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@19613.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_101 & _T_147) begin
          $fatal; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@19614.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_101 & _T_151) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel AcquirePerm smaller than a beat (connected at HasTiles.scala:49:43)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@19621.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_101 & _T_151) begin
          $fatal; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@19622.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_101 & _T_154) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel AcquirePerm address not aligned to size (connected at HasTiles.scala:49:43)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@19628.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_101 & _T_154) begin
          $fatal; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@19629.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_101 & _T_158) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel AcquirePerm carries invalid grow param (connected at HasTiles.scala:49:43)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@19636.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_101 & _T_158) begin
          $fatal; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@19637.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_101 & _T_252) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel AcquirePerm requests NtoB (connected at HasTiles.scala:49:43)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@19644.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_101 & _T_252) begin
          $fatal; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@19645.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_101 & _T_163) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel AcquirePerm contains invalid mask (connected at HasTiles.scala:49:43)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@19653.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_101 & _T_163) begin
          $fatal; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@19654.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_101 & _T_167) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel AcquirePerm is corrupt (connected at HasTiles.scala:49:43)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@19661.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_101 & _T_167) begin
          $fatal; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@19662.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_119 & _T_317) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel carries Get type unsupported by manager (connected at HasTiles.scala:49:43)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@19723.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_119 & _T_317) begin
          $fatal; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@19724.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_119 & _T_147) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel Get carries invalid source ID (connected at HasTiles.scala:49:43)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@19730.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_119 & _T_147) begin
          $fatal; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@19731.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_119 & _T_154) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel Get address not aligned to size (connected at HasTiles.scala:49:43)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@19737.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_119 & _T_154) begin
          $fatal; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@19738.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_119 & _T_327) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel Get carries invalid param (connected at HasTiles.scala:49:43)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@19745.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_119 & _T_327) begin
          $fatal; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@19746.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_119 & _T_331) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel Get contains invalid mask (connected at HasTiles.scala:49:43)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@19753.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_119 & _T_331) begin
          $fatal; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@19754.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_119 & _T_167) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel Get is corrupt (connected at HasTiles.scala:49:43)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@19761.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_119 & _T_167) begin
          $fatal; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@19762.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_131 & _T_398) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel carries PutFull type unsupported by manager (connected at HasTiles.scala:49:43)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@19830.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_131 & _T_398) begin
          $fatal; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@19831.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_131 & _T_147) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel PutFull carries invalid source ID (connected at HasTiles.scala:49:43)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@19837.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_131 & _T_147) begin
          $fatal; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@19838.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_131 & _T_154) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel PutFull address not aligned to size (connected at HasTiles.scala:49:43)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@19844.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_131 & _T_154) begin
          $fatal; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@19845.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_131 & _T_327) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel PutFull carries invalid param (connected at HasTiles.scala:49:43)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@19852.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_131 & _T_327) begin
          $fatal; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@19853.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_131 & _T_331) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel PutFull contains invalid mask (connected at HasTiles.scala:49:43)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@19860.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_131 & _T_331) begin
          $fatal; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@19861.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_141 & _T_398) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel carries PutPartial type unsupported by manager (connected at HasTiles.scala:49:43)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@19929.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_141 & _T_398) begin
          $fatal; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@19930.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_141 & _T_147) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel PutPartial carries invalid source ID (connected at HasTiles.scala:49:43)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@19936.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_141 & _T_147) begin
          $fatal; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@19937.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_141 & _T_154) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel PutPartial address not aligned to size (connected at HasTiles.scala:49:43)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@19943.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_141 & _T_154) begin
          $fatal; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@19944.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_141 & _T_327) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel PutPartial carries invalid param (connected at HasTiles.scala:49:43)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@19951.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_141 & _T_327) begin
          $fatal; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@19952.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_141 & _T_491) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel PutPartial contains invalid mask (connected at HasTiles.scala:49:43)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@19961.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_141 & _T_491) begin
          $fatal; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@19962.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_151 & _T_544) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel carries Arithmetic type unsupported by manager (connected at HasTiles.scala:49:43)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@20020.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_151 & _T_544) begin
          $fatal; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@20021.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_151 & _T_147) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel Arithmetic carries invalid source ID (connected at HasTiles.scala:49:43)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@20027.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_151 & _T_147) begin
          $fatal; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@20028.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_151 & _T_154) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel Arithmetic address not aligned to size (connected at HasTiles.scala:49:43)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@20034.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_151 & _T_154) begin
          $fatal; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@20035.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_151 & _T_554) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel Arithmetic carries invalid opcode param (connected at HasTiles.scala:49:43)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@20042.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_151 & _T_554) begin
          $fatal; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@20043.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_151 & _T_331) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel Arithmetic contains invalid mask (connected at HasTiles.scala:49:43)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@20050.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_151 & _T_331) begin
          $fatal; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@20051.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_161 & _T_544) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel carries Logical type unsupported by manager (connected at HasTiles.scala:49:43)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@20109.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_161 & _T_544) begin
          $fatal; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@20110.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_161 & _T_147) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel Logical carries invalid source ID (connected at HasTiles.scala:49:43)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@20116.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_161 & _T_147) begin
          $fatal; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@20117.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_161 & _T_154) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel Logical address not aligned to size (connected at HasTiles.scala:49:43)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@20123.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_161 & _T_154) begin
          $fatal; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@20124.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_161 & _T_621) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel Logical carries invalid opcode param (connected at HasTiles.scala:49:43)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@20131.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_161 & _T_621) begin
          $fatal; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@20132.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_161 & _T_331) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel Logical contains invalid mask (connected at HasTiles.scala:49:43)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@20139.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_161 & _T_331) begin
          $fatal; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@20140.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_171 & _T_678) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel carries Hint type unsupported by manager (connected at HasTiles.scala:49:43)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@20198.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_171 & _T_678) begin
          $fatal; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@20199.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_171 & _T_147) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel Hint carries invalid source ID (connected at HasTiles.scala:49:43)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@20205.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_171 & _T_147) begin
          $fatal; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@20206.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_171 & _T_154) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel Hint address not aligned to size (connected at HasTiles.scala:49:43)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@20212.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_171 & _T_154) begin
          $fatal; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@20213.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_171 & _T_688) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel Hint carries invalid opcode param (connected at HasTiles.scala:49:43)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@20220.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_171 & _T_688) begin
          $fatal; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@20221.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_171 & _T_331) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel Hint contains invalid mask (connected at HasTiles.scala:49:43)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@20228.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_171 & _T_331) begin
          $fatal; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@20229.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_171 & _T_167) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel Hint is corrupt (connected at HasTiles.scala:49:43)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@20236.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_171 & _T_167) begin
          $fatal; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@20237.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_d_valid & _T_700) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel has invalid opcode (connected at HasTiles.scala:49:43)\n    at Monitor.scala:51 assert(cond, message)\n"); // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@20247.8]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_d_valid & _T_700) begin
          $fatal; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@20248.8]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_183 & _T_711) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel ReleaseAck carries invalid source ID (connected at HasTiles.scala:49:43)\n    at Monitor.scala:51 assert(cond, message)\n"); // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@20267.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_183 & _T_711) begin
          $fatal; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@20268.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_183 & _T_715) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel ReleaseAck smaller than a beat (connected at HasTiles.scala:49:43)\n    at Monitor.scala:51 assert(cond, message)\n"); // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@20275.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_183 & _T_715) begin
          $fatal; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@20276.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_183 & _T_719) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel ReleaseeAck carries invalid param (connected at HasTiles.scala:49:43)\n    at Monitor.scala:51 assert(cond, message)\n"); // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@20283.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_183 & _T_719) begin
          $fatal; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@20284.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_183 & _T_723) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel ReleaseAck is corrupt (connected at HasTiles.scala:49:43)\n    at Monitor.scala:51 assert(cond, message)\n"); // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@20291.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_183 & _T_723) begin
          $fatal; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@20292.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_183 & _T_727) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel ReleaseAck is denied (connected at HasTiles.scala:49:43)\n    at Monitor.scala:51 assert(cond, message)\n"); // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@20299.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_183 & _T_727) begin
          $fatal; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@20300.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_193 & _T_711) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel Grant carries invalid source ID (connected at HasTiles.scala:49:43)\n    at Monitor.scala:51 assert(cond, message)\n"); // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@20309.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_193 & _T_711) begin
          $fatal; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@20310.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_193 & _T_715) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel Grant smaller than a beat (connected at HasTiles.scala:49:43)\n    at Monitor.scala:51 assert(cond, message)\n"); // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@20324.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_193 & _T_715) begin
          $fatal; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@20325.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_193 & _T_742) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel Grant carries invalid cap param (connected at HasTiles.scala:49:43)\n    at Monitor.scala:51 assert(cond, message)\n"); // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@20332.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_193 & _T_742) begin
          $fatal; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@20333.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_193 & _T_746) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel Grant carries toN param (connected at HasTiles.scala:49:43)\n    at Monitor.scala:51 assert(cond, message)\n"); // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@20340.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_193 & _T_746) begin
          $fatal; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@20341.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_193 & _T_723) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel Grant is corrupt (connected at HasTiles.scala:49:43)\n    at Monitor.scala:51 assert(cond, message)\n"); // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@20348.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_193 & _T_723) begin
          $fatal; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@20349.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_203 & _T_711) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel GrantData carries invalid source ID (connected at HasTiles.scala:49:43)\n    at Monitor.scala:51 assert(cond, message)\n"); // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@20367.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_203 & _T_711) begin
          $fatal; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@20368.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_203 & _T_715) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel GrantData smaller than a beat (connected at HasTiles.scala:49:43)\n    at Monitor.scala:51 assert(cond, message)\n"); // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@20382.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_203 & _T_715) begin
          $fatal; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@20383.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_203 & _T_742) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel GrantData carries invalid cap param (connected at HasTiles.scala:49:43)\n    at Monitor.scala:51 assert(cond, message)\n"); // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@20390.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_203 & _T_742) begin
          $fatal; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@20391.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_203 & _T_746) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel GrantData carries toN param (connected at HasTiles.scala:49:43)\n    at Monitor.scala:51 assert(cond, message)\n"); // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@20398.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_203 & _T_746) begin
          $fatal; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@20399.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_203 & _T_779) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel GrantData is denied but not corrupt (connected at HasTiles.scala:49:43)\n    at Monitor.scala:51 assert(cond, message)\n"); // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@20407.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_203 & _T_779) begin
          $fatal; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@20408.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_213 & _T_711) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel AccessAck carries invalid source ID (connected at HasTiles.scala:49:43)\n    at Monitor.scala:51 assert(cond, message)\n"); // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@20426.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_213 & _T_711) begin
          $fatal; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@20427.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_213 & _T_719) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel AccessAck carries invalid param (connected at HasTiles.scala:49:43)\n    at Monitor.scala:51 assert(cond, message)\n"); // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@20434.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_213 & _T_719) begin
          $fatal; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@20435.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_213 & _T_723) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel AccessAck is corrupt (connected at HasTiles.scala:49:43)\n    at Monitor.scala:51 assert(cond, message)\n"); // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@20442.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_213 & _T_723) begin
          $fatal; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@20443.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_219 & _T_711) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel AccessAckData carries invalid source ID (connected at HasTiles.scala:49:43)\n    at Monitor.scala:51 assert(cond, message)\n"); // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@20461.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_219 & _T_711) begin
          $fatal; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@20462.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_219 & _T_719) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel AccessAckData carries invalid param (connected at HasTiles.scala:49:43)\n    at Monitor.scala:51 assert(cond, message)\n"); // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@20469.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_219 & _T_719) begin
          $fatal; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@20470.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_219 & _T_779) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel AccessAckData is denied but not corrupt (connected at HasTiles.scala:49:43)\n    at Monitor.scala:51 assert(cond, message)\n"); // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@20478.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_219 & _T_779) begin
          $fatal; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@20479.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_225 & _T_711) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel HintAck carries invalid source ID (connected at HasTiles.scala:49:43)\n    at Monitor.scala:51 assert(cond, message)\n"); // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@20497.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_225 & _T_711) begin
          $fatal; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@20498.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_225 & _T_719) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel HintAck carries invalid param (connected at HasTiles.scala:49:43)\n    at Monitor.scala:51 assert(cond, message)\n"); // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@20505.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_225 & _T_719) begin
          $fatal; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@20506.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_225 & _T_723) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel HintAck is corrupt (connected at HasTiles.scala:49:43)\n    at Monitor.scala:51 assert(cond, message)\n"); // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@20513.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_225 & _T_723) begin
          $fatal; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@20514.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_b_valid & _T_979) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel Probe carries unmanaged address (connected at HasTiles.scala:49:43)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@20703.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_b_valid & _T_979) begin
          $fatal; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@20704.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_b_valid & _T_985) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel Probe address not aligned to size (connected at HasTiles.scala:49:43)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@20717.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_b_valid & _T_985) begin
          $fatal; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@20718.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_b_valid & _T_989) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel Probe carries invalid cap param (connected at HasTiles.scala:49:43)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@20725.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_b_valid & _T_989) begin
          $fatal; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@20726.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_231 & _T_1220) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel ProbeAck carries unmanaged address (connected at HasTiles.scala:49:43)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@21152.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_231 & _T_1220) begin
          $fatal; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@21153.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_231 & _T_1223) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel ProbeAck carries invalid source ID (connected at HasTiles.scala:49:43)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@21159.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_231 & _T_1223) begin
          $fatal; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@21160.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_231 & _T_1227) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel ProbeAck smaller than a beat (connected at HasTiles.scala:49:43)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@21167.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_231 & _T_1227) begin
          $fatal; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@21168.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_231 & _T_1230) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel ProbeAck address not aligned to size (connected at HasTiles.scala:49:43)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@21174.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_231 & _T_1230) begin
          $fatal; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@21175.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_231 & _T_1234) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel ProbeAck carries invalid report param (connected at HasTiles.scala:49:43)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@21182.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_231 & _T_1234) begin
          $fatal; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@21183.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_231 & _T_1238) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel ProbeAck is corrupt (connected at HasTiles.scala:49:43)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@21190.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_231 & _T_1238) begin
          $fatal; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@21191.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_243 & _T_1220) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel ProbeAckData carries unmanaged address (connected at HasTiles.scala:49:43)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@21200.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_243 & _T_1220) begin
          $fatal; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@21201.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_243 & _T_1223) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel ProbeAckData carries invalid source ID (connected at HasTiles.scala:49:43)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@21207.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_243 & _T_1223) begin
          $fatal; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@21208.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_243 & _T_1227) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel ProbeAckData smaller than a beat (connected at HasTiles.scala:49:43)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@21215.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_243 & _T_1227) begin
          $fatal; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@21216.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_243 & _T_1230) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel ProbeAckData address not aligned to size (connected at HasTiles.scala:49:43)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@21222.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_243 & _T_1230) begin
          $fatal; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@21223.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_243 & _T_1234) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel ProbeAckData carries invalid report param (connected at HasTiles.scala:49:43)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@21230.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_243 & _T_1234) begin
          $fatal; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@21231.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_253 & _T_1309) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel carries Release type unsupported by manager (connected at HasTiles.scala:49:43)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@21289.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_253 & _T_1309) begin
          $fatal; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@21290.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_253 & _T_1323) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel carries Release from a client which does not support Probe (connected at HasTiles.scala:49:43)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@21312.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_253 & _T_1323) begin
          $fatal; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@21313.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_253 & _T_1223) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel Release carries invalid source ID (connected at HasTiles.scala:49:43)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@21319.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_253 & _T_1223) begin
          $fatal; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@21320.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_253 & _T_1227) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel Release smaller than a beat (connected at HasTiles.scala:49:43)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@21327.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_253 & _T_1227) begin
          $fatal; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@21328.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_253 & _T_1230) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel Release address not aligned to size (connected at HasTiles.scala:49:43)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@21334.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_253 & _T_1230) begin
          $fatal; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@21335.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_253 & _T_1337) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel Release carries invalid shrink param (connected at HasTiles.scala:49:43)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@21342.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_253 & _T_1337) begin
          $fatal; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@21343.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_253 & _T_1238) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel Release is corrupt (connected at HasTiles.scala:49:43)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@21350.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_253 & _T_1238) begin
          $fatal; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@21351.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_267 & _T_1309) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel carries ReleaseData type unsupported by manager (connected at HasTiles.scala:49:43)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@21409.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_267 & _T_1309) begin
          $fatal; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@21410.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_267 & _T_1323) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel carries Release from a client which does not support Probe (connected at HasTiles.scala:49:43)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@21432.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_267 & _T_1323) begin
          $fatal; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@21433.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_267 & _T_1223) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel ReleaseData carries invalid source ID (connected at HasTiles.scala:49:43)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@21439.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_267 & _T_1223) begin
          $fatal; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@21440.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_267 & _T_1227) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel ReleaseData smaller than a beat (connected at HasTiles.scala:49:43)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@21447.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_267 & _T_1227) begin
          $fatal; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@21448.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_267 & _T_1230) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel ReleaseData address not aligned to size (connected at HasTiles.scala:49:43)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@21454.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_267 & _T_1230) begin
          $fatal; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@21455.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_267 & _T_1337) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel ReleaseData carries invalid shrink param (connected at HasTiles.scala:49:43)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@21462.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_267 & _T_1337) begin
          $fatal; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@21463.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_279 & _T_1220) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel AccessAck carries unmanaged address (connected at HasTiles.scala:49:43)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@21472.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_279 & _T_1220) begin
          $fatal; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@21473.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_279 & _T_1223) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel AccessAck carries invalid source ID (connected at HasTiles.scala:49:43)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@21479.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_279 & _T_1223) begin
          $fatal; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@21480.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_279 & _T_1230) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel AccessAck address not aligned to size (connected at HasTiles.scala:49:43)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@21486.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_279 & _T_1230) begin
          $fatal; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@21487.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_279 & _T_1436) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel AccessAck carries invalid param (connected at HasTiles.scala:49:43)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@21494.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_279 & _T_1436) begin
          $fatal; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@21495.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_279 & _T_1238) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel AccessAck is corrupt (connected at HasTiles.scala:49:43)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@21502.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_279 & _T_1238) begin
          $fatal; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@21503.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_289 & _T_1220) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel AccessAckData carries unmanaged address (connected at HasTiles.scala:49:43)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@21512.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_289 & _T_1220) begin
          $fatal; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@21513.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_289 & _T_1223) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel AccessAckData carries invalid source ID (connected at HasTiles.scala:49:43)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@21519.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_289 & _T_1223) begin
          $fatal; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@21520.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_289 & _T_1230) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel AccessAckData address not aligned to size (connected at HasTiles.scala:49:43)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@21526.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_289 & _T_1230) begin
          $fatal; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@21527.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_289 & _T_1436) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel AccessAckData carries invalid param (connected at HasTiles.scala:49:43)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@21534.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_289 & _T_1436) begin
          $fatal; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@21535.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_297 & _T_1220) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel HintAck carries unmanaged address (connected at HasTiles.scala:49:43)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@21544.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_297 & _T_1220) begin
          $fatal; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@21545.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_297 & _T_1223) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel HintAck carries invalid source ID (connected at HasTiles.scala:49:43)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@21551.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_297 & _T_1223) begin
          $fatal; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@21552.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_297 & _T_1230) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel HintAck address not aligned to size (connected at HasTiles.scala:49:43)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@21558.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_297 & _T_1230) begin
          $fatal; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@21559.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_297 & _T_1436) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel HintAck carries invalid param (connected at HasTiles.scala:49:43)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@21566.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_297 & _T_1436) begin
          $fatal; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@21567.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_297 & _T_1238) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel HintAck is corrupt (connected at HasTiles.scala:49:43)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@21574.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_297 & _T_1238) begin
          $fatal; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@21575.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1503 & _T_1507) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel opcode changed within multibeat operation (connected at HasTiles.scala:49:43)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@21625.8]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_1503 & _T_1507) begin
          $fatal; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@21626.8]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1503 & _T_1511) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel param changed within multibeat operation (connected at HasTiles.scala:49:43)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@21633.8]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_1503 & _T_1511) begin
          $fatal; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@21634.8]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1503 & _T_1515) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel size changed within multibeat operation (connected at HasTiles.scala:49:43)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@21641.8]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_1503 & _T_1515) begin
          $fatal; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@21642.8]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1503 & _T_1519) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel source changed within multibeat operation (connected at HasTiles.scala:49:43)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@21649.8]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_1503 & _T_1519) begin
          $fatal; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@21650.8]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1503 & _T_1523) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel address changed with multibeat operation (connected at HasTiles.scala:49:43)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@21657.8]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_1503 & _T_1523) begin
          $fatal; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@21658.8]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1552 & _T_1556) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel opcode changed within multibeat operation (connected at HasTiles.scala:49:43)\n    at Monitor.scala:51 assert(cond, message)\n"); // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@21706.8]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_1552 & _T_1556) begin
          $fatal; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@21707.8]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1552 & _T_1560) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel param changed within multibeat operation (connected at HasTiles.scala:49:43)\n    at Monitor.scala:51 assert(cond, message)\n"); // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@21714.8]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_1552 & _T_1560) begin
          $fatal; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@21715.8]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1552 & _T_1564) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel size changed within multibeat operation (connected at HasTiles.scala:49:43)\n    at Monitor.scala:51 assert(cond, message)\n"); // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@21722.8]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_1552 & _T_1564) begin
          $fatal; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@21723.8]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1552 & _T_1568) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel source changed within multibeat operation (connected at HasTiles.scala:49:43)\n    at Monitor.scala:51 assert(cond, message)\n"); // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@21730.8]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_1552 & _T_1568) begin
          $fatal; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@21731.8]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1552 & _T_1572) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel sink changed with multibeat operation (connected at HasTiles.scala:49:43)\n    at Monitor.scala:51 assert(cond, message)\n"); // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@21738.8]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_1552 & _T_1572) begin
          $fatal; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@21739.8]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1552 & _T_1576) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel denied changed with multibeat operation (connected at HasTiles.scala:49:43)\n    at Monitor.scala:51 assert(cond, message)\n"); // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@21746.8]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_1552 & _T_1576) begin
          $fatal; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@21747.8]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1605 & _T_1613) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel param changed within multibeat operation (connected at HasTiles.scala:49:43)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@21804.8]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_1605 & _T_1613) begin
          $fatal; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@21805.8]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1605 & _T_1625) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel addresss changed with multibeat operation (connected at HasTiles.scala:49:43)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@21828.8]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_1605 & _T_1625) begin
          $fatal; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@21829.8]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1653 & _T_1657) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel opcode changed within multibeat operation (connected at HasTiles.scala:49:43)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@21876.8]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_1653 & _T_1657) begin
          $fatal; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@21877.8]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1653 & _T_1661) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel param changed within multibeat operation (connected at HasTiles.scala:49:43)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@21884.8]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_1653 & _T_1661) begin
          $fatal; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@21885.8]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1653 & _T_1665) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel size changed within multibeat operation (connected at HasTiles.scala:49:43)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@21892.8]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_1653 & _T_1665) begin
          $fatal; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@21893.8]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1653 & _T_1669) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel source changed within multibeat operation (connected at HasTiles.scala:49:43)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@21900.8]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_1653 & _T_1669) begin
          $fatal; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@21901.8]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1653 & _T_1673) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel address changed with multibeat operation (connected at HasTiles.scala:49:43)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@21908.8]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_1653 & _T_1673) begin
          $fatal; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@21909.8]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1732 & _T_1748) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel re-used a source ID (connected at HasTiles.scala:49:43)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@22044.8]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_1732 & _T_1748) begin
          $fatal; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@22045.8]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1771 & _T_1782) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel acknowledged for nothing inflight (connected at HasTiles.scala:49:43)\n    at Monitor.scala:51 assert(cond, message)\n"); // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@22095.8]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_1771 & _T_1782) begin
          $fatal; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@22096.8]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1771 & _T_1795) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel contains improper opcode response (connected at HasTiles.scala:49:43)\n    at Monitor.scala:51 assert(cond, message)\n"); // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@22112.8]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_1771 & _T_1795) begin
          $fatal; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@22113.8]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1771 & _T_1802) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel contains improper response size (connected at HasTiles.scala:49:43)\n    at Monitor.scala:51 assert(cond, message)\n"); // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@22123.8]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_1771 & _T_1802) begin
          $fatal; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@22124.8]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1809 & _T_1814) begin
          $fwrite(32'h80000002,"Assertion failed: ready check\n    at Monitor.scala:51 assert(cond, message)\n"); // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@22141.8]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_1809 & _T_1814) begin
          $fatal; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@22142.8]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1821) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' and 'D' concurrent, despite minlatency 1 (connected at HasTiles.scala:49:43)\n    at Monitor.scala:51 assert(cond, message)\n"); // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@22153.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_1821) begin
          $fatal; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@22154.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1840) begin
          $fwrite(32'h80000002,"Assertion failed: TileLink timeout expired (connected at HasTiles.scala:49:43)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@22181.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_1840) begin
          $fatal; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@22182.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1873 & _T_1880) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel re-used a sink ID (connected at HasTiles.scala:49:43)\n    at Monitor.scala:51 assert(cond, message)\n"); // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@22235.8]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_1873 & _T_1880) begin
          $fatal; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@22236.8]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_e_valid & _T_1891) begin
          $fwrite(32'h80000002,"Assertion failed: 'E' channel acknowledged for nothing inflight (connected at HasTiles.scala:49:43)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@22254.8]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_e_valid & _T_1891) begin
          $fatal; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@22255.8]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
  end
endmodule
