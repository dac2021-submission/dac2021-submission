module OptimizationBarrier_117( // @[:freechips.rocketchip.system.DefaultRV32Config.fir@214049.2]
  input  [2:0] io_x, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@214052.4]
  output [2:0] io_y // @[:freechips.rocketchip.system.DefaultRV32Config.fir@214052.4]
);
  assign io_y = io_x; // @[package.scala 236:12:freechips.rocketchip.system.DefaultRV32Config.fir@214057.4]
endmodule
