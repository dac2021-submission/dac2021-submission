module DCache( // @[:freechips.rocketchip.system.DefaultRV32Config.fir@192092.2]
  input         gated_clock, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@192093.4]
  input         reset, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@192094.4]
  input         auto_out_a_ready, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@192095.4]
  output        auto_out_a_valid, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@192095.4]
  output [2:0]  auto_out_a_bits_opcode, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@192095.4]
  output [2:0]  auto_out_a_bits_param, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@192095.4]
  output [3:0]  auto_out_a_bits_size, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@192095.4]
  output        auto_out_a_bits_source, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@192095.4]
  output [31:0] auto_out_a_bits_address, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@192095.4]
  output [3:0]  auto_out_a_bits_mask, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@192095.4]
  output [31:0] auto_out_a_bits_data, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@192095.4]
  output        auto_out_b_ready, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@192095.4]
  input         auto_out_b_valid, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@192095.4]
  input  [1:0]  auto_out_b_bits_param, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@192095.4]
  input  [3:0]  auto_out_b_bits_size, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@192095.4]
  input         auto_out_b_bits_source, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@192095.4]
  input  [31:0] auto_out_b_bits_address, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@192095.4]
  input         auto_out_c_ready, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@192095.4]
  output        auto_out_c_valid, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@192095.4]
  output [2:0]  auto_out_c_bits_opcode, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@192095.4]
  output [2:0]  auto_out_c_bits_param, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@192095.4]
  output [3:0]  auto_out_c_bits_size, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@192095.4]
  output        auto_out_c_bits_source, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@192095.4]
  output [31:0] auto_out_c_bits_address, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@192095.4]
  output [31:0] auto_out_c_bits_data, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@192095.4]
  output        auto_out_d_ready, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@192095.4]
  input         auto_out_d_valid, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@192095.4]
  input  [2:0]  auto_out_d_bits_opcode, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@192095.4]
  input  [1:0]  auto_out_d_bits_param, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@192095.4]
  input  [3:0]  auto_out_d_bits_size, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@192095.4]
  input         auto_out_d_bits_source, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@192095.4]
  input  [1:0]  auto_out_d_bits_sink, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@192095.4]
  input         auto_out_d_bits_denied, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@192095.4]
  input  [31:0] auto_out_d_bits_data, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@192095.4]
  input         auto_out_e_ready, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@192095.4]
  output        auto_out_e_valid, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@192095.4]
  output [1:0]  auto_out_e_bits_sink, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@192095.4]
  output        io_cpu_req_ready, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@192096.4]
  input         io_cpu_req_valid, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@192096.4]
  input  [31:0] io_cpu_req_bits_addr, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@192096.4]
  input  [6:0]  io_cpu_req_bits_tag, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@192096.4]
  input  [4:0]  io_cpu_req_bits_cmd, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@192096.4]
  input  [1:0]  io_cpu_req_bits_size, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@192096.4]
  input         io_cpu_req_bits_signed, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@192096.4]
  input  [1:0]  io_cpu_req_bits_dprv, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@192096.4]
  input         io_cpu_req_bits_phys, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@192096.4]
  input         io_cpu_s1_kill, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@192096.4]
  input  [31:0] io_cpu_s1_data_data, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@192096.4]
  input  [3:0]  io_cpu_s1_data_mask, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@192096.4]
  output        io_cpu_s2_nack, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@192096.4]
  output        io_cpu_resp_valid, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@192096.4]
  output [31:0] io_cpu_resp_bits_addr, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@192096.4]
  output [6:0]  io_cpu_resp_bits_tag, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@192096.4]
  output [4:0]  io_cpu_resp_bits_cmd, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@192096.4]
  output [1:0]  io_cpu_resp_bits_size, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@192096.4]
  output        io_cpu_resp_bits_signed, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@192096.4]
  output [1:0]  io_cpu_resp_bits_dprv, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@192096.4]
  output [31:0] io_cpu_resp_bits_data, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@192096.4]
  output [3:0]  io_cpu_resp_bits_mask, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@192096.4]
  output        io_cpu_resp_bits_replay, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@192096.4]
  output        io_cpu_resp_bits_has_data, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@192096.4]
  output [31:0] io_cpu_resp_bits_data_word_bypass, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@192096.4]
  output [31:0] io_cpu_resp_bits_data_raw, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@192096.4]
  output [31:0] io_cpu_resp_bits_store_data, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@192096.4]
  output        io_cpu_replay_next, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@192096.4]
  output        io_cpu_s2_xcpt_ma_ld, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@192096.4]
  output        io_cpu_s2_xcpt_ma_st, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@192096.4]
  output        io_cpu_s2_xcpt_pf_ld, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@192096.4]
  output        io_cpu_s2_xcpt_pf_st, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@192096.4]
  output        io_cpu_s2_xcpt_ae_ld, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@192096.4]
  output        io_cpu_s2_xcpt_ae_st, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@192096.4]
  output        io_cpu_ordered, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@192096.4]
  output        io_cpu_perf_release, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@192096.4]
  output        io_cpu_perf_grant, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@192096.4]
  input         io_ptw_req_ready, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@192096.4]
  output        io_ptw_req_valid, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@192096.4]
  output [19:0] io_ptw_req_bits_bits_addr, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@192096.4]
  input         io_ptw_resp_valid, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@192096.4]
  input         io_ptw_resp_bits_ae, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@192096.4]
  input  [53:0] io_ptw_resp_bits_pte_ppn, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@192096.4]
  input         io_ptw_resp_bits_pte_d, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@192096.4]
  input         io_ptw_resp_bits_pte_a, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@192096.4]
  input         io_ptw_resp_bits_pte_g, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@192096.4]
  input         io_ptw_resp_bits_pte_u, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@192096.4]
  input         io_ptw_resp_bits_pte_x, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@192096.4]
  input         io_ptw_resp_bits_pte_w, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@192096.4]
  input         io_ptw_resp_bits_pte_r, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@192096.4]
  input         io_ptw_resp_bits_pte_v, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@192096.4]
  input         io_ptw_resp_bits_level, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@192096.4]
  input         io_ptw_resp_bits_homogeneous, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@192096.4]
  input         io_ptw_ptbr_mode, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@192096.4]
  input         io_ptw_status_debug, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@192096.4]
  input  [1:0]  io_ptw_status_dprv, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@192096.4]
  input         io_ptw_status_mxr, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@192096.4]
  input         io_ptw_status_sum, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@192096.4]
  input         io_ptw_pmp_0_cfg_l, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@192096.4]
  input  [1:0]  io_ptw_pmp_0_cfg_a, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@192096.4]
  input         io_ptw_pmp_0_cfg_x, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@192096.4]
  input         io_ptw_pmp_0_cfg_w, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@192096.4]
  input         io_ptw_pmp_0_cfg_r, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@192096.4]
  input  [29:0] io_ptw_pmp_0_addr, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@192096.4]
  input  [31:0] io_ptw_pmp_0_mask, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@192096.4]
  input         io_ptw_pmp_1_cfg_l, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@192096.4]
  input  [1:0]  io_ptw_pmp_1_cfg_a, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@192096.4]
  input         io_ptw_pmp_1_cfg_x, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@192096.4]
  input         io_ptw_pmp_1_cfg_w, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@192096.4]
  input         io_ptw_pmp_1_cfg_r, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@192096.4]
  input  [29:0] io_ptw_pmp_1_addr, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@192096.4]
  input  [31:0] io_ptw_pmp_1_mask, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@192096.4]
  input         io_ptw_pmp_2_cfg_l, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@192096.4]
  input  [1:0]  io_ptw_pmp_2_cfg_a, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@192096.4]
  input         io_ptw_pmp_2_cfg_x, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@192096.4]
  input         io_ptw_pmp_2_cfg_w, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@192096.4]
  input         io_ptw_pmp_2_cfg_r, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@192096.4]
  input  [29:0] io_ptw_pmp_2_addr, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@192096.4]
  input  [31:0] io_ptw_pmp_2_mask, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@192096.4]
  input         io_ptw_pmp_3_cfg_l, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@192096.4]
  input  [1:0]  io_ptw_pmp_3_cfg_a, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@192096.4]
  input         io_ptw_pmp_3_cfg_x, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@192096.4]
  input         io_ptw_pmp_3_cfg_w, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@192096.4]
  input         io_ptw_pmp_3_cfg_r, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@192096.4]
  input  [29:0] io_ptw_pmp_3_addr, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@192096.4]
  input  [31:0] io_ptw_pmp_3_mask, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@192096.4]
  input         io_ptw_pmp_4_cfg_l, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@192096.4]
  input  [1:0]  io_ptw_pmp_4_cfg_a, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@192096.4]
  input         io_ptw_pmp_4_cfg_x, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@192096.4]
  input         io_ptw_pmp_4_cfg_w, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@192096.4]
  input         io_ptw_pmp_4_cfg_r, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@192096.4]
  input  [29:0] io_ptw_pmp_4_addr, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@192096.4]
  input  [31:0] io_ptw_pmp_4_mask, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@192096.4]
  input         io_ptw_pmp_5_cfg_l, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@192096.4]
  input  [1:0]  io_ptw_pmp_5_cfg_a, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@192096.4]
  input         io_ptw_pmp_5_cfg_x, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@192096.4]
  input         io_ptw_pmp_5_cfg_w, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@192096.4]
  input         io_ptw_pmp_5_cfg_r, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@192096.4]
  input  [29:0] io_ptw_pmp_5_addr, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@192096.4]
  input  [31:0] io_ptw_pmp_5_mask, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@192096.4]
  input         io_ptw_pmp_6_cfg_l, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@192096.4]
  input  [1:0]  io_ptw_pmp_6_cfg_a, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@192096.4]
  input         io_ptw_pmp_6_cfg_x, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@192096.4]
  input         io_ptw_pmp_6_cfg_w, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@192096.4]
  input         io_ptw_pmp_6_cfg_r, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@192096.4]
  input  [29:0] io_ptw_pmp_6_addr, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@192096.4]
  input  [31:0] io_ptw_pmp_6_mask, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@192096.4]
  input         io_ptw_pmp_7_cfg_l, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@192096.4]
  input  [1:0]  io_ptw_pmp_7_cfg_a, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@192096.4]
  input         io_ptw_pmp_7_cfg_x, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@192096.4]
  input         io_ptw_pmp_7_cfg_w, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@192096.4]
  input         io_ptw_pmp_7_cfg_r, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@192096.4]
  input  [29:0] io_ptw_pmp_7_addr, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@192096.4]
  input  [31:0] io_ptw_pmp_7_mask // @[:freechips.rocketchip.system.DefaultRV32Config.fir@192096.4]
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [63:0] _RAND_1;
  reg [63:0] _RAND_2;
  reg [63:0] _RAND_3;
  reg [63:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [63:0] _RAND_10;
  reg [63:0] _RAND_11;
  reg [63:0] _RAND_12;
  reg [63:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [63:0] _RAND_19;
  reg [63:0] _RAND_20;
  reg [63:0] _RAND_21;
  reg [63:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [63:0] _RAND_28;
  reg [63:0] _RAND_29;
  reg [63:0] _RAND_30;
  reg [63:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [31:0] _RAND_34;
  reg [31:0] _RAND_35;
  reg [31:0] _RAND_36;
  reg [63:0] _RAND_37;
  reg [63:0] _RAND_38;
  reg [63:0] _RAND_39;
  reg [63:0] _RAND_40;
  reg [31:0] _RAND_41;
  reg [31:0] _RAND_42;
  reg [31:0] _RAND_43;
  reg [31:0] _RAND_44;
  reg [31:0] _RAND_45;
  reg [63:0] _RAND_46;
  reg [63:0] _RAND_47;
  reg [63:0] _RAND_48;
  reg [63:0] _RAND_49;
  reg [31:0] _RAND_50;
  reg [31:0] _RAND_51;
  reg [31:0] _RAND_52;
  reg [31:0] _RAND_53;
  reg [31:0] _RAND_54;
  reg [63:0] _RAND_55;
  reg [63:0] _RAND_56;
  reg [63:0] _RAND_57;
  reg [63:0] _RAND_58;
  reg [31:0] _RAND_59;
  reg [31:0] _RAND_60;
  reg [31:0] _RAND_61;
  reg [31:0] _RAND_62;
  reg [31:0] _RAND_63;
  reg [63:0] _RAND_64;
  reg [63:0] _RAND_65;
  reg [63:0] _RAND_66;
  reg [63:0] _RAND_67;
  reg [31:0] _RAND_68;
  reg [31:0] _RAND_69;
  reg [31:0] _RAND_70;
  reg [31:0] _RAND_71;
  reg [31:0] _RAND_72;
  reg [63:0] _RAND_73;
  reg [31:0] _RAND_74;
  reg [31:0] _RAND_75;
  reg [63:0] _RAND_76;
  reg [31:0] _RAND_77;
  reg [31:0] _RAND_78;
  reg [63:0] _RAND_79;
  reg [31:0] _RAND_80;
  reg [31:0] _RAND_81;
  reg [63:0] _RAND_82;
  reg [31:0] _RAND_83;
  reg [31:0] _RAND_84;
  reg [31:0] _RAND_85;
  reg [63:0] _RAND_86;
  reg [31:0] _RAND_87;
  reg [31:0] _RAND_88;
  reg [31:0] _RAND_89;
  reg [31:0] _RAND_90;
  reg [31:0] _RAND_91;
  reg [31:0] _RAND_92;
  reg [31:0] _RAND_93;
  reg [31:0] _RAND_94;
  reg [31:0] _RAND_95;
  reg [31:0] _RAND_96;
  reg [31:0] _RAND_97;
  reg [31:0] _RAND_98;
  reg [31:0] _RAND_99;
  reg [31:0] _RAND_100;
  reg [31:0] _RAND_101;
  reg [31:0] _RAND_102;
  reg [31:0] _RAND_103;
  reg [31:0] _RAND_104;
  reg [31:0] _RAND_105;
  reg [31:0] _RAND_106;
  reg [31:0] _RAND_107;
  reg [31:0] _RAND_108;
  reg [31:0] _RAND_109;
  reg [31:0] _RAND_110;
  reg [31:0] _RAND_111;
  reg [31:0] _RAND_112;
  reg [31:0] _RAND_113;
  reg [31:0] _RAND_114;
  reg [31:0] _RAND_115;
  reg [31:0] _RAND_116;
  reg [31:0] _RAND_117;
  reg [31:0] _RAND_118;
  reg [31:0] _RAND_119;
  reg [31:0] _RAND_120;
  reg [31:0] _RAND_121;
  reg [31:0] _RAND_122;
  reg [31:0] _RAND_123;
  reg [31:0] _RAND_124;
  reg [31:0] _RAND_125;
  reg [31:0] _RAND_126;
  reg [31:0] _RAND_127;
  reg [31:0] _RAND_128;
  reg [31:0] _RAND_129;
  reg [31:0] _RAND_130;
  reg [31:0] _RAND_131;
  reg [31:0] _RAND_132;
  reg [31:0] _RAND_133;
  reg [31:0] _RAND_134;
  reg [31:0] _RAND_135;
  reg [31:0] _RAND_136;
  reg [31:0] _RAND_137;
  reg [31:0] _RAND_138;
  reg [31:0] _RAND_139;
  reg [31:0] _RAND_140;
  reg [31:0] _RAND_141;
  reg [31:0] _RAND_142;
  reg [31:0] _RAND_143;
  reg [31:0] _RAND_144;
  reg [31:0] _RAND_145;
  reg [31:0] _RAND_146;
  reg [31:0] _RAND_147;
  reg [31:0] _RAND_148;
  reg [31:0] _RAND_149;
  reg [31:0] _RAND_150;
  reg [31:0] _RAND_151;
  reg [31:0] _RAND_152;
  reg [31:0] _RAND_153;
  reg [31:0] _RAND_154;
  reg [31:0] _RAND_155;
  reg [31:0] _RAND_156;
  reg [31:0] _RAND_157;
  reg [31:0] _RAND_158;
  reg [31:0] _RAND_159;
  reg [31:0] _RAND_160;
  reg [31:0] _RAND_161;
  reg [31:0] _RAND_162;
  reg [31:0] _RAND_163;
  reg [31:0] _RAND_164;
  reg [31:0] _RAND_165;
  reg [31:0] _RAND_166;
  reg [31:0] _RAND_167;
  reg [31:0] _RAND_168;
  reg [31:0] _RAND_169;
  reg [31:0] _RAND_170;
  reg [31:0] _RAND_171;
  reg [31:0] _RAND_172;
  reg [31:0] _RAND_173;
  reg [31:0] _RAND_174;
  reg [31:0] _RAND_175;
  reg [31:0] _RAND_176;
  reg [31:0] _RAND_177;
  reg [31:0] _RAND_178;
  reg [31:0] _RAND_179;
`endif // RANDOMIZE_REG_INIT
  wire  tlb_clock; // @[:freechips.rocketchip.system.DefaultRV32Config.fir@176840.4]
  wire  tlb_reset; // @[:freechips.rocketchip.system.DefaultRV32Config.fir@176841.4]
  wire  tlb_io_req_ready; // @[:freechips.rocketchip.system.DefaultRV32Config.fir@176842.4]
  wire  tlb_io_req_valid; // @[:freechips.rocketchip.system.DefaultRV32Config.fir@176842.4]
  wire [31:0] tlb_io_req_bits_vaddr; // @[:freechips.rocketchip.system.DefaultRV32Config.fir@176842.4]
  wire  tlb_io_req_bits_passthrough; // @[:freechips.rocketchip.system.DefaultRV32Config.fir@176842.4]
  wire [1:0] tlb_io_req_bits_size; // @[:freechips.rocketchip.system.DefaultRV32Config.fir@176842.4]
  wire [4:0] tlb_io_req_bits_cmd; // @[:freechips.rocketchip.system.DefaultRV32Config.fir@176842.4]
  wire  tlb_io_resp_miss; // @[:freechips.rocketchip.system.DefaultRV32Config.fir@176842.4]
  wire [31:0] tlb_io_resp_paddr; // @[:freechips.rocketchip.system.DefaultRV32Config.fir@176842.4]
  wire  tlb_io_resp_pf_ld; // @[:freechips.rocketchip.system.DefaultRV32Config.fir@176842.4]
  wire  tlb_io_resp_pf_st; // @[:freechips.rocketchip.system.DefaultRV32Config.fir@176842.4]
  wire  tlb_io_resp_ae_ld; // @[:freechips.rocketchip.system.DefaultRV32Config.fir@176842.4]
  wire  tlb_io_resp_ae_st; // @[:freechips.rocketchip.system.DefaultRV32Config.fir@176842.4]
  wire  tlb_io_resp_ma_ld; // @[:freechips.rocketchip.system.DefaultRV32Config.fir@176842.4]
  wire  tlb_io_resp_ma_st; // @[:freechips.rocketchip.system.DefaultRV32Config.fir@176842.4]
  wire  tlb_io_resp_cacheable; // @[:freechips.rocketchip.system.DefaultRV32Config.fir@176842.4]
  wire  tlb_io_sfence_valid; // @[:freechips.rocketchip.system.DefaultRV32Config.fir@176842.4]
  wire  tlb_io_sfence_bits_rs1; // @[:freechips.rocketchip.system.DefaultRV32Config.fir@176842.4]
  wire  tlb_io_sfence_bits_rs2; // @[:freechips.rocketchip.system.DefaultRV32Config.fir@176842.4]
  wire [31:0] tlb_io_sfence_bits_addr; // @[:freechips.rocketchip.system.DefaultRV32Config.fir@176842.4]
  wire  tlb_io_ptw_req_ready; // @[:freechips.rocketchip.system.DefaultRV32Config.fir@176842.4]
  wire  tlb_io_ptw_req_valid; // @[:freechips.rocketchip.system.DefaultRV32Config.fir@176842.4]
  wire [19:0] tlb_io_ptw_req_bits_bits_addr; // @[:freechips.rocketchip.system.DefaultRV32Config.fir@176842.4]
  wire  tlb_io_ptw_resp_valid; // @[:freechips.rocketchip.system.DefaultRV32Config.fir@176842.4]
  wire  tlb_io_ptw_resp_bits_ae; // @[:freechips.rocketchip.system.DefaultRV32Config.fir@176842.4]
  wire [53:0] tlb_io_ptw_resp_bits_pte_ppn; // @[:freechips.rocketchip.system.DefaultRV32Config.fir@176842.4]
  wire  tlb_io_ptw_resp_bits_pte_d; // @[:freechips.rocketchip.system.DefaultRV32Config.fir@176842.4]
  wire  tlb_io_ptw_resp_bits_pte_a; // @[:freechips.rocketchip.system.DefaultRV32Config.fir@176842.4]
  wire  tlb_io_ptw_resp_bits_pte_g; // @[:freechips.rocketchip.system.DefaultRV32Config.fir@176842.4]
  wire  tlb_io_ptw_resp_bits_pte_u; // @[:freechips.rocketchip.system.DefaultRV32Config.fir@176842.4]
  wire  tlb_io_ptw_resp_bits_pte_x; // @[:freechips.rocketchip.system.DefaultRV32Config.fir@176842.4]
  wire  tlb_io_ptw_resp_bits_pte_w; // @[:freechips.rocketchip.system.DefaultRV32Config.fir@176842.4]
  wire  tlb_io_ptw_resp_bits_pte_r; // @[:freechips.rocketchip.system.DefaultRV32Config.fir@176842.4]
  wire  tlb_io_ptw_resp_bits_pte_v; // @[:freechips.rocketchip.system.DefaultRV32Config.fir@176842.4]
  wire  tlb_io_ptw_resp_bits_level; // @[:freechips.rocketchip.system.DefaultRV32Config.fir@176842.4]
  wire  tlb_io_ptw_resp_bits_homogeneous; // @[:freechips.rocketchip.system.DefaultRV32Config.fir@176842.4]
  wire  tlb_io_ptw_ptbr_mode; // @[:freechips.rocketchip.system.DefaultRV32Config.fir@176842.4]
  wire  tlb_io_ptw_status_debug; // @[:freechips.rocketchip.system.DefaultRV32Config.fir@176842.4]
  wire [1:0] tlb_io_ptw_status_dprv; // @[:freechips.rocketchip.system.DefaultRV32Config.fir@176842.4]
  wire  tlb_io_ptw_status_mxr; // @[:freechips.rocketchip.system.DefaultRV32Config.fir@176842.4]
  wire  tlb_io_ptw_status_sum; // @[:freechips.rocketchip.system.DefaultRV32Config.fir@176842.4]
  wire  tlb_io_ptw_pmp_0_cfg_l; // @[:freechips.rocketchip.system.DefaultRV32Config.fir@176842.4]
  wire [1:0] tlb_io_ptw_pmp_0_cfg_a; // @[:freechips.rocketchip.system.DefaultRV32Config.fir@176842.4]
  wire  tlb_io_ptw_pmp_0_cfg_x; // @[:freechips.rocketchip.system.DefaultRV32Config.fir@176842.4]
  wire  tlb_io_ptw_pmp_0_cfg_w; // @[:freechips.rocketchip.system.DefaultRV32Config.fir@176842.4]
  wire  tlb_io_ptw_pmp_0_cfg_r; // @[:freechips.rocketchip.system.DefaultRV32Config.fir@176842.4]
  wire [29:0] tlb_io_ptw_pmp_0_addr; // @[:freechips.rocketchip.system.DefaultRV32Config.fir@176842.4]
  wire [31:0] tlb_io_ptw_pmp_0_mask; // @[:freechips.rocketchip.system.DefaultRV32Config.fir@176842.4]
  wire  tlb_io_ptw_pmp_1_cfg_l; // @[:freechips.rocketchip.system.DefaultRV32Config.fir@176842.4]
  wire [1:0] tlb_io_ptw_pmp_1_cfg_a; // @[:freechips.rocketchip.system.DefaultRV32Config.fir@176842.4]
  wire  tlb_io_ptw_pmp_1_cfg_x; // @[:freechips.rocketchip.system.DefaultRV32Config.fir@176842.4]
  wire  tlb_io_ptw_pmp_1_cfg_w; // @[:freechips.rocketchip.system.DefaultRV32Config.fir@176842.4]
  wire  tlb_io_ptw_pmp_1_cfg_r; // @[:freechips.rocketchip.system.DefaultRV32Config.fir@176842.4]
  wire [29:0] tlb_io_ptw_pmp_1_addr; // @[:freechips.rocketchip.system.DefaultRV32Config.fir@176842.4]
  wire [31:0] tlb_io_ptw_pmp_1_mask; // @[:freechips.rocketchip.system.DefaultRV32Config.fir@176842.4]
  wire  tlb_io_ptw_pmp_2_cfg_l; // @[:freechips.rocketchip.system.DefaultRV32Config.fir@176842.4]
  wire [1:0] tlb_io_ptw_pmp_2_cfg_a; // @[:freechips.rocketchip.system.DefaultRV32Config.fir@176842.4]
  wire  tlb_io_ptw_pmp_2_cfg_x; // @[:freechips.rocketchip.system.DefaultRV32Config.fir@176842.4]
  wire  tlb_io_ptw_pmp_2_cfg_w; // @[:freechips.rocketchip.system.DefaultRV32Config.fir@176842.4]
  wire  tlb_io_ptw_pmp_2_cfg_r; // @[:freechips.rocketchip.system.DefaultRV32Config.fir@176842.4]
  wire [29:0] tlb_io_ptw_pmp_2_addr; // @[:freechips.rocketchip.system.DefaultRV32Config.fir@176842.4]
  wire [31:0] tlb_io_ptw_pmp_2_mask; // @[:freechips.rocketchip.system.DefaultRV32Config.fir@176842.4]
  wire  tlb_io_ptw_pmp_3_cfg_l; // @[:freechips.rocketchip.system.DefaultRV32Config.fir@176842.4]
  wire [1:0] tlb_io_ptw_pmp_3_cfg_a; // @[:freechips.rocketchip.system.DefaultRV32Config.fir@176842.4]
  wire  tlb_io_ptw_pmp_3_cfg_x; // @[:freechips.rocketchip.system.DefaultRV32Config.fir@176842.4]
  wire  tlb_io_ptw_pmp_3_cfg_w; // @[:freechips.rocketchip.system.DefaultRV32Config.fir@176842.4]
  wire  tlb_io_ptw_pmp_3_cfg_r; // @[:freechips.rocketchip.system.DefaultRV32Config.fir@176842.4]
  wire [29:0] tlb_io_ptw_pmp_3_addr; // @[:freechips.rocketchip.system.DefaultRV32Config.fir@176842.4]
  wire [31:0] tlb_io_ptw_pmp_3_mask; // @[:freechips.rocketchip.system.DefaultRV32Config.fir@176842.4]
  wire  tlb_io_ptw_pmp_4_cfg_l; // @[:freechips.rocketchip.system.DefaultRV32Config.fir@176842.4]
  wire [1:0] tlb_io_ptw_pmp_4_cfg_a; // @[:freechips.rocketchip.system.DefaultRV32Config.fir@176842.4]
  wire  tlb_io_ptw_pmp_4_cfg_x; // @[:freechips.rocketchip.system.DefaultRV32Config.fir@176842.4]
  wire  tlb_io_ptw_pmp_4_cfg_w; // @[:freechips.rocketchip.system.DefaultRV32Config.fir@176842.4]
  wire  tlb_io_ptw_pmp_4_cfg_r; // @[:freechips.rocketchip.system.DefaultRV32Config.fir@176842.4]
  wire [29:0] tlb_io_ptw_pmp_4_addr; // @[:freechips.rocketchip.system.DefaultRV32Config.fir@176842.4]
  wire [31:0] tlb_io_ptw_pmp_4_mask; // @[:freechips.rocketchip.system.DefaultRV32Config.fir@176842.4]
  wire  tlb_io_ptw_pmp_5_cfg_l; // @[:freechips.rocketchip.system.DefaultRV32Config.fir@176842.4]
  wire [1:0] tlb_io_ptw_pmp_5_cfg_a; // @[:freechips.rocketchip.system.DefaultRV32Config.fir@176842.4]
  wire  tlb_io_ptw_pmp_5_cfg_x; // @[:freechips.rocketchip.system.DefaultRV32Config.fir@176842.4]
  wire  tlb_io_ptw_pmp_5_cfg_w; // @[:freechips.rocketchip.system.DefaultRV32Config.fir@176842.4]
  wire  tlb_io_ptw_pmp_5_cfg_r; // @[:freechips.rocketchip.system.DefaultRV32Config.fir@176842.4]
  wire [29:0] tlb_io_ptw_pmp_5_addr; // @[:freechips.rocketchip.system.DefaultRV32Config.fir@176842.4]
  wire [31:0] tlb_io_ptw_pmp_5_mask; // @[:freechips.rocketchip.system.DefaultRV32Config.fir@176842.4]
  wire  tlb_io_ptw_pmp_6_cfg_l; // @[:freechips.rocketchip.system.DefaultRV32Config.fir@176842.4]
  wire [1:0] tlb_io_ptw_pmp_6_cfg_a; // @[:freechips.rocketchip.system.DefaultRV32Config.fir@176842.4]
  wire  tlb_io_ptw_pmp_6_cfg_x; // @[:freechips.rocketchip.system.DefaultRV32Config.fir@176842.4]
  wire  tlb_io_ptw_pmp_6_cfg_w; // @[:freechips.rocketchip.system.DefaultRV32Config.fir@176842.4]
  wire  tlb_io_ptw_pmp_6_cfg_r; // @[:freechips.rocketchip.system.DefaultRV32Config.fir@176842.4]
  wire [29:0] tlb_io_ptw_pmp_6_addr; // @[:freechips.rocketchip.system.DefaultRV32Config.fir@176842.4]
  wire [31:0] tlb_io_ptw_pmp_6_mask; // @[:freechips.rocketchip.system.DefaultRV32Config.fir@176842.4]
  wire  tlb_io_ptw_pmp_7_cfg_l; // @[:freechips.rocketchip.system.DefaultRV32Config.fir@176842.4]
  wire [1:0] tlb_io_ptw_pmp_7_cfg_a; // @[:freechips.rocketchip.system.DefaultRV32Config.fir@176842.4]
  wire  tlb_io_ptw_pmp_7_cfg_x; // @[:freechips.rocketchip.system.DefaultRV32Config.fir@176842.4]
  wire  tlb_io_ptw_pmp_7_cfg_w; // @[:freechips.rocketchip.system.DefaultRV32Config.fir@176842.4]
  wire  tlb_io_ptw_pmp_7_cfg_r; // @[:freechips.rocketchip.system.DefaultRV32Config.fir@176842.4]
  wire [29:0] tlb_io_ptw_pmp_7_addr; // @[:freechips.rocketchip.system.DefaultRV32Config.fir@176842.4]
  wire [31:0] tlb_io_ptw_pmp_7_mask; // @[:freechips.rocketchip.system.DefaultRV32Config.fir@176842.4]
  wire [19:0] tlb_OptimizationBarrier_io_x_ppn; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@176907.4]
  wire  tlb_OptimizationBarrier_io_x_u; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@176907.4]
  wire  tlb_OptimizationBarrier_io_x_ae; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@176907.4]
  wire  tlb_OptimizationBarrier_io_x_sw; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@176907.4]
  wire  tlb_OptimizationBarrier_io_x_sx; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@176907.4]
  wire  tlb_OptimizationBarrier_io_x_sr; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@176907.4]
  wire  tlb_OptimizationBarrier_io_x_pw; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@176907.4]
  wire  tlb_OptimizationBarrier_io_x_px; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@176907.4]
  wire  tlb_OptimizationBarrier_io_x_pr; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@176907.4]
  wire  tlb_OptimizationBarrier_io_x_ppp; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@176907.4]
  wire  tlb_OptimizationBarrier_io_x_pal; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@176907.4]
  wire  tlb_OptimizationBarrier_io_x_paa; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@176907.4]
  wire  tlb_OptimizationBarrier_io_x_eff; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@176907.4]
  wire  tlb_OptimizationBarrier_io_x_c; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@176907.4]
  wire [19:0] tlb_OptimizationBarrier_io_y_ppn; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@176907.4]
  wire  tlb_OptimizationBarrier_io_y_u; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@176907.4]
  wire  tlb_OptimizationBarrier_io_y_ae; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@176907.4]
  wire  tlb_OptimizationBarrier_io_y_sw; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@176907.4]
  wire  tlb_OptimizationBarrier_io_y_sx; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@176907.4]
  wire  tlb_OptimizationBarrier_io_y_sr; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@176907.4]
  wire  tlb_OptimizationBarrier_io_y_pw; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@176907.4]
  wire  tlb_OptimizationBarrier_io_y_px; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@176907.4]
  wire  tlb_OptimizationBarrier_io_y_pr; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@176907.4]
  wire  tlb_OptimizationBarrier_io_y_ppp; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@176907.4]
  wire  tlb_OptimizationBarrier_io_y_pal; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@176907.4]
  wire  tlb_OptimizationBarrier_io_y_paa; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@176907.4]
  wire  tlb_OptimizationBarrier_io_y_eff; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@176907.4]
  wire  tlb_OptimizationBarrier_io_y_c; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@176907.4]
  wire [1:0] tlb_pmp_io_prv; // @[TLB.scala 190:19:freechips.rocketchip.system.DefaultRV32Config.fir@176928.4]
  wire  tlb_pmp_io_pmp_0_cfg_l; // @[TLB.scala 190:19:freechips.rocketchip.system.DefaultRV32Config.fir@176928.4]
  wire [1:0] tlb_pmp_io_pmp_0_cfg_a; // @[TLB.scala 190:19:freechips.rocketchip.system.DefaultRV32Config.fir@176928.4]
  wire  tlb_pmp_io_pmp_0_cfg_x; // @[TLB.scala 190:19:freechips.rocketchip.system.DefaultRV32Config.fir@176928.4]
  wire  tlb_pmp_io_pmp_0_cfg_w; // @[TLB.scala 190:19:freechips.rocketchip.system.DefaultRV32Config.fir@176928.4]
  wire  tlb_pmp_io_pmp_0_cfg_r; // @[TLB.scala 190:19:freechips.rocketchip.system.DefaultRV32Config.fir@176928.4]
  wire [29:0] tlb_pmp_io_pmp_0_addr; // @[TLB.scala 190:19:freechips.rocketchip.system.DefaultRV32Config.fir@176928.4]
  wire [31:0] tlb_pmp_io_pmp_0_mask; // @[TLB.scala 190:19:freechips.rocketchip.system.DefaultRV32Config.fir@176928.4]
  wire  tlb_pmp_io_pmp_1_cfg_l; // @[TLB.scala 190:19:freechips.rocketchip.system.DefaultRV32Config.fir@176928.4]
  wire [1:0] tlb_pmp_io_pmp_1_cfg_a; // @[TLB.scala 190:19:freechips.rocketchip.system.DefaultRV32Config.fir@176928.4]
  wire  tlb_pmp_io_pmp_1_cfg_x; // @[TLB.scala 190:19:freechips.rocketchip.system.DefaultRV32Config.fir@176928.4]
  wire  tlb_pmp_io_pmp_1_cfg_w; // @[TLB.scala 190:19:freechips.rocketchip.system.DefaultRV32Config.fir@176928.4]
  wire  tlb_pmp_io_pmp_1_cfg_r; // @[TLB.scala 190:19:freechips.rocketchip.system.DefaultRV32Config.fir@176928.4]
  wire [29:0] tlb_pmp_io_pmp_1_addr; // @[TLB.scala 190:19:freechips.rocketchip.system.DefaultRV32Config.fir@176928.4]
  wire [31:0] tlb_pmp_io_pmp_1_mask; // @[TLB.scala 190:19:freechips.rocketchip.system.DefaultRV32Config.fir@176928.4]
  wire  tlb_pmp_io_pmp_2_cfg_l; // @[TLB.scala 190:19:freechips.rocketchip.system.DefaultRV32Config.fir@176928.4]
  wire [1:0] tlb_pmp_io_pmp_2_cfg_a; // @[TLB.scala 190:19:freechips.rocketchip.system.DefaultRV32Config.fir@176928.4]
  wire  tlb_pmp_io_pmp_2_cfg_x; // @[TLB.scala 190:19:freechips.rocketchip.system.DefaultRV32Config.fir@176928.4]
  wire  tlb_pmp_io_pmp_2_cfg_w; // @[TLB.scala 190:19:freechips.rocketchip.system.DefaultRV32Config.fir@176928.4]
  wire  tlb_pmp_io_pmp_2_cfg_r; // @[TLB.scala 190:19:freechips.rocketchip.system.DefaultRV32Config.fir@176928.4]
  wire [29:0] tlb_pmp_io_pmp_2_addr; // @[TLB.scala 190:19:freechips.rocketchip.system.DefaultRV32Config.fir@176928.4]
  wire [31:0] tlb_pmp_io_pmp_2_mask; // @[TLB.scala 190:19:freechips.rocketchip.system.DefaultRV32Config.fir@176928.4]
  wire  tlb_pmp_io_pmp_3_cfg_l; // @[TLB.scala 190:19:freechips.rocketchip.system.DefaultRV32Config.fir@176928.4]
  wire [1:0] tlb_pmp_io_pmp_3_cfg_a; // @[TLB.scala 190:19:freechips.rocketchip.system.DefaultRV32Config.fir@176928.4]
  wire  tlb_pmp_io_pmp_3_cfg_x; // @[TLB.scala 190:19:freechips.rocketchip.system.DefaultRV32Config.fir@176928.4]
  wire  tlb_pmp_io_pmp_3_cfg_w; // @[TLB.scala 190:19:freechips.rocketchip.system.DefaultRV32Config.fir@176928.4]
  wire  tlb_pmp_io_pmp_3_cfg_r; // @[TLB.scala 190:19:freechips.rocketchip.system.DefaultRV32Config.fir@176928.4]
  wire [29:0] tlb_pmp_io_pmp_3_addr; // @[TLB.scala 190:19:freechips.rocketchip.system.DefaultRV32Config.fir@176928.4]
  wire [31:0] tlb_pmp_io_pmp_3_mask; // @[TLB.scala 190:19:freechips.rocketchip.system.DefaultRV32Config.fir@176928.4]
  wire  tlb_pmp_io_pmp_4_cfg_l; // @[TLB.scala 190:19:freechips.rocketchip.system.DefaultRV32Config.fir@176928.4]
  wire [1:0] tlb_pmp_io_pmp_4_cfg_a; // @[TLB.scala 190:19:freechips.rocketchip.system.DefaultRV32Config.fir@176928.4]
  wire  tlb_pmp_io_pmp_4_cfg_x; // @[TLB.scala 190:19:freechips.rocketchip.system.DefaultRV32Config.fir@176928.4]
  wire  tlb_pmp_io_pmp_4_cfg_w; // @[TLB.scala 190:19:freechips.rocketchip.system.DefaultRV32Config.fir@176928.4]
  wire  tlb_pmp_io_pmp_4_cfg_r; // @[TLB.scala 190:19:freechips.rocketchip.system.DefaultRV32Config.fir@176928.4]
  wire [29:0] tlb_pmp_io_pmp_4_addr; // @[TLB.scala 190:19:freechips.rocketchip.system.DefaultRV32Config.fir@176928.4]
  wire [31:0] tlb_pmp_io_pmp_4_mask; // @[TLB.scala 190:19:freechips.rocketchip.system.DefaultRV32Config.fir@176928.4]
  wire  tlb_pmp_io_pmp_5_cfg_l; // @[TLB.scala 190:19:freechips.rocketchip.system.DefaultRV32Config.fir@176928.4]
  wire [1:0] tlb_pmp_io_pmp_5_cfg_a; // @[TLB.scala 190:19:freechips.rocketchip.system.DefaultRV32Config.fir@176928.4]
  wire  tlb_pmp_io_pmp_5_cfg_x; // @[TLB.scala 190:19:freechips.rocketchip.system.DefaultRV32Config.fir@176928.4]
  wire  tlb_pmp_io_pmp_5_cfg_w; // @[TLB.scala 190:19:freechips.rocketchip.system.DefaultRV32Config.fir@176928.4]
  wire  tlb_pmp_io_pmp_5_cfg_r; // @[TLB.scala 190:19:freechips.rocketchip.system.DefaultRV32Config.fir@176928.4]
  wire [29:0] tlb_pmp_io_pmp_5_addr; // @[TLB.scala 190:19:freechips.rocketchip.system.DefaultRV32Config.fir@176928.4]
  wire [31:0] tlb_pmp_io_pmp_5_mask; // @[TLB.scala 190:19:freechips.rocketchip.system.DefaultRV32Config.fir@176928.4]
  wire  tlb_pmp_io_pmp_6_cfg_l; // @[TLB.scala 190:19:freechips.rocketchip.system.DefaultRV32Config.fir@176928.4]
  wire [1:0] tlb_pmp_io_pmp_6_cfg_a; // @[TLB.scala 190:19:freechips.rocketchip.system.DefaultRV32Config.fir@176928.4]
  wire  tlb_pmp_io_pmp_6_cfg_x; // @[TLB.scala 190:19:freechips.rocketchip.system.DefaultRV32Config.fir@176928.4]
  wire  tlb_pmp_io_pmp_6_cfg_w; // @[TLB.scala 190:19:freechips.rocketchip.system.DefaultRV32Config.fir@176928.4]
  wire  tlb_pmp_io_pmp_6_cfg_r; // @[TLB.scala 190:19:freechips.rocketchip.system.DefaultRV32Config.fir@176928.4]
  wire [29:0] tlb_pmp_io_pmp_6_addr; // @[TLB.scala 190:19:freechips.rocketchip.system.DefaultRV32Config.fir@176928.4]
  wire [31:0] tlb_pmp_io_pmp_6_mask; // @[TLB.scala 190:19:freechips.rocketchip.system.DefaultRV32Config.fir@176928.4]
  wire  tlb_pmp_io_pmp_7_cfg_l; // @[TLB.scala 190:19:freechips.rocketchip.system.DefaultRV32Config.fir@176928.4]
  wire [1:0] tlb_pmp_io_pmp_7_cfg_a; // @[TLB.scala 190:19:freechips.rocketchip.system.DefaultRV32Config.fir@176928.4]
  wire  tlb_pmp_io_pmp_7_cfg_x; // @[TLB.scala 190:19:freechips.rocketchip.system.DefaultRV32Config.fir@176928.4]
  wire  tlb_pmp_io_pmp_7_cfg_w; // @[TLB.scala 190:19:freechips.rocketchip.system.DefaultRV32Config.fir@176928.4]
  wire  tlb_pmp_io_pmp_7_cfg_r; // @[TLB.scala 190:19:freechips.rocketchip.system.DefaultRV32Config.fir@176928.4]
  wire [29:0] tlb_pmp_io_pmp_7_addr; // @[TLB.scala 190:19:freechips.rocketchip.system.DefaultRV32Config.fir@176928.4]
  wire [31:0] tlb_pmp_io_pmp_7_mask; // @[TLB.scala 190:19:freechips.rocketchip.system.DefaultRV32Config.fir@176928.4]
  wire [31:0] tlb_pmp_io_addr; // @[TLB.scala 190:19:freechips.rocketchip.system.DefaultRV32Config.fir@176928.4]
  wire  tlb_pmp_io_r; // @[TLB.scala 190:19:freechips.rocketchip.system.DefaultRV32Config.fir@176928.4]
  wire  tlb_pmp_io_w; // @[TLB.scala 190:19:freechips.rocketchip.system.DefaultRV32Config.fir@176928.4]
  wire  tlb_pmp_io_x; // @[TLB.scala 190:19:freechips.rocketchip.system.DefaultRV32Config.fir@176928.4]
  wire [19:0] tlb_OptimizationBarrier_1_io_x_ppn; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@177629.4]
  wire  tlb_OptimizationBarrier_1_io_x_u; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@177629.4]
  wire  tlb_OptimizationBarrier_1_io_x_ae; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@177629.4]
  wire  tlb_OptimizationBarrier_1_io_x_sw; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@177629.4]
  wire  tlb_OptimizationBarrier_1_io_x_sx; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@177629.4]
  wire  tlb_OptimizationBarrier_1_io_x_sr; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@177629.4]
  wire  tlb_OptimizationBarrier_1_io_x_pw; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@177629.4]
  wire  tlb_OptimizationBarrier_1_io_x_px; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@177629.4]
  wire  tlb_OptimizationBarrier_1_io_x_pr; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@177629.4]
  wire  tlb_OptimizationBarrier_1_io_x_ppp; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@177629.4]
  wire  tlb_OptimizationBarrier_1_io_x_pal; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@177629.4]
  wire  tlb_OptimizationBarrier_1_io_x_paa; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@177629.4]
  wire  tlb_OptimizationBarrier_1_io_x_eff; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@177629.4]
  wire  tlb_OptimizationBarrier_1_io_x_c; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@177629.4]
  wire [19:0] tlb_OptimizationBarrier_1_io_y_ppn; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@177629.4]
  wire  tlb_OptimizationBarrier_1_io_y_u; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@177629.4]
  wire  tlb_OptimizationBarrier_1_io_y_ae; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@177629.4]
  wire  tlb_OptimizationBarrier_1_io_y_sw; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@177629.4]
  wire  tlb_OptimizationBarrier_1_io_y_sx; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@177629.4]
  wire  tlb_OptimizationBarrier_1_io_y_sr; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@177629.4]
  wire  tlb_OptimizationBarrier_1_io_y_pw; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@177629.4]
  wire  tlb_OptimizationBarrier_1_io_y_px; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@177629.4]
  wire  tlb_OptimizationBarrier_1_io_y_pr; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@177629.4]
  wire  tlb_OptimizationBarrier_1_io_y_ppp; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@177629.4]
  wire  tlb_OptimizationBarrier_1_io_y_pal; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@177629.4]
  wire  tlb_OptimizationBarrier_1_io_y_paa; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@177629.4]
  wire  tlb_OptimizationBarrier_1_io_y_eff; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@177629.4]
  wire  tlb_OptimizationBarrier_1_io_y_c; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@177629.4]
  wire [19:0] tlb_OptimizationBarrier_2_io_x_ppn; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@177672.4]
  wire  tlb_OptimizationBarrier_2_io_x_u; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@177672.4]
  wire  tlb_OptimizationBarrier_2_io_x_ae; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@177672.4]
  wire  tlb_OptimizationBarrier_2_io_x_sw; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@177672.4]
  wire  tlb_OptimizationBarrier_2_io_x_sx; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@177672.4]
  wire  tlb_OptimizationBarrier_2_io_x_sr; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@177672.4]
  wire  tlb_OptimizationBarrier_2_io_x_pw; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@177672.4]
  wire  tlb_OptimizationBarrier_2_io_x_px; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@177672.4]
  wire  tlb_OptimizationBarrier_2_io_x_pr; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@177672.4]
  wire  tlb_OptimizationBarrier_2_io_x_ppp; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@177672.4]
  wire  tlb_OptimizationBarrier_2_io_x_pal; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@177672.4]
  wire  tlb_OptimizationBarrier_2_io_x_paa; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@177672.4]
  wire  tlb_OptimizationBarrier_2_io_x_eff; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@177672.4]
  wire  tlb_OptimizationBarrier_2_io_x_c; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@177672.4]
  wire [19:0] tlb_OptimizationBarrier_2_io_y_ppn; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@177672.4]
  wire  tlb_OptimizationBarrier_2_io_y_u; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@177672.4]
  wire  tlb_OptimizationBarrier_2_io_y_ae; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@177672.4]
  wire  tlb_OptimizationBarrier_2_io_y_sw; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@177672.4]
  wire  tlb_OptimizationBarrier_2_io_y_sx; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@177672.4]
  wire  tlb_OptimizationBarrier_2_io_y_sr; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@177672.4]
  wire  tlb_OptimizationBarrier_2_io_y_pw; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@177672.4]
  wire  tlb_OptimizationBarrier_2_io_y_px; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@177672.4]
  wire  tlb_OptimizationBarrier_2_io_y_pr; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@177672.4]
  wire  tlb_OptimizationBarrier_2_io_y_ppp; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@177672.4]
  wire  tlb_OptimizationBarrier_2_io_y_pal; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@177672.4]
  wire  tlb_OptimizationBarrier_2_io_y_paa; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@177672.4]
  wire  tlb_OptimizationBarrier_2_io_y_eff; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@177672.4]
  wire  tlb_OptimizationBarrier_2_io_y_c; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@177672.4]
  wire [19:0] tlb_OptimizationBarrier_3_io_x_ppn; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@177715.4]
  wire  tlb_OptimizationBarrier_3_io_x_u; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@177715.4]
  wire  tlb_OptimizationBarrier_3_io_x_ae; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@177715.4]
  wire  tlb_OptimizationBarrier_3_io_x_sw; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@177715.4]
  wire  tlb_OptimizationBarrier_3_io_x_sx; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@177715.4]
  wire  tlb_OptimizationBarrier_3_io_x_sr; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@177715.4]
  wire  tlb_OptimizationBarrier_3_io_x_pw; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@177715.4]
  wire  tlb_OptimizationBarrier_3_io_x_px; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@177715.4]
  wire  tlb_OptimizationBarrier_3_io_x_pr; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@177715.4]
  wire  tlb_OptimizationBarrier_3_io_x_ppp; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@177715.4]
  wire  tlb_OptimizationBarrier_3_io_x_pal; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@177715.4]
  wire  tlb_OptimizationBarrier_3_io_x_paa; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@177715.4]
  wire  tlb_OptimizationBarrier_3_io_x_eff; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@177715.4]
  wire  tlb_OptimizationBarrier_3_io_x_c; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@177715.4]
  wire [19:0] tlb_OptimizationBarrier_3_io_y_ppn; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@177715.4]
  wire  tlb_OptimizationBarrier_3_io_y_u; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@177715.4]
  wire  tlb_OptimizationBarrier_3_io_y_ae; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@177715.4]
  wire  tlb_OptimizationBarrier_3_io_y_sw; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@177715.4]
  wire  tlb_OptimizationBarrier_3_io_y_sx; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@177715.4]
  wire  tlb_OptimizationBarrier_3_io_y_sr; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@177715.4]
  wire  tlb_OptimizationBarrier_3_io_y_pw; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@177715.4]
  wire  tlb_OptimizationBarrier_3_io_y_px; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@177715.4]
  wire  tlb_OptimizationBarrier_3_io_y_pr; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@177715.4]
  wire  tlb_OptimizationBarrier_3_io_y_ppp; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@177715.4]
  wire  tlb_OptimizationBarrier_3_io_y_pal; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@177715.4]
  wire  tlb_OptimizationBarrier_3_io_y_paa; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@177715.4]
  wire  tlb_OptimizationBarrier_3_io_y_eff; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@177715.4]
  wire  tlb_OptimizationBarrier_3_io_y_c; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@177715.4]
  wire [19:0] tlb_OptimizationBarrier_4_io_x_ppn; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@177758.4]
  wire  tlb_OptimizationBarrier_4_io_x_u; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@177758.4]
  wire  tlb_OptimizationBarrier_4_io_x_ae; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@177758.4]
  wire  tlb_OptimizationBarrier_4_io_x_sw; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@177758.4]
  wire  tlb_OptimizationBarrier_4_io_x_sx; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@177758.4]
  wire  tlb_OptimizationBarrier_4_io_x_sr; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@177758.4]
  wire  tlb_OptimizationBarrier_4_io_x_pw; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@177758.4]
  wire  tlb_OptimizationBarrier_4_io_x_px; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@177758.4]
  wire  tlb_OptimizationBarrier_4_io_x_pr; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@177758.4]
  wire  tlb_OptimizationBarrier_4_io_x_ppp; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@177758.4]
  wire  tlb_OptimizationBarrier_4_io_x_pal; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@177758.4]
  wire  tlb_OptimizationBarrier_4_io_x_paa; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@177758.4]
  wire  tlb_OptimizationBarrier_4_io_x_eff; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@177758.4]
  wire  tlb_OptimizationBarrier_4_io_x_c; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@177758.4]
  wire [19:0] tlb_OptimizationBarrier_4_io_y_ppn; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@177758.4]
  wire  tlb_OptimizationBarrier_4_io_y_u; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@177758.4]
  wire  tlb_OptimizationBarrier_4_io_y_ae; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@177758.4]
  wire  tlb_OptimizationBarrier_4_io_y_sw; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@177758.4]
  wire  tlb_OptimizationBarrier_4_io_y_sx; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@177758.4]
  wire  tlb_OptimizationBarrier_4_io_y_sr; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@177758.4]
  wire  tlb_OptimizationBarrier_4_io_y_pw; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@177758.4]
  wire  tlb_OptimizationBarrier_4_io_y_px; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@177758.4]
  wire  tlb_OptimizationBarrier_4_io_y_pr; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@177758.4]
  wire  tlb_OptimizationBarrier_4_io_y_ppp; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@177758.4]
  wire  tlb_OptimizationBarrier_4_io_y_pal; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@177758.4]
  wire  tlb_OptimizationBarrier_4_io_y_paa; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@177758.4]
  wire  tlb_OptimizationBarrier_4_io_y_eff; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@177758.4]
  wire  tlb_OptimizationBarrier_4_io_y_c; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@177758.4]
  wire [19:0] tlb_OptimizationBarrier_5_io_x_ppn; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@177801.4]
  wire  tlb_OptimizationBarrier_5_io_x_u; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@177801.4]
  wire  tlb_OptimizationBarrier_5_io_x_ae; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@177801.4]
  wire  tlb_OptimizationBarrier_5_io_x_sw; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@177801.4]
  wire  tlb_OptimizationBarrier_5_io_x_sx; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@177801.4]
  wire  tlb_OptimizationBarrier_5_io_x_sr; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@177801.4]
  wire  tlb_OptimizationBarrier_5_io_x_pw; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@177801.4]
  wire  tlb_OptimizationBarrier_5_io_x_px; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@177801.4]
  wire  tlb_OptimizationBarrier_5_io_x_pr; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@177801.4]
  wire  tlb_OptimizationBarrier_5_io_x_ppp; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@177801.4]
  wire  tlb_OptimizationBarrier_5_io_x_pal; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@177801.4]
  wire  tlb_OptimizationBarrier_5_io_x_paa; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@177801.4]
  wire  tlb_OptimizationBarrier_5_io_x_eff; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@177801.4]
  wire  tlb_OptimizationBarrier_5_io_x_c; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@177801.4]
  wire [19:0] tlb_OptimizationBarrier_5_io_y_ppn; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@177801.4]
  wire  tlb_OptimizationBarrier_5_io_y_u; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@177801.4]
  wire  tlb_OptimizationBarrier_5_io_y_ae; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@177801.4]
  wire  tlb_OptimizationBarrier_5_io_y_sw; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@177801.4]
  wire  tlb_OptimizationBarrier_5_io_y_sx; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@177801.4]
  wire  tlb_OptimizationBarrier_5_io_y_sr; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@177801.4]
  wire  tlb_OptimizationBarrier_5_io_y_pw; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@177801.4]
  wire  tlb_OptimizationBarrier_5_io_y_px; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@177801.4]
  wire  tlb_OptimizationBarrier_5_io_y_pr; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@177801.4]
  wire  tlb_OptimizationBarrier_5_io_y_ppp; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@177801.4]
  wire  tlb_OptimizationBarrier_5_io_y_pal; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@177801.4]
  wire  tlb_OptimizationBarrier_5_io_y_paa; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@177801.4]
  wire  tlb_OptimizationBarrier_5_io_y_eff; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@177801.4]
  wire  tlb_OptimizationBarrier_5_io_y_c; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@177801.4]
  wire [19:0] tlb_OptimizationBarrier_6_io_x_ppn; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@177844.4]
  wire  tlb_OptimizationBarrier_6_io_x_u; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@177844.4]
  wire  tlb_OptimizationBarrier_6_io_x_ae; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@177844.4]
  wire  tlb_OptimizationBarrier_6_io_x_sw; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@177844.4]
  wire  tlb_OptimizationBarrier_6_io_x_sx; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@177844.4]
  wire  tlb_OptimizationBarrier_6_io_x_sr; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@177844.4]
  wire  tlb_OptimizationBarrier_6_io_x_pw; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@177844.4]
  wire  tlb_OptimizationBarrier_6_io_x_px; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@177844.4]
  wire  tlb_OptimizationBarrier_6_io_x_pr; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@177844.4]
  wire  tlb_OptimizationBarrier_6_io_x_ppp; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@177844.4]
  wire  tlb_OptimizationBarrier_6_io_x_pal; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@177844.4]
  wire  tlb_OptimizationBarrier_6_io_x_paa; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@177844.4]
  wire  tlb_OptimizationBarrier_6_io_x_eff; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@177844.4]
  wire  tlb_OptimizationBarrier_6_io_x_c; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@177844.4]
  wire [19:0] tlb_OptimizationBarrier_6_io_y_ppn; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@177844.4]
  wire  tlb_OptimizationBarrier_6_io_y_u; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@177844.4]
  wire  tlb_OptimizationBarrier_6_io_y_ae; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@177844.4]
  wire  tlb_OptimizationBarrier_6_io_y_sw; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@177844.4]
  wire  tlb_OptimizationBarrier_6_io_y_sx; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@177844.4]
  wire  tlb_OptimizationBarrier_6_io_y_sr; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@177844.4]
  wire  tlb_OptimizationBarrier_6_io_y_pw; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@177844.4]
  wire  tlb_OptimizationBarrier_6_io_y_px; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@177844.4]
  wire  tlb_OptimizationBarrier_6_io_y_pr; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@177844.4]
  wire  tlb_OptimizationBarrier_6_io_y_ppp; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@177844.4]
  wire  tlb_OptimizationBarrier_6_io_y_pal; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@177844.4]
  wire  tlb_OptimizationBarrier_6_io_y_paa; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@177844.4]
  wire  tlb_OptimizationBarrier_6_io_y_eff; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@177844.4]
  wire  tlb_OptimizationBarrier_6_io_y_c; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@177844.4]
  wire [19:0] tlb_OptimizationBarrier_7_io_x_ppn; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@177887.4]
  wire  tlb_OptimizationBarrier_7_io_x_u; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@177887.4]
  wire  tlb_OptimizationBarrier_7_io_x_ae; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@177887.4]
  wire  tlb_OptimizationBarrier_7_io_x_sw; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@177887.4]
  wire  tlb_OptimizationBarrier_7_io_x_sx; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@177887.4]
  wire  tlb_OptimizationBarrier_7_io_x_sr; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@177887.4]
  wire  tlb_OptimizationBarrier_7_io_x_pw; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@177887.4]
  wire  tlb_OptimizationBarrier_7_io_x_px; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@177887.4]
  wire  tlb_OptimizationBarrier_7_io_x_pr; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@177887.4]
  wire  tlb_OptimizationBarrier_7_io_x_ppp; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@177887.4]
  wire  tlb_OptimizationBarrier_7_io_x_pal; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@177887.4]
  wire  tlb_OptimizationBarrier_7_io_x_paa; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@177887.4]
  wire  tlb_OptimizationBarrier_7_io_x_eff; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@177887.4]
  wire  tlb_OptimizationBarrier_7_io_x_c; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@177887.4]
  wire [19:0] tlb_OptimizationBarrier_7_io_y_ppn; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@177887.4]
  wire  tlb_OptimizationBarrier_7_io_y_u; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@177887.4]
  wire  tlb_OptimizationBarrier_7_io_y_ae; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@177887.4]
  wire  tlb_OptimizationBarrier_7_io_y_sw; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@177887.4]
  wire  tlb_OptimizationBarrier_7_io_y_sx; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@177887.4]
  wire  tlb_OptimizationBarrier_7_io_y_sr; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@177887.4]
  wire  tlb_OptimizationBarrier_7_io_y_pw; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@177887.4]
  wire  tlb_OptimizationBarrier_7_io_y_px; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@177887.4]
  wire  tlb_OptimizationBarrier_7_io_y_pr; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@177887.4]
  wire  tlb_OptimizationBarrier_7_io_y_ppp; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@177887.4]
  wire  tlb_OptimizationBarrier_7_io_y_pal; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@177887.4]
  wire  tlb_OptimizationBarrier_7_io_y_paa; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@177887.4]
  wire  tlb_OptimizationBarrier_7_io_y_eff; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@177887.4]
  wire  tlb_OptimizationBarrier_7_io_y_c; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@177887.4]
  wire [19:0] tlb_OptimizationBarrier_8_io_x_ppn; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@177930.4]
  wire  tlb_OptimizationBarrier_8_io_x_u; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@177930.4]
  wire  tlb_OptimizationBarrier_8_io_x_ae; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@177930.4]
  wire  tlb_OptimizationBarrier_8_io_x_sw; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@177930.4]
  wire  tlb_OptimizationBarrier_8_io_x_sx; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@177930.4]
  wire  tlb_OptimizationBarrier_8_io_x_sr; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@177930.4]
  wire  tlb_OptimizationBarrier_8_io_x_pw; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@177930.4]
  wire  tlb_OptimizationBarrier_8_io_x_px; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@177930.4]
  wire  tlb_OptimizationBarrier_8_io_x_pr; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@177930.4]
  wire  tlb_OptimizationBarrier_8_io_x_ppp; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@177930.4]
  wire  tlb_OptimizationBarrier_8_io_x_pal; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@177930.4]
  wire  tlb_OptimizationBarrier_8_io_x_paa; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@177930.4]
  wire  tlb_OptimizationBarrier_8_io_x_eff; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@177930.4]
  wire  tlb_OptimizationBarrier_8_io_x_c; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@177930.4]
  wire [19:0] tlb_OptimizationBarrier_8_io_y_ppn; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@177930.4]
  wire  tlb_OptimizationBarrier_8_io_y_u; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@177930.4]
  wire  tlb_OptimizationBarrier_8_io_y_ae; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@177930.4]
  wire  tlb_OptimizationBarrier_8_io_y_sw; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@177930.4]
  wire  tlb_OptimizationBarrier_8_io_y_sx; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@177930.4]
  wire  tlb_OptimizationBarrier_8_io_y_sr; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@177930.4]
  wire  tlb_OptimizationBarrier_8_io_y_pw; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@177930.4]
  wire  tlb_OptimizationBarrier_8_io_y_px; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@177930.4]
  wire  tlb_OptimizationBarrier_8_io_y_pr; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@177930.4]
  wire  tlb_OptimizationBarrier_8_io_y_ppp; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@177930.4]
  wire  tlb_OptimizationBarrier_8_io_y_pal; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@177930.4]
  wire  tlb_OptimizationBarrier_8_io_y_paa; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@177930.4]
  wire  tlb_OptimizationBarrier_8_io_y_eff; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@177930.4]
  wire  tlb_OptimizationBarrier_8_io_y_c; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@177930.4]
  wire [19:0] tlb_OptimizationBarrier_9_io_x_ppn; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@177972.4]
  wire  tlb_OptimizationBarrier_9_io_x_u; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@177972.4]
  wire  tlb_OptimizationBarrier_9_io_x_ae; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@177972.4]
  wire  tlb_OptimizationBarrier_9_io_x_sw; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@177972.4]
  wire  tlb_OptimizationBarrier_9_io_x_sx; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@177972.4]
  wire  tlb_OptimizationBarrier_9_io_x_sr; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@177972.4]
  wire  tlb_OptimizationBarrier_9_io_x_pw; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@177972.4]
  wire  tlb_OptimizationBarrier_9_io_x_px; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@177972.4]
  wire  tlb_OptimizationBarrier_9_io_x_pr; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@177972.4]
  wire  tlb_OptimizationBarrier_9_io_x_ppp; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@177972.4]
  wire  tlb_OptimizationBarrier_9_io_x_pal; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@177972.4]
  wire  tlb_OptimizationBarrier_9_io_x_paa; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@177972.4]
  wire  tlb_OptimizationBarrier_9_io_x_eff; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@177972.4]
  wire  tlb_OptimizationBarrier_9_io_x_c; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@177972.4]
  wire [19:0] tlb_OptimizationBarrier_9_io_y_ppn; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@177972.4]
  wire  tlb_OptimizationBarrier_9_io_y_u; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@177972.4]
  wire  tlb_OptimizationBarrier_9_io_y_ae; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@177972.4]
  wire  tlb_OptimizationBarrier_9_io_y_sw; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@177972.4]
  wire  tlb_OptimizationBarrier_9_io_y_sx; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@177972.4]
  wire  tlb_OptimizationBarrier_9_io_y_sr; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@177972.4]
  wire  tlb_OptimizationBarrier_9_io_y_pw; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@177972.4]
  wire  tlb_OptimizationBarrier_9_io_y_px; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@177972.4]
  wire  tlb_OptimizationBarrier_9_io_y_pr; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@177972.4]
  wire  tlb_OptimizationBarrier_9_io_y_ppp; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@177972.4]
  wire  tlb_OptimizationBarrier_9_io_y_pal; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@177972.4]
  wire  tlb_OptimizationBarrier_9_io_y_paa; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@177972.4]
  wire  tlb_OptimizationBarrier_9_io_y_eff; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@177972.4]
  wire  tlb_OptimizationBarrier_9_io_y_c; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@177972.4]
  wire [19:0] tlb_OptimizationBarrier_10_io_x_ppn; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178021.4]
  wire  tlb_OptimizationBarrier_10_io_x_u; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178021.4]
  wire  tlb_OptimizationBarrier_10_io_x_ae; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178021.4]
  wire  tlb_OptimizationBarrier_10_io_x_sw; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178021.4]
  wire  tlb_OptimizationBarrier_10_io_x_sx; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178021.4]
  wire  tlb_OptimizationBarrier_10_io_x_sr; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178021.4]
  wire  tlb_OptimizationBarrier_10_io_x_pw; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178021.4]
  wire  tlb_OptimizationBarrier_10_io_x_px; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178021.4]
  wire  tlb_OptimizationBarrier_10_io_x_pr; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178021.4]
  wire  tlb_OptimizationBarrier_10_io_x_ppp; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178021.4]
  wire  tlb_OptimizationBarrier_10_io_x_pal; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178021.4]
  wire  tlb_OptimizationBarrier_10_io_x_paa; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178021.4]
  wire  tlb_OptimizationBarrier_10_io_x_eff; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178021.4]
  wire  tlb_OptimizationBarrier_10_io_x_c; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178021.4]
  wire [19:0] tlb_OptimizationBarrier_10_io_y_ppn; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178021.4]
  wire  tlb_OptimizationBarrier_10_io_y_u; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178021.4]
  wire  tlb_OptimizationBarrier_10_io_y_ae; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178021.4]
  wire  tlb_OptimizationBarrier_10_io_y_sw; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178021.4]
  wire  tlb_OptimizationBarrier_10_io_y_sx; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178021.4]
  wire  tlb_OptimizationBarrier_10_io_y_sr; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178021.4]
  wire  tlb_OptimizationBarrier_10_io_y_pw; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178021.4]
  wire  tlb_OptimizationBarrier_10_io_y_px; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178021.4]
  wire  tlb_OptimizationBarrier_10_io_y_pr; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178021.4]
  wire  tlb_OptimizationBarrier_10_io_y_ppp; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178021.4]
  wire  tlb_OptimizationBarrier_10_io_y_pal; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178021.4]
  wire  tlb_OptimizationBarrier_10_io_y_paa; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178021.4]
  wire  tlb_OptimizationBarrier_10_io_y_eff; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178021.4]
  wire  tlb_OptimizationBarrier_10_io_y_c; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178021.4]
  wire [19:0] tlb_OptimizationBarrier_11_io_x_ppn; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178070.4]
  wire  tlb_OptimizationBarrier_11_io_x_u; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178070.4]
  wire  tlb_OptimizationBarrier_11_io_x_ae; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178070.4]
  wire  tlb_OptimizationBarrier_11_io_x_sw; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178070.4]
  wire  tlb_OptimizationBarrier_11_io_x_sx; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178070.4]
  wire  tlb_OptimizationBarrier_11_io_x_sr; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178070.4]
  wire  tlb_OptimizationBarrier_11_io_x_pw; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178070.4]
  wire  tlb_OptimizationBarrier_11_io_x_px; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178070.4]
  wire  tlb_OptimizationBarrier_11_io_x_pr; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178070.4]
  wire  tlb_OptimizationBarrier_11_io_x_ppp; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178070.4]
  wire  tlb_OptimizationBarrier_11_io_x_pal; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178070.4]
  wire  tlb_OptimizationBarrier_11_io_x_paa; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178070.4]
  wire  tlb_OptimizationBarrier_11_io_x_eff; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178070.4]
  wire  tlb_OptimizationBarrier_11_io_x_c; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178070.4]
  wire [19:0] tlb_OptimizationBarrier_11_io_y_ppn; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178070.4]
  wire  tlb_OptimizationBarrier_11_io_y_u; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178070.4]
  wire  tlb_OptimizationBarrier_11_io_y_ae; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178070.4]
  wire  tlb_OptimizationBarrier_11_io_y_sw; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178070.4]
  wire  tlb_OptimizationBarrier_11_io_y_sx; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178070.4]
  wire  tlb_OptimizationBarrier_11_io_y_sr; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178070.4]
  wire  tlb_OptimizationBarrier_11_io_y_pw; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178070.4]
  wire  tlb_OptimizationBarrier_11_io_y_px; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178070.4]
  wire  tlb_OptimizationBarrier_11_io_y_pr; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178070.4]
  wire  tlb_OptimizationBarrier_11_io_y_ppp; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178070.4]
  wire  tlb_OptimizationBarrier_11_io_y_pal; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178070.4]
  wire  tlb_OptimizationBarrier_11_io_y_paa; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178070.4]
  wire  tlb_OptimizationBarrier_11_io_y_eff; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178070.4]
  wire  tlb_OptimizationBarrier_11_io_y_c; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178070.4]
  wire [19:0] tlb_OptimizationBarrier_12_io_x_ppn; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178119.4]
  wire  tlb_OptimizationBarrier_12_io_x_u; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178119.4]
  wire  tlb_OptimizationBarrier_12_io_x_ae; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178119.4]
  wire  tlb_OptimizationBarrier_12_io_x_sw; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178119.4]
  wire  tlb_OptimizationBarrier_12_io_x_sx; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178119.4]
  wire  tlb_OptimizationBarrier_12_io_x_sr; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178119.4]
  wire  tlb_OptimizationBarrier_12_io_x_pw; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178119.4]
  wire  tlb_OptimizationBarrier_12_io_x_px; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178119.4]
  wire  tlb_OptimizationBarrier_12_io_x_pr; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178119.4]
  wire  tlb_OptimizationBarrier_12_io_x_ppp; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178119.4]
  wire  tlb_OptimizationBarrier_12_io_x_pal; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178119.4]
  wire  tlb_OptimizationBarrier_12_io_x_paa; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178119.4]
  wire  tlb_OptimizationBarrier_12_io_x_eff; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178119.4]
  wire  tlb_OptimizationBarrier_12_io_x_c; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178119.4]
  wire [19:0] tlb_OptimizationBarrier_12_io_y_ppn; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178119.4]
  wire  tlb_OptimizationBarrier_12_io_y_u; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178119.4]
  wire  tlb_OptimizationBarrier_12_io_y_ae; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178119.4]
  wire  tlb_OptimizationBarrier_12_io_y_sw; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178119.4]
  wire  tlb_OptimizationBarrier_12_io_y_sx; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178119.4]
  wire  tlb_OptimizationBarrier_12_io_y_sr; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178119.4]
  wire  tlb_OptimizationBarrier_12_io_y_pw; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178119.4]
  wire  tlb_OptimizationBarrier_12_io_y_px; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178119.4]
  wire  tlb_OptimizationBarrier_12_io_y_pr; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178119.4]
  wire  tlb_OptimizationBarrier_12_io_y_ppp; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178119.4]
  wire  tlb_OptimizationBarrier_12_io_y_pal; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178119.4]
  wire  tlb_OptimizationBarrier_12_io_y_paa; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178119.4]
  wire  tlb_OptimizationBarrier_12_io_y_eff; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178119.4]
  wire  tlb_OptimizationBarrier_12_io_y_c; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178119.4]
  wire [19:0] tlb_OptimizationBarrier_13_io_x_ppn; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178168.4]
  wire  tlb_OptimizationBarrier_13_io_x_u; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178168.4]
  wire  tlb_OptimizationBarrier_13_io_x_ae; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178168.4]
  wire  tlb_OptimizationBarrier_13_io_x_sw; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178168.4]
  wire  tlb_OptimizationBarrier_13_io_x_sx; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178168.4]
  wire  tlb_OptimizationBarrier_13_io_x_sr; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178168.4]
  wire  tlb_OptimizationBarrier_13_io_x_pw; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178168.4]
  wire  tlb_OptimizationBarrier_13_io_x_px; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178168.4]
  wire  tlb_OptimizationBarrier_13_io_x_pr; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178168.4]
  wire  tlb_OptimizationBarrier_13_io_x_ppp; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178168.4]
  wire  tlb_OptimizationBarrier_13_io_x_pal; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178168.4]
  wire  tlb_OptimizationBarrier_13_io_x_paa; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178168.4]
  wire  tlb_OptimizationBarrier_13_io_x_eff; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178168.4]
  wire  tlb_OptimizationBarrier_13_io_x_c; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178168.4]
  wire [19:0] tlb_OptimizationBarrier_13_io_y_ppn; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178168.4]
  wire  tlb_OptimizationBarrier_13_io_y_u; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178168.4]
  wire  tlb_OptimizationBarrier_13_io_y_ae; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178168.4]
  wire  tlb_OptimizationBarrier_13_io_y_sw; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178168.4]
  wire  tlb_OptimizationBarrier_13_io_y_sx; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178168.4]
  wire  tlb_OptimizationBarrier_13_io_y_sr; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178168.4]
  wire  tlb_OptimizationBarrier_13_io_y_pw; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178168.4]
  wire  tlb_OptimizationBarrier_13_io_y_px; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178168.4]
  wire  tlb_OptimizationBarrier_13_io_y_pr; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178168.4]
  wire  tlb_OptimizationBarrier_13_io_y_ppp; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178168.4]
  wire  tlb_OptimizationBarrier_13_io_y_pal; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178168.4]
  wire  tlb_OptimizationBarrier_13_io_y_paa; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178168.4]
  wire  tlb_OptimizationBarrier_13_io_y_eff; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178168.4]
  wire  tlb_OptimizationBarrier_13_io_y_c; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178168.4]
  wire [19:0] tlb_OptimizationBarrier_14_io_x_ppn; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178649.4]
  wire  tlb_OptimizationBarrier_14_io_x_u; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178649.4]
  wire  tlb_OptimizationBarrier_14_io_x_ae; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178649.4]
  wire  tlb_OptimizationBarrier_14_io_x_sw; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178649.4]
  wire  tlb_OptimizationBarrier_14_io_x_sx; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178649.4]
  wire  tlb_OptimizationBarrier_14_io_x_sr; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178649.4]
  wire  tlb_OptimizationBarrier_14_io_x_pw; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178649.4]
  wire  tlb_OptimizationBarrier_14_io_x_px; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178649.4]
  wire  tlb_OptimizationBarrier_14_io_x_pr; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178649.4]
  wire  tlb_OptimizationBarrier_14_io_x_ppp; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178649.4]
  wire  tlb_OptimizationBarrier_14_io_x_pal; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178649.4]
  wire  tlb_OptimizationBarrier_14_io_x_paa; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178649.4]
  wire  tlb_OptimizationBarrier_14_io_x_eff; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178649.4]
  wire  tlb_OptimizationBarrier_14_io_x_c; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178649.4]
  wire [19:0] tlb_OptimizationBarrier_14_io_y_ppn; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178649.4]
  wire  tlb_OptimizationBarrier_14_io_y_u; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178649.4]
  wire  tlb_OptimizationBarrier_14_io_y_ae; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178649.4]
  wire  tlb_OptimizationBarrier_14_io_y_sw; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178649.4]
  wire  tlb_OptimizationBarrier_14_io_y_sx; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178649.4]
  wire  tlb_OptimizationBarrier_14_io_y_sr; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178649.4]
  wire  tlb_OptimizationBarrier_14_io_y_pw; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178649.4]
  wire  tlb_OptimizationBarrier_14_io_y_px; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178649.4]
  wire  tlb_OptimizationBarrier_14_io_y_pr; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178649.4]
  wire  tlb_OptimizationBarrier_14_io_y_ppp; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178649.4]
  wire  tlb_OptimizationBarrier_14_io_y_pal; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178649.4]
  wire  tlb_OptimizationBarrier_14_io_y_paa; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178649.4]
  wire  tlb_OptimizationBarrier_14_io_y_eff; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178649.4]
  wire  tlb_OptimizationBarrier_14_io_y_c; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178649.4]
  wire [19:0] tlb_OptimizationBarrier_15_io_x_ppn; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178692.4]
  wire  tlb_OptimizationBarrier_15_io_x_u; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178692.4]
  wire  tlb_OptimizationBarrier_15_io_x_ae; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178692.4]
  wire  tlb_OptimizationBarrier_15_io_x_sw; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178692.4]
  wire  tlb_OptimizationBarrier_15_io_x_sx; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178692.4]
  wire  tlb_OptimizationBarrier_15_io_x_sr; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178692.4]
  wire  tlb_OptimizationBarrier_15_io_x_pw; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178692.4]
  wire  tlb_OptimizationBarrier_15_io_x_px; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178692.4]
  wire  tlb_OptimizationBarrier_15_io_x_pr; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178692.4]
  wire  tlb_OptimizationBarrier_15_io_x_ppp; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178692.4]
  wire  tlb_OptimizationBarrier_15_io_x_pal; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178692.4]
  wire  tlb_OptimizationBarrier_15_io_x_paa; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178692.4]
  wire  tlb_OptimizationBarrier_15_io_x_eff; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178692.4]
  wire  tlb_OptimizationBarrier_15_io_x_c; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178692.4]
  wire [19:0] tlb_OptimizationBarrier_15_io_y_ppn; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178692.4]
  wire  tlb_OptimizationBarrier_15_io_y_u; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178692.4]
  wire  tlb_OptimizationBarrier_15_io_y_ae; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178692.4]
  wire  tlb_OptimizationBarrier_15_io_y_sw; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178692.4]
  wire  tlb_OptimizationBarrier_15_io_y_sx; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178692.4]
  wire  tlb_OptimizationBarrier_15_io_y_sr; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178692.4]
  wire  tlb_OptimizationBarrier_15_io_y_pw; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178692.4]
  wire  tlb_OptimizationBarrier_15_io_y_px; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178692.4]
  wire  tlb_OptimizationBarrier_15_io_y_pr; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178692.4]
  wire  tlb_OptimizationBarrier_15_io_y_ppp; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178692.4]
  wire  tlb_OptimizationBarrier_15_io_y_pal; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178692.4]
  wire  tlb_OptimizationBarrier_15_io_y_paa; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178692.4]
  wire  tlb_OptimizationBarrier_15_io_y_eff; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178692.4]
  wire  tlb_OptimizationBarrier_15_io_y_c; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178692.4]
  wire [19:0] tlb_OptimizationBarrier_16_io_x_ppn; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178735.4]
  wire  tlb_OptimizationBarrier_16_io_x_u; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178735.4]
  wire  tlb_OptimizationBarrier_16_io_x_ae; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178735.4]
  wire  tlb_OptimizationBarrier_16_io_x_sw; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178735.4]
  wire  tlb_OptimizationBarrier_16_io_x_sx; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178735.4]
  wire  tlb_OptimizationBarrier_16_io_x_sr; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178735.4]
  wire  tlb_OptimizationBarrier_16_io_x_pw; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178735.4]
  wire  tlb_OptimizationBarrier_16_io_x_px; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178735.4]
  wire  tlb_OptimizationBarrier_16_io_x_pr; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178735.4]
  wire  tlb_OptimizationBarrier_16_io_x_ppp; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178735.4]
  wire  tlb_OptimizationBarrier_16_io_x_pal; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178735.4]
  wire  tlb_OptimizationBarrier_16_io_x_paa; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178735.4]
  wire  tlb_OptimizationBarrier_16_io_x_eff; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178735.4]
  wire  tlb_OptimizationBarrier_16_io_x_c; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178735.4]
  wire [19:0] tlb_OptimizationBarrier_16_io_y_ppn; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178735.4]
  wire  tlb_OptimizationBarrier_16_io_y_u; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178735.4]
  wire  tlb_OptimizationBarrier_16_io_y_ae; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178735.4]
  wire  tlb_OptimizationBarrier_16_io_y_sw; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178735.4]
  wire  tlb_OptimizationBarrier_16_io_y_sx; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178735.4]
  wire  tlb_OptimizationBarrier_16_io_y_sr; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178735.4]
  wire  tlb_OptimizationBarrier_16_io_y_pw; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178735.4]
  wire  tlb_OptimizationBarrier_16_io_y_px; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178735.4]
  wire  tlb_OptimizationBarrier_16_io_y_pr; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178735.4]
  wire  tlb_OptimizationBarrier_16_io_y_ppp; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178735.4]
  wire  tlb_OptimizationBarrier_16_io_y_pal; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178735.4]
  wire  tlb_OptimizationBarrier_16_io_y_paa; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178735.4]
  wire  tlb_OptimizationBarrier_16_io_y_eff; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178735.4]
  wire  tlb_OptimizationBarrier_16_io_y_c; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178735.4]
  wire [19:0] tlb_OptimizationBarrier_17_io_x_ppn; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178778.4]
  wire  tlb_OptimizationBarrier_17_io_x_u; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178778.4]
  wire  tlb_OptimizationBarrier_17_io_x_ae; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178778.4]
  wire  tlb_OptimizationBarrier_17_io_x_sw; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178778.4]
  wire  tlb_OptimizationBarrier_17_io_x_sx; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178778.4]
  wire  tlb_OptimizationBarrier_17_io_x_sr; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178778.4]
  wire  tlb_OptimizationBarrier_17_io_x_pw; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178778.4]
  wire  tlb_OptimizationBarrier_17_io_x_px; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178778.4]
  wire  tlb_OptimizationBarrier_17_io_x_pr; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178778.4]
  wire  tlb_OptimizationBarrier_17_io_x_ppp; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178778.4]
  wire  tlb_OptimizationBarrier_17_io_x_pal; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178778.4]
  wire  tlb_OptimizationBarrier_17_io_x_paa; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178778.4]
  wire  tlb_OptimizationBarrier_17_io_x_eff; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178778.4]
  wire  tlb_OptimizationBarrier_17_io_x_c; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178778.4]
  wire [19:0] tlb_OptimizationBarrier_17_io_y_ppn; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178778.4]
  wire  tlb_OptimizationBarrier_17_io_y_u; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178778.4]
  wire  tlb_OptimizationBarrier_17_io_y_ae; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178778.4]
  wire  tlb_OptimizationBarrier_17_io_y_sw; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178778.4]
  wire  tlb_OptimizationBarrier_17_io_y_sx; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178778.4]
  wire  tlb_OptimizationBarrier_17_io_y_sr; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178778.4]
  wire  tlb_OptimizationBarrier_17_io_y_pw; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178778.4]
  wire  tlb_OptimizationBarrier_17_io_y_px; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178778.4]
  wire  tlb_OptimizationBarrier_17_io_y_pr; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178778.4]
  wire  tlb_OptimizationBarrier_17_io_y_ppp; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178778.4]
  wire  tlb_OptimizationBarrier_17_io_y_pal; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178778.4]
  wire  tlb_OptimizationBarrier_17_io_y_paa; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178778.4]
  wire  tlb_OptimizationBarrier_17_io_y_eff; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178778.4]
  wire  tlb_OptimizationBarrier_17_io_y_c; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178778.4]
  wire [19:0] tlb_OptimizationBarrier_18_io_x_ppn; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178821.4]
  wire  tlb_OptimizationBarrier_18_io_x_u; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178821.4]
  wire  tlb_OptimizationBarrier_18_io_x_ae; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178821.4]
  wire  tlb_OptimizationBarrier_18_io_x_sw; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178821.4]
  wire  tlb_OptimizationBarrier_18_io_x_sx; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178821.4]
  wire  tlb_OptimizationBarrier_18_io_x_sr; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178821.4]
  wire  tlb_OptimizationBarrier_18_io_x_pw; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178821.4]
  wire  tlb_OptimizationBarrier_18_io_x_px; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178821.4]
  wire  tlb_OptimizationBarrier_18_io_x_pr; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178821.4]
  wire  tlb_OptimizationBarrier_18_io_x_ppp; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178821.4]
  wire  tlb_OptimizationBarrier_18_io_x_pal; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178821.4]
  wire  tlb_OptimizationBarrier_18_io_x_paa; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178821.4]
  wire  tlb_OptimizationBarrier_18_io_x_eff; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178821.4]
  wire  tlb_OptimizationBarrier_18_io_x_c; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178821.4]
  wire [19:0] tlb_OptimizationBarrier_18_io_y_ppn; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178821.4]
  wire  tlb_OptimizationBarrier_18_io_y_u; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178821.4]
  wire  tlb_OptimizationBarrier_18_io_y_ae; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178821.4]
  wire  tlb_OptimizationBarrier_18_io_y_sw; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178821.4]
  wire  tlb_OptimizationBarrier_18_io_y_sx; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178821.4]
  wire  tlb_OptimizationBarrier_18_io_y_sr; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178821.4]
  wire  tlb_OptimizationBarrier_18_io_y_pw; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178821.4]
  wire  tlb_OptimizationBarrier_18_io_y_px; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178821.4]
  wire  tlb_OptimizationBarrier_18_io_y_pr; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178821.4]
  wire  tlb_OptimizationBarrier_18_io_y_ppp; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178821.4]
  wire  tlb_OptimizationBarrier_18_io_y_pal; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178821.4]
  wire  tlb_OptimizationBarrier_18_io_y_paa; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178821.4]
  wire  tlb_OptimizationBarrier_18_io_y_eff; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178821.4]
  wire  tlb_OptimizationBarrier_18_io_y_c; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178821.4]
  wire [19:0] tlb_OptimizationBarrier_19_io_x_ppn; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178864.4]
  wire  tlb_OptimizationBarrier_19_io_x_u; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178864.4]
  wire  tlb_OptimizationBarrier_19_io_x_ae; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178864.4]
  wire  tlb_OptimizationBarrier_19_io_x_sw; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178864.4]
  wire  tlb_OptimizationBarrier_19_io_x_sx; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178864.4]
  wire  tlb_OptimizationBarrier_19_io_x_sr; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178864.4]
  wire  tlb_OptimizationBarrier_19_io_x_pw; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178864.4]
  wire  tlb_OptimizationBarrier_19_io_x_px; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178864.4]
  wire  tlb_OptimizationBarrier_19_io_x_pr; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178864.4]
  wire  tlb_OptimizationBarrier_19_io_x_ppp; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178864.4]
  wire  tlb_OptimizationBarrier_19_io_x_pal; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178864.4]
  wire  tlb_OptimizationBarrier_19_io_x_paa; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178864.4]
  wire  tlb_OptimizationBarrier_19_io_x_eff; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178864.4]
  wire  tlb_OptimizationBarrier_19_io_x_c; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178864.4]
  wire [19:0] tlb_OptimizationBarrier_19_io_y_ppn; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178864.4]
  wire  tlb_OptimizationBarrier_19_io_y_u; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178864.4]
  wire  tlb_OptimizationBarrier_19_io_y_ae; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178864.4]
  wire  tlb_OptimizationBarrier_19_io_y_sw; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178864.4]
  wire  tlb_OptimizationBarrier_19_io_y_sx; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178864.4]
  wire  tlb_OptimizationBarrier_19_io_y_sr; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178864.4]
  wire  tlb_OptimizationBarrier_19_io_y_pw; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178864.4]
  wire  tlb_OptimizationBarrier_19_io_y_px; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178864.4]
  wire  tlb_OptimizationBarrier_19_io_y_pr; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178864.4]
  wire  tlb_OptimizationBarrier_19_io_y_ppp; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178864.4]
  wire  tlb_OptimizationBarrier_19_io_y_pal; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178864.4]
  wire  tlb_OptimizationBarrier_19_io_y_paa; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178864.4]
  wire  tlb_OptimizationBarrier_19_io_y_eff; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178864.4]
  wire  tlb_OptimizationBarrier_19_io_y_c; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178864.4]
  wire [19:0] tlb_OptimizationBarrier_20_io_x_ppn; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178907.4]
  wire  tlb_OptimizationBarrier_20_io_x_u; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178907.4]
  wire  tlb_OptimizationBarrier_20_io_x_ae; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178907.4]
  wire  tlb_OptimizationBarrier_20_io_x_sw; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178907.4]
  wire  tlb_OptimizationBarrier_20_io_x_sx; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178907.4]
  wire  tlb_OptimizationBarrier_20_io_x_sr; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178907.4]
  wire  tlb_OptimizationBarrier_20_io_x_pw; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178907.4]
  wire  tlb_OptimizationBarrier_20_io_x_px; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178907.4]
  wire  tlb_OptimizationBarrier_20_io_x_pr; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178907.4]
  wire  tlb_OptimizationBarrier_20_io_x_ppp; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178907.4]
  wire  tlb_OptimizationBarrier_20_io_x_pal; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178907.4]
  wire  tlb_OptimizationBarrier_20_io_x_paa; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178907.4]
  wire  tlb_OptimizationBarrier_20_io_x_eff; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178907.4]
  wire  tlb_OptimizationBarrier_20_io_x_c; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178907.4]
  wire [19:0] tlb_OptimizationBarrier_20_io_y_ppn; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178907.4]
  wire  tlb_OptimizationBarrier_20_io_y_u; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178907.4]
  wire  tlb_OptimizationBarrier_20_io_y_ae; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178907.4]
  wire  tlb_OptimizationBarrier_20_io_y_sw; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178907.4]
  wire  tlb_OptimizationBarrier_20_io_y_sx; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178907.4]
  wire  tlb_OptimizationBarrier_20_io_y_sr; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178907.4]
  wire  tlb_OptimizationBarrier_20_io_y_pw; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178907.4]
  wire  tlb_OptimizationBarrier_20_io_y_px; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178907.4]
  wire  tlb_OptimizationBarrier_20_io_y_pr; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178907.4]
  wire  tlb_OptimizationBarrier_20_io_y_ppp; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178907.4]
  wire  tlb_OptimizationBarrier_20_io_y_pal; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178907.4]
  wire  tlb_OptimizationBarrier_20_io_y_paa; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178907.4]
  wire  tlb_OptimizationBarrier_20_io_y_eff; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178907.4]
  wire  tlb_OptimizationBarrier_20_io_y_c; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178907.4]
  wire [19:0] tlb_OptimizationBarrier_21_io_x_ppn; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178950.4]
  wire  tlb_OptimizationBarrier_21_io_x_u; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178950.4]
  wire  tlb_OptimizationBarrier_21_io_x_ae; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178950.4]
  wire  tlb_OptimizationBarrier_21_io_x_sw; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178950.4]
  wire  tlb_OptimizationBarrier_21_io_x_sx; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178950.4]
  wire  tlb_OptimizationBarrier_21_io_x_sr; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178950.4]
  wire  tlb_OptimizationBarrier_21_io_x_pw; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178950.4]
  wire  tlb_OptimizationBarrier_21_io_x_px; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178950.4]
  wire  tlb_OptimizationBarrier_21_io_x_pr; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178950.4]
  wire  tlb_OptimizationBarrier_21_io_x_ppp; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178950.4]
  wire  tlb_OptimizationBarrier_21_io_x_pal; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178950.4]
  wire  tlb_OptimizationBarrier_21_io_x_paa; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178950.4]
  wire  tlb_OptimizationBarrier_21_io_x_eff; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178950.4]
  wire  tlb_OptimizationBarrier_21_io_x_c; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178950.4]
  wire [19:0] tlb_OptimizationBarrier_21_io_y_ppn; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178950.4]
  wire  tlb_OptimizationBarrier_21_io_y_u; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178950.4]
  wire  tlb_OptimizationBarrier_21_io_y_ae; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178950.4]
  wire  tlb_OptimizationBarrier_21_io_y_sw; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178950.4]
  wire  tlb_OptimizationBarrier_21_io_y_sx; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178950.4]
  wire  tlb_OptimizationBarrier_21_io_y_sr; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178950.4]
  wire  tlb_OptimizationBarrier_21_io_y_pw; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178950.4]
  wire  tlb_OptimizationBarrier_21_io_y_px; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178950.4]
  wire  tlb_OptimizationBarrier_21_io_y_pr; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178950.4]
  wire  tlb_OptimizationBarrier_21_io_y_ppp; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178950.4]
  wire  tlb_OptimizationBarrier_21_io_y_pal; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178950.4]
  wire  tlb_OptimizationBarrier_21_io_y_paa; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178950.4]
  wire  tlb_OptimizationBarrier_21_io_y_eff; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178950.4]
  wire  tlb_OptimizationBarrier_21_io_y_c; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178950.4]
  wire [19:0] tlb_OptimizationBarrier_22_io_x_ppn; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178992.4]
  wire  tlb_OptimizationBarrier_22_io_x_u; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178992.4]
  wire  tlb_OptimizationBarrier_22_io_x_ae; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178992.4]
  wire  tlb_OptimizationBarrier_22_io_x_sw; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178992.4]
  wire  tlb_OptimizationBarrier_22_io_x_sx; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178992.4]
  wire  tlb_OptimizationBarrier_22_io_x_sr; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178992.4]
  wire  tlb_OptimizationBarrier_22_io_x_pw; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178992.4]
  wire  tlb_OptimizationBarrier_22_io_x_px; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178992.4]
  wire  tlb_OptimizationBarrier_22_io_x_pr; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178992.4]
  wire  tlb_OptimizationBarrier_22_io_x_ppp; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178992.4]
  wire  tlb_OptimizationBarrier_22_io_x_pal; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178992.4]
  wire  tlb_OptimizationBarrier_22_io_x_paa; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178992.4]
  wire  tlb_OptimizationBarrier_22_io_x_eff; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178992.4]
  wire  tlb_OptimizationBarrier_22_io_x_c; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178992.4]
  wire [19:0] tlb_OptimizationBarrier_22_io_y_ppn; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178992.4]
  wire  tlb_OptimizationBarrier_22_io_y_u; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178992.4]
  wire  tlb_OptimizationBarrier_22_io_y_ae; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178992.4]
  wire  tlb_OptimizationBarrier_22_io_y_sw; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178992.4]
  wire  tlb_OptimizationBarrier_22_io_y_sx; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178992.4]
  wire  tlb_OptimizationBarrier_22_io_y_sr; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178992.4]
  wire  tlb_OptimizationBarrier_22_io_y_pw; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178992.4]
  wire  tlb_OptimizationBarrier_22_io_y_px; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178992.4]
  wire  tlb_OptimizationBarrier_22_io_y_pr; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178992.4]
  wire  tlb_OptimizationBarrier_22_io_y_ppp; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178992.4]
  wire  tlb_OptimizationBarrier_22_io_y_pal; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178992.4]
  wire  tlb_OptimizationBarrier_22_io_y_paa; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178992.4]
  wire  tlb_OptimizationBarrier_22_io_y_eff; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178992.4]
  wire  tlb_OptimizationBarrier_22_io_y_c; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178992.4]
  wire [19:0] tlb_OptimizationBarrier_23_io_x_ppn; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179034.4]
  wire  tlb_OptimizationBarrier_23_io_x_u; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179034.4]
  wire  tlb_OptimizationBarrier_23_io_x_ae; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179034.4]
  wire  tlb_OptimizationBarrier_23_io_x_sw; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179034.4]
  wire  tlb_OptimizationBarrier_23_io_x_sx; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179034.4]
  wire  tlb_OptimizationBarrier_23_io_x_sr; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179034.4]
  wire  tlb_OptimizationBarrier_23_io_x_pw; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179034.4]
  wire  tlb_OptimizationBarrier_23_io_x_px; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179034.4]
  wire  tlb_OptimizationBarrier_23_io_x_pr; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179034.4]
  wire  tlb_OptimizationBarrier_23_io_x_ppp; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179034.4]
  wire  tlb_OptimizationBarrier_23_io_x_pal; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179034.4]
  wire  tlb_OptimizationBarrier_23_io_x_paa; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179034.4]
  wire  tlb_OptimizationBarrier_23_io_x_eff; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179034.4]
  wire  tlb_OptimizationBarrier_23_io_x_c; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179034.4]
  wire [19:0] tlb_OptimizationBarrier_23_io_y_ppn; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179034.4]
  wire  tlb_OptimizationBarrier_23_io_y_u; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179034.4]
  wire  tlb_OptimizationBarrier_23_io_y_ae; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179034.4]
  wire  tlb_OptimizationBarrier_23_io_y_sw; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179034.4]
  wire  tlb_OptimizationBarrier_23_io_y_sx; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179034.4]
  wire  tlb_OptimizationBarrier_23_io_y_sr; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179034.4]
  wire  tlb_OptimizationBarrier_23_io_y_pw; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179034.4]
  wire  tlb_OptimizationBarrier_23_io_y_px; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179034.4]
  wire  tlb_OptimizationBarrier_23_io_y_pr; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179034.4]
  wire  tlb_OptimizationBarrier_23_io_y_ppp; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179034.4]
  wire  tlb_OptimizationBarrier_23_io_y_pal; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179034.4]
  wire  tlb_OptimizationBarrier_23_io_y_paa; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179034.4]
  wire  tlb_OptimizationBarrier_23_io_y_eff; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179034.4]
  wire  tlb_OptimizationBarrier_23_io_y_c; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179034.4]
  wire [19:0] tlb_OptimizationBarrier_24_io_x_ppn; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179076.4]
  wire  tlb_OptimizationBarrier_24_io_x_u; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179076.4]
  wire  tlb_OptimizationBarrier_24_io_x_ae; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179076.4]
  wire  tlb_OptimizationBarrier_24_io_x_sw; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179076.4]
  wire  tlb_OptimizationBarrier_24_io_x_sx; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179076.4]
  wire  tlb_OptimizationBarrier_24_io_x_sr; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179076.4]
  wire  tlb_OptimizationBarrier_24_io_x_pw; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179076.4]
  wire  tlb_OptimizationBarrier_24_io_x_px; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179076.4]
  wire  tlb_OptimizationBarrier_24_io_x_pr; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179076.4]
  wire  tlb_OptimizationBarrier_24_io_x_ppp; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179076.4]
  wire  tlb_OptimizationBarrier_24_io_x_pal; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179076.4]
  wire  tlb_OptimizationBarrier_24_io_x_paa; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179076.4]
  wire  tlb_OptimizationBarrier_24_io_x_eff; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179076.4]
  wire  tlb_OptimizationBarrier_24_io_x_c; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179076.4]
  wire [19:0] tlb_OptimizationBarrier_24_io_y_ppn; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179076.4]
  wire  tlb_OptimizationBarrier_24_io_y_u; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179076.4]
  wire  tlb_OptimizationBarrier_24_io_y_ae; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179076.4]
  wire  tlb_OptimizationBarrier_24_io_y_sw; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179076.4]
  wire  tlb_OptimizationBarrier_24_io_y_sx; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179076.4]
  wire  tlb_OptimizationBarrier_24_io_y_sr; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179076.4]
  wire  tlb_OptimizationBarrier_24_io_y_pw; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179076.4]
  wire  tlb_OptimizationBarrier_24_io_y_px; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179076.4]
  wire  tlb_OptimizationBarrier_24_io_y_pr; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179076.4]
  wire  tlb_OptimizationBarrier_24_io_y_ppp; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179076.4]
  wire  tlb_OptimizationBarrier_24_io_y_pal; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179076.4]
  wire  tlb_OptimizationBarrier_24_io_y_paa; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179076.4]
  wire  tlb_OptimizationBarrier_24_io_y_eff; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179076.4]
  wire  tlb_OptimizationBarrier_24_io_y_c; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179076.4]
  wire [19:0] tlb_OptimizationBarrier_25_io_x_ppn; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179118.4]
  wire  tlb_OptimizationBarrier_25_io_x_u; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179118.4]
  wire  tlb_OptimizationBarrier_25_io_x_ae; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179118.4]
  wire  tlb_OptimizationBarrier_25_io_x_sw; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179118.4]
  wire  tlb_OptimizationBarrier_25_io_x_sx; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179118.4]
  wire  tlb_OptimizationBarrier_25_io_x_sr; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179118.4]
  wire  tlb_OptimizationBarrier_25_io_x_pw; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179118.4]
  wire  tlb_OptimizationBarrier_25_io_x_px; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179118.4]
  wire  tlb_OptimizationBarrier_25_io_x_pr; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179118.4]
  wire  tlb_OptimizationBarrier_25_io_x_ppp; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179118.4]
  wire  tlb_OptimizationBarrier_25_io_x_pal; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179118.4]
  wire  tlb_OptimizationBarrier_25_io_x_paa; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179118.4]
  wire  tlb_OptimizationBarrier_25_io_x_eff; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179118.4]
  wire  tlb_OptimizationBarrier_25_io_x_c; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179118.4]
  wire [19:0] tlb_OptimizationBarrier_25_io_y_ppn; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179118.4]
  wire  tlb_OptimizationBarrier_25_io_y_u; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179118.4]
  wire  tlb_OptimizationBarrier_25_io_y_ae; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179118.4]
  wire  tlb_OptimizationBarrier_25_io_y_sw; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179118.4]
  wire  tlb_OptimizationBarrier_25_io_y_sx; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179118.4]
  wire  tlb_OptimizationBarrier_25_io_y_sr; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179118.4]
  wire  tlb_OptimizationBarrier_25_io_y_pw; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179118.4]
  wire  tlb_OptimizationBarrier_25_io_y_px; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179118.4]
  wire  tlb_OptimizationBarrier_25_io_y_pr; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179118.4]
  wire  tlb_OptimizationBarrier_25_io_y_ppp; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179118.4]
  wire  tlb_OptimizationBarrier_25_io_y_pal; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179118.4]
  wire  tlb_OptimizationBarrier_25_io_y_paa; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179118.4]
  wire  tlb_OptimizationBarrier_25_io_y_eff; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179118.4]
  wire  tlb_OptimizationBarrier_25_io_y_c; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179118.4]
  wire [19:0] tlb_OptimizationBarrier_26_io_x_ppn; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179160.4]
  wire  tlb_OptimizationBarrier_26_io_x_u; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179160.4]
  wire  tlb_OptimizationBarrier_26_io_x_ae; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179160.4]
  wire  tlb_OptimizationBarrier_26_io_x_sw; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179160.4]
  wire  tlb_OptimizationBarrier_26_io_x_sx; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179160.4]
  wire  tlb_OptimizationBarrier_26_io_x_sr; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179160.4]
  wire  tlb_OptimizationBarrier_26_io_x_pw; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179160.4]
  wire  tlb_OptimizationBarrier_26_io_x_px; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179160.4]
  wire  tlb_OptimizationBarrier_26_io_x_pr; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179160.4]
  wire  tlb_OptimizationBarrier_26_io_x_ppp; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179160.4]
  wire  tlb_OptimizationBarrier_26_io_x_pal; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179160.4]
  wire  tlb_OptimizationBarrier_26_io_x_paa; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179160.4]
  wire  tlb_OptimizationBarrier_26_io_x_eff; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179160.4]
  wire  tlb_OptimizationBarrier_26_io_x_c; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179160.4]
  wire [19:0] tlb_OptimizationBarrier_26_io_y_ppn; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179160.4]
  wire  tlb_OptimizationBarrier_26_io_y_u; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179160.4]
  wire  tlb_OptimizationBarrier_26_io_y_ae; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179160.4]
  wire  tlb_OptimizationBarrier_26_io_y_sw; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179160.4]
  wire  tlb_OptimizationBarrier_26_io_y_sx; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179160.4]
  wire  tlb_OptimizationBarrier_26_io_y_sr; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179160.4]
  wire  tlb_OptimizationBarrier_26_io_y_pw; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179160.4]
  wire  tlb_OptimizationBarrier_26_io_y_px; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179160.4]
  wire  tlb_OptimizationBarrier_26_io_y_pr; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179160.4]
  wire  tlb_OptimizationBarrier_26_io_y_ppp; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179160.4]
  wire  tlb_OptimizationBarrier_26_io_y_pal; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179160.4]
  wire  tlb_OptimizationBarrier_26_io_y_paa; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179160.4]
  wire  tlb_OptimizationBarrier_26_io_y_eff; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179160.4]
  wire  tlb_OptimizationBarrier_26_io_y_c; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179160.4]
  wire [19:0] tlb_OptimizationBarrier_27_io_x_ppn; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179203.4]
  wire  tlb_OptimizationBarrier_27_io_x_u; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179203.4]
  wire  tlb_OptimizationBarrier_27_io_x_ae; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179203.4]
  wire  tlb_OptimizationBarrier_27_io_x_sw; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179203.4]
  wire  tlb_OptimizationBarrier_27_io_x_sx; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179203.4]
  wire  tlb_OptimizationBarrier_27_io_x_sr; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179203.4]
  wire  tlb_OptimizationBarrier_27_io_x_pw; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179203.4]
  wire  tlb_OptimizationBarrier_27_io_x_px; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179203.4]
  wire  tlb_OptimizationBarrier_27_io_x_pr; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179203.4]
  wire  tlb_OptimizationBarrier_27_io_x_ppp; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179203.4]
  wire  tlb_OptimizationBarrier_27_io_x_pal; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179203.4]
  wire  tlb_OptimizationBarrier_27_io_x_paa; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179203.4]
  wire  tlb_OptimizationBarrier_27_io_x_eff; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179203.4]
  wire  tlb_OptimizationBarrier_27_io_x_c; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179203.4]
  wire [19:0] tlb_OptimizationBarrier_27_io_y_ppn; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179203.4]
  wire  tlb_OptimizationBarrier_27_io_y_u; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179203.4]
  wire  tlb_OptimizationBarrier_27_io_y_ae; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179203.4]
  wire  tlb_OptimizationBarrier_27_io_y_sw; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179203.4]
  wire  tlb_OptimizationBarrier_27_io_y_sx; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179203.4]
  wire  tlb_OptimizationBarrier_27_io_y_sr; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179203.4]
  wire  tlb_OptimizationBarrier_27_io_y_pw; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179203.4]
  wire  tlb_OptimizationBarrier_27_io_y_px; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179203.4]
  wire  tlb_OptimizationBarrier_27_io_y_pr; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179203.4]
  wire  tlb_OptimizationBarrier_27_io_y_ppp; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179203.4]
  wire  tlb_OptimizationBarrier_27_io_y_pal; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179203.4]
  wire  tlb_OptimizationBarrier_27_io_y_paa; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179203.4]
  wire  tlb_OptimizationBarrier_27_io_y_eff; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179203.4]
  wire  tlb_OptimizationBarrier_27_io_y_c; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179203.4]
  wire [19:0] tlb_OptimizationBarrier_28_io_x_ppn; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179246.4]
  wire  tlb_OptimizationBarrier_28_io_x_u; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179246.4]
  wire  tlb_OptimizationBarrier_28_io_x_ae; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179246.4]
  wire  tlb_OptimizationBarrier_28_io_x_sw; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179246.4]
  wire  tlb_OptimizationBarrier_28_io_x_sx; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179246.4]
  wire  tlb_OptimizationBarrier_28_io_x_sr; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179246.4]
  wire  tlb_OptimizationBarrier_28_io_x_pw; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179246.4]
  wire  tlb_OptimizationBarrier_28_io_x_px; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179246.4]
  wire  tlb_OptimizationBarrier_28_io_x_pr; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179246.4]
  wire  tlb_OptimizationBarrier_28_io_x_ppp; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179246.4]
  wire  tlb_OptimizationBarrier_28_io_x_pal; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179246.4]
  wire  tlb_OptimizationBarrier_28_io_x_paa; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179246.4]
  wire  tlb_OptimizationBarrier_28_io_x_eff; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179246.4]
  wire  tlb_OptimizationBarrier_28_io_x_c; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179246.4]
  wire [19:0] tlb_OptimizationBarrier_28_io_y_ppn; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179246.4]
  wire  tlb_OptimizationBarrier_28_io_y_u; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179246.4]
  wire  tlb_OptimizationBarrier_28_io_y_ae; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179246.4]
  wire  tlb_OptimizationBarrier_28_io_y_sw; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179246.4]
  wire  tlb_OptimizationBarrier_28_io_y_sx; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179246.4]
  wire  tlb_OptimizationBarrier_28_io_y_sr; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179246.4]
  wire  tlb_OptimizationBarrier_28_io_y_pw; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179246.4]
  wire  tlb_OptimizationBarrier_28_io_y_px; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179246.4]
  wire  tlb_OptimizationBarrier_28_io_y_pr; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179246.4]
  wire  tlb_OptimizationBarrier_28_io_y_ppp; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179246.4]
  wire  tlb_OptimizationBarrier_28_io_y_pal; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179246.4]
  wire  tlb_OptimizationBarrier_28_io_y_paa; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179246.4]
  wire  tlb_OptimizationBarrier_28_io_y_eff; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179246.4]
  wire  tlb_OptimizationBarrier_28_io_y_c; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179246.4]
  wire [19:0] tlb_OptimizationBarrier_29_io_x_ppn; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179289.4]
  wire  tlb_OptimizationBarrier_29_io_x_u; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179289.4]
  wire  tlb_OptimizationBarrier_29_io_x_ae; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179289.4]
  wire  tlb_OptimizationBarrier_29_io_x_sw; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179289.4]
  wire  tlb_OptimizationBarrier_29_io_x_sx; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179289.4]
  wire  tlb_OptimizationBarrier_29_io_x_sr; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179289.4]
  wire  tlb_OptimizationBarrier_29_io_x_pw; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179289.4]
  wire  tlb_OptimizationBarrier_29_io_x_px; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179289.4]
  wire  tlb_OptimizationBarrier_29_io_x_pr; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179289.4]
  wire  tlb_OptimizationBarrier_29_io_x_ppp; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179289.4]
  wire  tlb_OptimizationBarrier_29_io_x_pal; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179289.4]
  wire  tlb_OptimizationBarrier_29_io_x_paa; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179289.4]
  wire  tlb_OptimizationBarrier_29_io_x_eff; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179289.4]
  wire  tlb_OptimizationBarrier_29_io_x_c; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179289.4]
  wire [19:0] tlb_OptimizationBarrier_29_io_y_ppn; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179289.4]
  wire  tlb_OptimizationBarrier_29_io_y_u; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179289.4]
  wire  tlb_OptimizationBarrier_29_io_y_ae; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179289.4]
  wire  tlb_OptimizationBarrier_29_io_y_sw; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179289.4]
  wire  tlb_OptimizationBarrier_29_io_y_sx; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179289.4]
  wire  tlb_OptimizationBarrier_29_io_y_sr; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179289.4]
  wire  tlb_OptimizationBarrier_29_io_y_pw; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179289.4]
  wire  tlb_OptimizationBarrier_29_io_y_px; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179289.4]
  wire  tlb_OptimizationBarrier_29_io_y_pr; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179289.4]
  wire  tlb_OptimizationBarrier_29_io_y_ppp; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179289.4]
  wire  tlb_OptimizationBarrier_29_io_y_pal; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179289.4]
  wire  tlb_OptimizationBarrier_29_io_y_paa; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179289.4]
  wire  tlb_OptimizationBarrier_29_io_y_eff; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179289.4]
  wire  tlb_OptimizationBarrier_29_io_y_c; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179289.4]
  wire [19:0] tlb_OptimizationBarrier_30_io_x_ppn; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179332.4]
  wire  tlb_OptimizationBarrier_30_io_x_u; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179332.4]
  wire  tlb_OptimizationBarrier_30_io_x_ae; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179332.4]
  wire  tlb_OptimizationBarrier_30_io_x_sw; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179332.4]
  wire  tlb_OptimizationBarrier_30_io_x_sx; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179332.4]
  wire  tlb_OptimizationBarrier_30_io_x_sr; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179332.4]
  wire  tlb_OptimizationBarrier_30_io_x_pw; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179332.4]
  wire  tlb_OptimizationBarrier_30_io_x_px; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179332.4]
  wire  tlb_OptimizationBarrier_30_io_x_pr; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179332.4]
  wire  tlb_OptimizationBarrier_30_io_x_ppp; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179332.4]
  wire  tlb_OptimizationBarrier_30_io_x_pal; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179332.4]
  wire  tlb_OptimizationBarrier_30_io_x_paa; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179332.4]
  wire  tlb_OptimizationBarrier_30_io_x_eff; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179332.4]
  wire  tlb_OptimizationBarrier_30_io_x_c; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179332.4]
  wire [19:0] tlb_OptimizationBarrier_30_io_y_ppn; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179332.4]
  wire  tlb_OptimizationBarrier_30_io_y_u; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179332.4]
  wire  tlb_OptimizationBarrier_30_io_y_ae; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179332.4]
  wire  tlb_OptimizationBarrier_30_io_y_sw; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179332.4]
  wire  tlb_OptimizationBarrier_30_io_y_sx; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179332.4]
  wire  tlb_OptimizationBarrier_30_io_y_sr; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179332.4]
  wire  tlb_OptimizationBarrier_30_io_y_pw; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179332.4]
  wire  tlb_OptimizationBarrier_30_io_y_px; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179332.4]
  wire  tlb_OptimizationBarrier_30_io_y_pr; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179332.4]
  wire  tlb_OptimizationBarrier_30_io_y_ppp; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179332.4]
  wire  tlb_OptimizationBarrier_30_io_y_pal; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179332.4]
  wire  tlb_OptimizationBarrier_30_io_y_paa; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179332.4]
  wire  tlb_OptimizationBarrier_30_io_y_eff; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179332.4]
  wire  tlb_OptimizationBarrier_30_io_y_c; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179332.4]
  wire [19:0] tlb_OptimizationBarrier_31_io_x_ppn; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179375.4]
  wire  tlb_OptimizationBarrier_31_io_x_u; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179375.4]
  wire  tlb_OptimizationBarrier_31_io_x_ae; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179375.4]
  wire  tlb_OptimizationBarrier_31_io_x_sw; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179375.4]
  wire  tlb_OptimizationBarrier_31_io_x_sx; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179375.4]
  wire  tlb_OptimizationBarrier_31_io_x_sr; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179375.4]
  wire  tlb_OptimizationBarrier_31_io_x_pw; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179375.4]
  wire  tlb_OptimizationBarrier_31_io_x_px; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179375.4]
  wire  tlb_OptimizationBarrier_31_io_x_pr; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179375.4]
  wire  tlb_OptimizationBarrier_31_io_x_ppp; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179375.4]
  wire  tlb_OptimizationBarrier_31_io_x_pal; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179375.4]
  wire  tlb_OptimizationBarrier_31_io_x_paa; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179375.4]
  wire  tlb_OptimizationBarrier_31_io_x_eff; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179375.4]
  wire  tlb_OptimizationBarrier_31_io_x_c; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179375.4]
  wire [19:0] tlb_OptimizationBarrier_31_io_y_ppn; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179375.4]
  wire  tlb_OptimizationBarrier_31_io_y_u; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179375.4]
  wire  tlb_OptimizationBarrier_31_io_y_ae; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179375.4]
  wire  tlb_OptimizationBarrier_31_io_y_sw; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179375.4]
  wire  tlb_OptimizationBarrier_31_io_y_sx; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179375.4]
  wire  tlb_OptimizationBarrier_31_io_y_sr; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179375.4]
  wire  tlb_OptimizationBarrier_31_io_y_pw; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179375.4]
  wire  tlb_OptimizationBarrier_31_io_y_px; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179375.4]
  wire  tlb_OptimizationBarrier_31_io_y_pr; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179375.4]
  wire  tlb_OptimizationBarrier_31_io_y_ppp; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179375.4]
  wire  tlb_OptimizationBarrier_31_io_y_pal; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179375.4]
  wire  tlb_OptimizationBarrier_31_io_y_paa; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179375.4]
  wire  tlb_OptimizationBarrier_31_io_y_eff; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179375.4]
  wire  tlb_OptimizationBarrier_31_io_y_c; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179375.4]
  wire [19:0] tlb_OptimizationBarrier_32_io_x_ppn; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179418.4]
  wire  tlb_OptimizationBarrier_32_io_x_u; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179418.4]
  wire  tlb_OptimizationBarrier_32_io_x_ae; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179418.4]
  wire  tlb_OptimizationBarrier_32_io_x_sw; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179418.4]
  wire  tlb_OptimizationBarrier_32_io_x_sx; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179418.4]
  wire  tlb_OptimizationBarrier_32_io_x_sr; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179418.4]
  wire  tlb_OptimizationBarrier_32_io_x_pw; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179418.4]
  wire  tlb_OptimizationBarrier_32_io_x_px; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179418.4]
  wire  tlb_OptimizationBarrier_32_io_x_pr; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179418.4]
  wire  tlb_OptimizationBarrier_32_io_x_ppp; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179418.4]
  wire  tlb_OptimizationBarrier_32_io_x_pal; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179418.4]
  wire  tlb_OptimizationBarrier_32_io_x_paa; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179418.4]
  wire  tlb_OptimizationBarrier_32_io_x_eff; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179418.4]
  wire  tlb_OptimizationBarrier_32_io_x_c; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179418.4]
  wire [19:0] tlb_OptimizationBarrier_32_io_y_ppn; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179418.4]
  wire  tlb_OptimizationBarrier_32_io_y_u; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179418.4]
  wire  tlb_OptimizationBarrier_32_io_y_ae; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179418.4]
  wire  tlb_OptimizationBarrier_32_io_y_sw; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179418.4]
  wire  tlb_OptimizationBarrier_32_io_y_sx; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179418.4]
  wire  tlb_OptimizationBarrier_32_io_y_sr; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179418.4]
  wire  tlb_OptimizationBarrier_32_io_y_pw; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179418.4]
  wire  tlb_OptimizationBarrier_32_io_y_px; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179418.4]
  wire  tlb_OptimizationBarrier_32_io_y_pr; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179418.4]
  wire  tlb_OptimizationBarrier_32_io_y_ppp; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179418.4]
  wire  tlb_OptimizationBarrier_32_io_y_pal; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179418.4]
  wire  tlb_OptimizationBarrier_32_io_y_paa; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179418.4]
  wire  tlb_OptimizationBarrier_32_io_y_eff; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179418.4]
  wire  tlb_OptimizationBarrier_32_io_y_c; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179418.4]
  wire [19:0] tlb_OptimizationBarrier_33_io_x_ppn; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179461.4]
  wire  tlb_OptimizationBarrier_33_io_x_u; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179461.4]
  wire  tlb_OptimizationBarrier_33_io_x_ae; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179461.4]
  wire  tlb_OptimizationBarrier_33_io_x_sw; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179461.4]
  wire  tlb_OptimizationBarrier_33_io_x_sx; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179461.4]
  wire  tlb_OptimizationBarrier_33_io_x_sr; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179461.4]
  wire  tlb_OptimizationBarrier_33_io_x_pw; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179461.4]
  wire  tlb_OptimizationBarrier_33_io_x_px; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179461.4]
  wire  tlb_OptimizationBarrier_33_io_x_pr; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179461.4]
  wire  tlb_OptimizationBarrier_33_io_x_ppp; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179461.4]
  wire  tlb_OptimizationBarrier_33_io_x_pal; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179461.4]
  wire  tlb_OptimizationBarrier_33_io_x_paa; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179461.4]
  wire  tlb_OptimizationBarrier_33_io_x_eff; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179461.4]
  wire  tlb_OptimizationBarrier_33_io_x_c; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179461.4]
  wire [19:0] tlb_OptimizationBarrier_33_io_y_ppn; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179461.4]
  wire  tlb_OptimizationBarrier_33_io_y_u; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179461.4]
  wire  tlb_OptimizationBarrier_33_io_y_ae; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179461.4]
  wire  tlb_OptimizationBarrier_33_io_y_sw; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179461.4]
  wire  tlb_OptimizationBarrier_33_io_y_sx; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179461.4]
  wire  tlb_OptimizationBarrier_33_io_y_sr; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179461.4]
  wire  tlb_OptimizationBarrier_33_io_y_pw; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179461.4]
  wire  tlb_OptimizationBarrier_33_io_y_px; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179461.4]
  wire  tlb_OptimizationBarrier_33_io_y_pr; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179461.4]
  wire  tlb_OptimizationBarrier_33_io_y_ppp; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179461.4]
  wire  tlb_OptimizationBarrier_33_io_y_pal; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179461.4]
  wire  tlb_OptimizationBarrier_33_io_y_paa; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179461.4]
  wire  tlb_OptimizationBarrier_33_io_y_eff; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179461.4]
  wire  tlb_OptimizationBarrier_33_io_y_c; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179461.4]
  wire [19:0] tlb_OptimizationBarrier_34_io_x_ppn; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179504.4]
  wire  tlb_OptimizationBarrier_34_io_x_u; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179504.4]
  wire  tlb_OptimizationBarrier_34_io_x_ae; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179504.4]
  wire  tlb_OptimizationBarrier_34_io_x_sw; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179504.4]
  wire  tlb_OptimizationBarrier_34_io_x_sx; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179504.4]
  wire  tlb_OptimizationBarrier_34_io_x_sr; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179504.4]
  wire  tlb_OptimizationBarrier_34_io_x_pw; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179504.4]
  wire  tlb_OptimizationBarrier_34_io_x_px; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179504.4]
  wire  tlb_OptimizationBarrier_34_io_x_pr; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179504.4]
  wire  tlb_OptimizationBarrier_34_io_x_ppp; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179504.4]
  wire  tlb_OptimizationBarrier_34_io_x_pal; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179504.4]
  wire  tlb_OptimizationBarrier_34_io_x_paa; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179504.4]
  wire  tlb_OptimizationBarrier_34_io_x_eff; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179504.4]
  wire  tlb_OptimizationBarrier_34_io_x_c; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179504.4]
  wire [19:0] tlb_OptimizationBarrier_34_io_y_ppn; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179504.4]
  wire  tlb_OptimizationBarrier_34_io_y_u; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179504.4]
  wire  tlb_OptimizationBarrier_34_io_y_ae; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179504.4]
  wire  tlb_OptimizationBarrier_34_io_y_sw; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179504.4]
  wire  tlb_OptimizationBarrier_34_io_y_sx; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179504.4]
  wire  tlb_OptimizationBarrier_34_io_y_sr; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179504.4]
  wire  tlb_OptimizationBarrier_34_io_y_pw; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179504.4]
  wire  tlb_OptimizationBarrier_34_io_y_px; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179504.4]
  wire  tlb_OptimizationBarrier_34_io_y_pr; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179504.4]
  wire  tlb_OptimizationBarrier_34_io_y_ppp; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179504.4]
  wire  tlb_OptimizationBarrier_34_io_y_pal; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179504.4]
  wire  tlb_OptimizationBarrier_34_io_y_paa; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179504.4]
  wire  tlb_OptimizationBarrier_34_io_y_eff; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179504.4]
  wire  tlb_OptimizationBarrier_34_io_y_c; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179504.4]
  wire [19:0] tlb_OptimizationBarrier_35_io_x_ppn; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179546.4]
  wire  tlb_OptimizationBarrier_35_io_x_u; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179546.4]
  wire  tlb_OptimizationBarrier_35_io_x_ae; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179546.4]
  wire  tlb_OptimizationBarrier_35_io_x_sw; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179546.4]
  wire  tlb_OptimizationBarrier_35_io_x_sx; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179546.4]
  wire  tlb_OptimizationBarrier_35_io_x_sr; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179546.4]
  wire  tlb_OptimizationBarrier_35_io_x_pw; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179546.4]
  wire  tlb_OptimizationBarrier_35_io_x_px; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179546.4]
  wire  tlb_OptimizationBarrier_35_io_x_pr; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179546.4]
  wire  tlb_OptimizationBarrier_35_io_x_ppp; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179546.4]
  wire  tlb_OptimizationBarrier_35_io_x_pal; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179546.4]
  wire  tlb_OptimizationBarrier_35_io_x_paa; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179546.4]
  wire  tlb_OptimizationBarrier_35_io_x_eff; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179546.4]
  wire  tlb_OptimizationBarrier_35_io_x_c; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179546.4]
  wire [19:0] tlb_OptimizationBarrier_35_io_y_ppn; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179546.4]
  wire  tlb_OptimizationBarrier_35_io_y_u; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179546.4]
  wire  tlb_OptimizationBarrier_35_io_y_ae; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179546.4]
  wire  tlb_OptimizationBarrier_35_io_y_sw; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179546.4]
  wire  tlb_OptimizationBarrier_35_io_y_sx; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179546.4]
  wire  tlb_OptimizationBarrier_35_io_y_sr; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179546.4]
  wire  tlb_OptimizationBarrier_35_io_y_pw; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179546.4]
  wire  tlb_OptimizationBarrier_35_io_y_px; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179546.4]
  wire  tlb_OptimizationBarrier_35_io_y_pr; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179546.4]
  wire  tlb_OptimizationBarrier_35_io_y_ppp; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179546.4]
  wire  tlb_OptimizationBarrier_35_io_y_pal; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179546.4]
  wire  tlb_OptimizationBarrier_35_io_y_paa; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179546.4]
  wire  tlb_OptimizationBarrier_35_io_y_eff; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179546.4]
  wire  tlb_OptimizationBarrier_35_io_y_c; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179546.4]
  wire [19:0] tlb_OptimizationBarrier_36_io_x_ppn; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179588.4]
  wire  tlb_OptimizationBarrier_36_io_x_u; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179588.4]
  wire  tlb_OptimizationBarrier_36_io_x_ae; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179588.4]
  wire  tlb_OptimizationBarrier_36_io_x_sw; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179588.4]
  wire  tlb_OptimizationBarrier_36_io_x_sx; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179588.4]
  wire  tlb_OptimizationBarrier_36_io_x_sr; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179588.4]
  wire  tlb_OptimizationBarrier_36_io_x_pw; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179588.4]
  wire  tlb_OptimizationBarrier_36_io_x_px; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179588.4]
  wire  tlb_OptimizationBarrier_36_io_x_pr; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179588.4]
  wire  tlb_OptimizationBarrier_36_io_x_ppp; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179588.4]
  wire  tlb_OptimizationBarrier_36_io_x_pal; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179588.4]
  wire  tlb_OptimizationBarrier_36_io_x_paa; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179588.4]
  wire  tlb_OptimizationBarrier_36_io_x_eff; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179588.4]
  wire  tlb_OptimizationBarrier_36_io_x_c; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179588.4]
  wire [19:0] tlb_OptimizationBarrier_36_io_y_ppn; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179588.4]
  wire  tlb_OptimizationBarrier_36_io_y_u; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179588.4]
  wire  tlb_OptimizationBarrier_36_io_y_ae; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179588.4]
  wire  tlb_OptimizationBarrier_36_io_y_sw; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179588.4]
  wire  tlb_OptimizationBarrier_36_io_y_sx; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179588.4]
  wire  tlb_OptimizationBarrier_36_io_y_sr; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179588.4]
  wire  tlb_OptimizationBarrier_36_io_y_pw; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179588.4]
  wire  tlb_OptimizationBarrier_36_io_y_px; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179588.4]
  wire  tlb_OptimizationBarrier_36_io_y_pr; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179588.4]
  wire  tlb_OptimizationBarrier_36_io_y_ppp; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179588.4]
  wire  tlb_OptimizationBarrier_36_io_y_pal; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179588.4]
  wire  tlb_OptimizationBarrier_36_io_y_paa; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179588.4]
  wire  tlb_OptimizationBarrier_36_io_y_eff; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179588.4]
  wire  tlb_OptimizationBarrier_36_io_y_c; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179588.4]
  wire [19:0] tlb_OptimizationBarrier_37_io_x_ppn; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179630.4]
  wire  tlb_OptimizationBarrier_37_io_x_u; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179630.4]
  wire  tlb_OptimizationBarrier_37_io_x_ae; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179630.4]
  wire  tlb_OptimizationBarrier_37_io_x_sw; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179630.4]
  wire  tlb_OptimizationBarrier_37_io_x_sx; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179630.4]
  wire  tlb_OptimizationBarrier_37_io_x_sr; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179630.4]
  wire  tlb_OptimizationBarrier_37_io_x_pw; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179630.4]
  wire  tlb_OptimizationBarrier_37_io_x_px; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179630.4]
  wire  tlb_OptimizationBarrier_37_io_x_pr; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179630.4]
  wire  tlb_OptimizationBarrier_37_io_x_ppp; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179630.4]
  wire  tlb_OptimizationBarrier_37_io_x_pal; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179630.4]
  wire  tlb_OptimizationBarrier_37_io_x_paa; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179630.4]
  wire  tlb_OptimizationBarrier_37_io_x_eff; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179630.4]
  wire  tlb_OptimizationBarrier_37_io_x_c; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179630.4]
  wire [19:0] tlb_OptimizationBarrier_37_io_y_ppn; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179630.4]
  wire  tlb_OptimizationBarrier_37_io_y_u; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179630.4]
  wire  tlb_OptimizationBarrier_37_io_y_ae; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179630.4]
  wire  tlb_OptimizationBarrier_37_io_y_sw; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179630.4]
  wire  tlb_OptimizationBarrier_37_io_y_sx; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179630.4]
  wire  tlb_OptimizationBarrier_37_io_y_sr; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179630.4]
  wire  tlb_OptimizationBarrier_37_io_y_pw; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179630.4]
  wire  tlb_OptimizationBarrier_37_io_y_px; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179630.4]
  wire  tlb_OptimizationBarrier_37_io_y_pr; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179630.4]
  wire  tlb_OptimizationBarrier_37_io_y_ppp; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179630.4]
  wire  tlb_OptimizationBarrier_37_io_y_pal; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179630.4]
  wire  tlb_OptimizationBarrier_37_io_y_paa; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179630.4]
  wire  tlb_OptimizationBarrier_37_io_y_eff; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179630.4]
  wire  tlb_OptimizationBarrier_37_io_y_c; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179630.4]
  wire [19:0] tlb_OptimizationBarrier_38_io_x_ppn; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179672.4]
  wire  tlb_OptimizationBarrier_38_io_x_u; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179672.4]
  wire  tlb_OptimizationBarrier_38_io_x_ae; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179672.4]
  wire  tlb_OptimizationBarrier_38_io_x_sw; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179672.4]
  wire  tlb_OptimizationBarrier_38_io_x_sx; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179672.4]
  wire  tlb_OptimizationBarrier_38_io_x_sr; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179672.4]
  wire  tlb_OptimizationBarrier_38_io_x_pw; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179672.4]
  wire  tlb_OptimizationBarrier_38_io_x_px; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179672.4]
  wire  tlb_OptimizationBarrier_38_io_x_pr; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179672.4]
  wire  tlb_OptimizationBarrier_38_io_x_ppp; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179672.4]
  wire  tlb_OptimizationBarrier_38_io_x_pal; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179672.4]
  wire  tlb_OptimizationBarrier_38_io_x_paa; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179672.4]
  wire  tlb_OptimizationBarrier_38_io_x_eff; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179672.4]
  wire  tlb_OptimizationBarrier_38_io_x_c; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179672.4]
  wire [19:0] tlb_OptimizationBarrier_38_io_y_ppn; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179672.4]
  wire  tlb_OptimizationBarrier_38_io_y_u; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179672.4]
  wire  tlb_OptimizationBarrier_38_io_y_ae; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179672.4]
  wire  tlb_OptimizationBarrier_38_io_y_sw; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179672.4]
  wire  tlb_OptimizationBarrier_38_io_y_sx; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179672.4]
  wire  tlb_OptimizationBarrier_38_io_y_sr; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179672.4]
  wire  tlb_OptimizationBarrier_38_io_y_pw; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179672.4]
  wire  tlb_OptimizationBarrier_38_io_y_px; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179672.4]
  wire  tlb_OptimizationBarrier_38_io_y_pr; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179672.4]
  wire  tlb_OptimizationBarrier_38_io_y_ppp; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179672.4]
  wire  tlb_OptimizationBarrier_38_io_y_pal; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179672.4]
  wire  tlb_OptimizationBarrier_38_io_y_paa; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179672.4]
  wire  tlb_OptimizationBarrier_38_io_y_eff; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179672.4]
  wire  tlb_OptimizationBarrier_38_io_y_c; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179672.4]
  reg [19:0] tlb_sectored_entries_0_tag; // @[TLB.scala 162:29:freechips.rocketchip.system.DefaultRV32Config.fir@176847.4]
  reg [34:0] tlb_sectored_entries_0_data_0; // @[TLB.scala 162:29:freechips.rocketchip.system.DefaultRV32Config.fir@176847.4]
  reg [34:0] tlb_sectored_entries_0_data_1; // @[TLB.scala 162:29:freechips.rocketchip.system.DefaultRV32Config.fir@176847.4]
  reg [34:0] tlb_sectored_entries_0_data_2; // @[TLB.scala 162:29:freechips.rocketchip.system.DefaultRV32Config.fir@176847.4]
  reg [34:0] tlb_sectored_entries_0_data_3; // @[TLB.scala 162:29:freechips.rocketchip.system.DefaultRV32Config.fir@176847.4]
  reg  tlb_sectored_entries_0_valid_0; // @[TLB.scala 162:29:freechips.rocketchip.system.DefaultRV32Config.fir@176847.4]
  reg  tlb_sectored_entries_0_valid_1; // @[TLB.scala 162:29:freechips.rocketchip.system.DefaultRV32Config.fir@176847.4]
  reg  tlb_sectored_entries_0_valid_2; // @[TLB.scala 162:29:freechips.rocketchip.system.DefaultRV32Config.fir@176847.4]
  reg  tlb_sectored_entries_0_valid_3; // @[TLB.scala 162:29:freechips.rocketchip.system.DefaultRV32Config.fir@176847.4]
  reg [19:0] tlb_sectored_entries_1_tag; // @[TLB.scala 162:29:freechips.rocketchip.system.DefaultRV32Config.fir@176847.4]
  reg [34:0] tlb_sectored_entries_1_data_0; // @[TLB.scala 162:29:freechips.rocketchip.system.DefaultRV32Config.fir@176847.4]
  reg [34:0] tlb_sectored_entries_1_data_1; // @[TLB.scala 162:29:freechips.rocketchip.system.DefaultRV32Config.fir@176847.4]
  reg [34:0] tlb_sectored_entries_1_data_2; // @[TLB.scala 162:29:freechips.rocketchip.system.DefaultRV32Config.fir@176847.4]
  reg [34:0] tlb_sectored_entries_1_data_3; // @[TLB.scala 162:29:freechips.rocketchip.system.DefaultRV32Config.fir@176847.4]
  reg  tlb_sectored_entries_1_valid_0; // @[TLB.scala 162:29:freechips.rocketchip.system.DefaultRV32Config.fir@176847.4]
  reg  tlb_sectored_entries_1_valid_1; // @[TLB.scala 162:29:freechips.rocketchip.system.DefaultRV32Config.fir@176847.4]
  reg  tlb_sectored_entries_1_valid_2; // @[TLB.scala 162:29:freechips.rocketchip.system.DefaultRV32Config.fir@176847.4]
  reg  tlb_sectored_entries_1_valid_3; // @[TLB.scala 162:29:freechips.rocketchip.system.DefaultRV32Config.fir@176847.4]
  reg [19:0] tlb_sectored_entries_2_tag; // @[TLB.scala 162:29:freechips.rocketchip.system.DefaultRV32Config.fir@176847.4]
  reg [34:0] tlb_sectored_entries_2_data_0; // @[TLB.scala 162:29:freechips.rocketchip.system.DefaultRV32Config.fir@176847.4]
  reg [34:0] tlb_sectored_entries_2_data_1; // @[TLB.scala 162:29:freechips.rocketchip.system.DefaultRV32Config.fir@176847.4]
  reg [34:0] tlb_sectored_entries_2_data_2; // @[TLB.scala 162:29:freechips.rocketchip.system.DefaultRV32Config.fir@176847.4]
  reg [34:0] tlb_sectored_entries_2_data_3; // @[TLB.scala 162:29:freechips.rocketchip.system.DefaultRV32Config.fir@176847.4]
  reg  tlb_sectored_entries_2_valid_0; // @[TLB.scala 162:29:freechips.rocketchip.system.DefaultRV32Config.fir@176847.4]
  reg  tlb_sectored_entries_2_valid_1; // @[TLB.scala 162:29:freechips.rocketchip.system.DefaultRV32Config.fir@176847.4]
  reg  tlb_sectored_entries_2_valid_2; // @[TLB.scala 162:29:freechips.rocketchip.system.DefaultRV32Config.fir@176847.4]
  reg  tlb_sectored_entries_2_valid_3; // @[TLB.scala 162:29:freechips.rocketchip.system.DefaultRV32Config.fir@176847.4]
  reg [19:0] tlb_sectored_entries_3_tag; // @[TLB.scala 162:29:freechips.rocketchip.system.DefaultRV32Config.fir@176847.4]
  reg [34:0] tlb_sectored_entries_3_data_0; // @[TLB.scala 162:29:freechips.rocketchip.system.DefaultRV32Config.fir@176847.4]
  reg [34:0] tlb_sectored_entries_3_data_1; // @[TLB.scala 162:29:freechips.rocketchip.system.DefaultRV32Config.fir@176847.4]
  reg [34:0] tlb_sectored_entries_3_data_2; // @[TLB.scala 162:29:freechips.rocketchip.system.DefaultRV32Config.fir@176847.4]
  reg [34:0] tlb_sectored_entries_3_data_3; // @[TLB.scala 162:29:freechips.rocketchip.system.DefaultRV32Config.fir@176847.4]
  reg  tlb_sectored_entries_3_valid_0; // @[TLB.scala 162:29:freechips.rocketchip.system.DefaultRV32Config.fir@176847.4]
  reg  tlb_sectored_entries_3_valid_1; // @[TLB.scala 162:29:freechips.rocketchip.system.DefaultRV32Config.fir@176847.4]
  reg  tlb_sectored_entries_3_valid_2; // @[TLB.scala 162:29:freechips.rocketchip.system.DefaultRV32Config.fir@176847.4]
  reg  tlb_sectored_entries_3_valid_3; // @[TLB.scala 162:29:freechips.rocketchip.system.DefaultRV32Config.fir@176847.4]
  reg [19:0] tlb_sectored_entries_4_tag; // @[TLB.scala 162:29:freechips.rocketchip.system.DefaultRV32Config.fir@176847.4]
  reg [34:0] tlb_sectored_entries_4_data_0; // @[TLB.scala 162:29:freechips.rocketchip.system.DefaultRV32Config.fir@176847.4]
  reg [34:0] tlb_sectored_entries_4_data_1; // @[TLB.scala 162:29:freechips.rocketchip.system.DefaultRV32Config.fir@176847.4]
  reg [34:0] tlb_sectored_entries_4_data_2; // @[TLB.scala 162:29:freechips.rocketchip.system.DefaultRV32Config.fir@176847.4]
  reg [34:0] tlb_sectored_entries_4_data_3; // @[TLB.scala 162:29:freechips.rocketchip.system.DefaultRV32Config.fir@176847.4]
  reg  tlb_sectored_entries_4_valid_0; // @[TLB.scala 162:29:freechips.rocketchip.system.DefaultRV32Config.fir@176847.4]
  reg  tlb_sectored_entries_4_valid_1; // @[TLB.scala 162:29:freechips.rocketchip.system.DefaultRV32Config.fir@176847.4]
  reg  tlb_sectored_entries_4_valid_2; // @[TLB.scala 162:29:freechips.rocketchip.system.DefaultRV32Config.fir@176847.4]
  reg  tlb_sectored_entries_4_valid_3; // @[TLB.scala 162:29:freechips.rocketchip.system.DefaultRV32Config.fir@176847.4]
  reg [19:0] tlb_sectored_entries_5_tag; // @[TLB.scala 162:29:freechips.rocketchip.system.DefaultRV32Config.fir@176847.4]
  reg [34:0] tlb_sectored_entries_5_data_0; // @[TLB.scala 162:29:freechips.rocketchip.system.DefaultRV32Config.fir@176847.4]
  reg [34:0] tlb_sectored_entries_5_data_1; // @[TLB.scala 162:29:freechips.rocketchip.system.DefaultRV32Config.fir@176847.4]
  reg [34:0] tlb_sectored_entries_5_data_2; // @[TLB.scala 162:29:freechips.rocketchip.system.DefaultRV32Config.fir@176847.4]
  reg [34:0] tlb_sectored_entries_5_data_3; // @[TLB.scala 162:29:freechips.rocketchip.system.DefaultRV32Config.fir@176847.4]
  reg  tlb_sectored_entries_5_valid_0; // @[TLB.scala 162:29:freechips.rocketchip.system.DefaultRV32Config.fir@176847.4]
  reg  tlb_sectored_entries_5_valid_1; // @[TLB.scala 162:29:freechips.rocketchip.system.DefaultRV32Config.fir@176847.4]
  reg  tlb_sectored_entries_5_valid_2; // @[TLB.scala 162:29:freechips.rocketchip.system.DefaultRV32Config.fir@176847.4]
  reg  tlb_sectored_entries_5_valid_3; // @[TLB.scala 162:29:freechips.rocketchip.system.DefaultRV32Config.fir@176847.4]
  reg [19:0] tlb_sectored_entries_6_tag; // @[TLB.scala 162:29:freechips.rocketchip.system.DefaultRV32Config.fir@176847.4]
  reg [34:0] tlb_sectored_entries_6_data_0; // @[TLB.scala 162:29:freechips.rocketchip.system.DefaultRV32Config.fir@176847.4]
  reg [34:0] tlb_sectored_entries_6_data_1; // @[TLB.scala 162:29:freechips.rocketchip.system.DefaultRV32Config.fir@176847.4]
  reg [34:0] tlb_sectored_entries_6_data_2; // @[TLB.scala 162:29:freechips.rocketchip.system.DefaultRV32Config.fir@176847.4]
  reg [34:0] tlb_sectored_entries_6_data_3; // @[TLB.scala 162:29:freechips.rocketchip.system.DefaultRV32Config.fir@176847.4]
  reg  tlb_sectored_entries_6_valid_0; // @[TLB.scala 162:29:freechips.rocketchip.system.DefaultRV32Config.fir@176847.4]
  reg  tlb_sectored_entries_6_valid_1; // @[TLB.scala 162:29:freechips.rocketchip.system.DefaultRV32Config.fir@176847.4]
  reg  tlb_sectored_entries_6_valid_2; // @[TLB.scala 162:29:freechips.rocketchip.system.DefaultRV32Config.fir@176847.4]
  reg  tlb_sectored_entries_6_valid_3; // @[TLB.scala 162:29:freechips.rocketchip.system.DefaultRV32Config.fir@176847.4]
  reg [19:0] tlb_sectored_entries_7_tag; // @[TLB.scala 162:29:freechips.rocketchip.system.DefaultRV32Config.fir@176847.4]
  reg [34:0] tlb_sectored_entries_7_data_0; // @[TLB.scala 162:29:freechips.rocketchip.system.DefaultRV32Config.fir@176847.4]
  reg [34:0] tlb_sectored_entries_7_data_1; // @[TLB.scala 162:29:freechips.rocketchip.system.DefaultRV32Config.fir@176847.4]
  reg [34:0] tlb_sectored_entries_7_data_2; // @[TLB.scala 162:29:freechips.rocketchip.system.DefaultRV32Config.fir@176847.4]
  reg [34:0] tlb_sectored_entries_7_data_3; // @[TLB.scala 162:29:freechips.rocketchip.system.DefaultRV32Config.fir@176847.4]
  reg  tlb_sectored_entries_7_valid_0; // @[TLB.scala 162:29:freechips.rocketchip.system.DefaultRV32Config.fir@176847.4]
  reg  tlb_sectored_entries_7_valid_1; // @[TLB.scala 162:29:freechips.rocketchip.system.DefaultRV32Config.fir@176847.4]
  reg  tlb_sectored_entries_7_valid_2; // @[TLB.scala 162:29:freechips.rocketchip.system.DefaultRV32Config.fir@176847.4]
  reg  tlb_sectored_entries_7_valid_3; // @[TLB.scala 162:29:freechips.rocketchip.system.DefaultRV32Config.fir@176847.4]
  reg [19:0] tlb_superpage_entries_0_tag; // @[TLB.scala 163:30:freechips.rocketchip.system.DefaultRV32Config.fir@176848.4]
  reg [34:0] tlb_superpage_entries_0_data_0; // @[TLB.scala 163:30:freechips.rocketchip.system.DefaultRV32Config.fir@176848.4]
  reg  tlb_superpage_entries_0_valid_0; // @[TLB.scala 163:30:freechips.rocketchip.system.DefaultRV32Config.fir@176848.4]
  reg [19:0] tlb_superpage_entries_1_tag; // @[TLB.scala 163:30:freechips.rocketchip.system.DefaultRV32Config.fir@176848.4]
  reg [34:0] tlb_superpage_entries_1_data_0; // @[TLB.scala 163:30:freechips.rocketchip.system.DefaultRV32Config.fir@176848.4]
  reg  tlb_superpage_entries_1_valid_0; // @[TLB.scala 163:30:freechips.rocketchip.system.DefaultRV32Config.fir@176848.4]
  reg [19:0] tlb_superpage_entries_2_tag; // @[TLB.scala 163:30:freechips.rocketchip.system.DefaultRV32Config.fir@176848.4]
  reg [34:0] tlb_superpage_entries_2_data_0; // @[TLB.scala 163:30:freechips.rocketchip.system.DefaultRV32Config.fir@176848.4]
  reg  tlb_superpage_entries_2_valid_0; // @[TLB.scala 163:30:freechips.rocketchip.system.DefaultRV32Config.fir@176848.4]
  reg [19:0] tlb_superpage_entries_3_tag; // @[TLB.scala 163:30:freechips.rocketchip.system.DefaultRV32Config.fir@176848.4]
  reg [34:0] tlb_superpage_entries_3_data_0; // @[TLB.scala 163:30:freechips.rocketchip.system.DefaultRV32Config.fir@176848.4]
  reg  tlb_superpage_entries_3_valid_0; // @[TLB.scala 163:30:freechips.rocketchip.system.DefaultRV32Config.fir@176848.4]
  reg  tlb_special_entry_level; // @[TLB.scala 164:56:freechips.rocketchip.system.DefaultRV32Config.fir@176849.4]
  reg [19:0] tlb_special_entry_tag; // @[TLB.scala 164:56:freechips.rocketchip.system.DefaultRV32Config.fir@176849.4]
  reg [34:0] tlb_special_entry_data_0; // @[TLB.scala 164:56:freechips.rocketchip.system.DefaultRV32Config.fir@176849.4]
  reg  tlb_special_entry_valid_0; // @[TLB.scala 164:56:freechips.rocketchip.system.DefaultRV32Config.fir@176849.4]
  reg [1:0] tlb_state; // @[TLB.scala 169:18:freechips.rocketchip.system.DefaultRV32Config.fir@176850.4]
  reg [19:0] tlb_r_refill_tag; // @[TLB.scala 170:25:freechips.rocketchip.system.DefaultRV32Config.fir@176851.4]
  reg [1:0] tlb_r_superpage_repl_addr; // @[TLB.scala 171:34:freechips.rocketchip.system.DefaultRV32Config.fir@176852.4]
  reg [2:0] tlb_r_sectored_repl_addr; // @[TLB.scala 172:33:freechips.rocketchip.system.DefaultRV32Config.fir@176853.4]
  reg [2:0] tlb_r_sectored_hit_addr; // @[TLB.scala 173:32:freechips.rocketchip.system.DefaultRV32Config.fir@176854.4]
  reg  tlb_r_sectored_hit; // @[TLB.scala 174:27:freechips.rocketchip.system.DefaultRV32Config.fir@176855.4]
  wire  tlb_priv_s; // @[TLB.scala 177:20:freechips.rocketchip.system.DefaultRV32Config.fir@176856.4]
  wire  tlb_priv_uses_vm; // @[TLB.scala 178:27:freechips.rocketchip.system.DefaultRV32Config.fir@176857.4]
  wire  tlb__T_2; // @[TLB.scala 179:83:freechips.rocketchip.system.DefaultRV32Config.fir@176860.4]
  wire  tlb__T_3; // @[TLB.scala 179:102:freechips.rocketchip.system.DefaultRV32Config.fir@176861.4]
  wire  tlb_vm_enabled; // @[TLB.scala 179:99:freechips.rocketchip.system.DefaultRV32Config.fir@176862.4]
  wire [19:0] tlb_vpn; // @[TLB.scala 182:30:freechips.rocketchip.system.DefaultRV32Config.fir@176863.4]
  wire [19:0] tlb_refill_ppn; // @[TLB.scala 183:44:freechips.rocketchip.system.DefaultRV32Config.fir@176864.4]
  wire  tlb__T_4; // @[package.scala 15:47:freechips.rocketchip.system.DefaultRV32Config.fir@176866.4]
  wire  tlb__T_5; // @[package.scala 15:47:freechips.rocketchip.system.DefaultRV32Config.fir@176867.4]
  wire  tlb_invalidate_refill; // @[package.scala 64:59:freechips.rocketchip.system.DefaultRV32Config.fir@176868.4]
  wire  tlb__T_22; // @[TLB.scala 86:77:freechips.rocketchip.system.DefaultRV32Config.fir@176901.4]
  wire [9:0] tlb__T_25; // @[TLB.scala 106:26:freechips.rocketchip.system.DefaultRV32Config.fir@176912.4]
  wire  tlb__T_26; // @[TLB.scala 108:28:freechips.rocketchip.system.DefaultRV32Config.fir@176913.4]
  wire [19:0] tlb__T_28; // @[TLB.scala 109:28:freechips.rocketchip.system.DefaultRV32Config.fir@176915.4]
  wire [19:0] tlb__T_29; // @[TLB.scala 109:47:freechips.rocketchip.system.DefaultRV32Config.fir@176916.4]
  wire [9:0] tlb__T_30; // @[TLB.scala 109:58:freechips.rocketchip.system.DefaultRV32Config.fir@176917.4]
  wire [19:0] tlb__T_31; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@176918.4]
  wire [19:0] tlb__T_32; // @[TLB.scala 187:123:freechips.rocketchip.system.DefaultRV32Config.fir@176919.4]
  wire [19:0] tlb__T_33; // @[TLB.scala 187:20:freechips.rocketchip.system.DefaultRV32Config.fir@176920.4]
  wire [19:0] tlb_mpu_ppn; // @[TLB.scala 186:20:freechips.rocketchip.system.DefaultRV32Config.fir@176921.4]
  wire [11:0] tlb__T_34; // @[TLB.scala 188:52:freechips.rocketchip.system.DefaultRV32Config.fir@176922.4]
  wire [31:0] tlb_mpu_physaddr; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@176923.4]
  wire  tlb__T_35; // @[TLB.scala 189:56:freechips.rocketchip.system.DefaultRV32Config.fir@176924.4]
  wire [2:0] tlb__T_37; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@176926.4]
  wire [2:0] tlb_mpu_priv; // @[TLB.scala 189:27:freechips.rocketchip.system.DefaultRV32Config.fir@176927.4]
  wire [31:0] tlb__T_38; // @[Parameters.scala 137:31:freechips.rocketchip.system.DefaultRV32Config.fir@176943.4]
  wire [32:0] tlb__T_39; // @[Parameters.scala 137:49:freechips.rocketchip.system.DefaultRV32Config.fir@176944.4]
  wire [32:0] tlb__T_41; // @[Parameters.scala 137:52:freechips.rocketchip.system.DefaultRV32Config.fir@176946.4]
  wire  tlb__T_42; // @[Parameters.scala 137:67:freechips.rocketchip.system.DefaultRV32Config.fir@176947.4]
  wire [31:0] tlb__T_43; // @[Parameters.scala 137:31:freechips.rocketchip.system.DefaultRV32Config.fir@176948.4]
  wire [32:0] tlb__T_44; // @[Parameters.scala 137:49:freechips.rocketchip.system.DefaultRV32Config.fir@176949.4]
  wire [32:0] tlb__T_46; // @[Parameters.scala 137:52:freechips.rocketchip.system.DefaultRV32Config.fir@176951.4]
  wire  tlb__T_47; // @[Parameters.scala 137:67:freechips.rocketchip.system.DefaultRV32Config.fir@176952.4]
  wire [31:0] tlb__T_48; // @[Parameters.scala 137:31:freechips.rocketchip.system.DefaultRV32Config.fir@176953.4]
  wire [32:0] tlb__T_49; // @[Parameters.scala 137:49:freechips.rocketchip.system.DefaultRV32Config.fir@176954.4]
  wire [32:0] tlb__T_51; // @[Parameters.scala 137:52:freechips.rocketchip.system.DefaultRV32Config.fir@176956.4]
  wire  tlb__T_52; // @[Parameters.scala 137:67:freechips.rocketchip.system.DefaultRV32Config.fir@176957.4]
  wire [32:0] tlb__T_54; // @[Parameters.scala 137:49:freechips.rocketchip.system.DefaultRV32Config.fir@176959.4]
  wire [32:0] tlb__T_56; // @[Parameters.scala 137:52:freechips.rocketchip.system.DefaultRV32Config.fir@176961.4]
  wire  tlb__T_57; // @[Parameters.scala 137:67:freechips.rocketchip.system.DefaultRV32Config.fir@176962.4]
  wire [31:0] tlb__T_58; // @[Parameters.scala 137:31:freechips.rocketchip.system.DefaultRV32Config.fir@176963.4]
  wire [32:0] tlb__T_59; // @[Parameters.scala 137:49:freechips.rocketchip.system.DefaultRV32Config.fir@176964.4]
  wire [32:0] tlb__T_61; // @[Parameters.scala 137:52:freechips.rocketchip.system.DefaultRV32Config.fir@176966.4]
  wire  tlb__T_62; // @[Parameters.scala 137:67:freechips.rocketchip.system.DefaultRV32Config.fir@176967.4]
  wire [31:0] tlb__T_63; // @[Parameters.scala 137:31:freechips.rocketchip.system.DefaultRV32Config.fir@176968.4]
  wire [32:0] tlb__T_64; // @[Parameters.scala 137:49:freechips.rocketchip.system.DefaultRV32Config.fir@176969.4]
  wire [32:0] tlb__T_66; // @[Parameters.scala 137:52:freechips.rocketchip.system.DefaultRV32Config.fir@176971.4]
  wire  tlb__T_67; // @[Parameters.scala 137:67:freechips.rocketchip.system.DefaultRV32Config.fir@176972.4]
  wire [31:0] tlb__T_68; // @[Parameters.scala 137:31:freechips.rocketchip.system.DefaultRV32Config.fir@176973.4]
  wire [32:0] tlb__T_69; // @[Parameters.scala 137:49:freechips.rocketchip.system.DefaultRV32Config.fir@176974.4]
  wire [32:0] tlb__T_71; // @[Parameters.scala 137:52:freechips.rocketchip.system.DefaultRV32Config.fir@176976.4]
  wire  tlb__T_72; // @[Parameters.scala 137:67:freechips.rocketchip.system.DefaultRV32Config.fir@176977.4]
  wire  tlb__T_74; // @[TLB.scala 195:67:freechips.rocketchip.system.DefaultRV32Config.fir@176987.4]
  wire  tlb__T_75; // @[TLB.scala 195:67:freechips.rocketchip.system.DefaultRV32Config.fir@176988.4]
  wire  tlb__T_76; // @[TLB.scala 195:67:freechips.rocketchip.system.DefaultRV32Config.fir@176989.4]
  wire  tlb__T_77; // @[TLB.scala 195:67:freechips.rocketchip.system.DefaultRV32Config.fir@176990.4]
  wire  tlb__T_78; // @[TLB.scala 195:67:freechips.rocketchip.system.DefaultRV32Config.fir@176991.4]
  wire  tlb_legal_address; // @[TLB.scala 195:67:freechips.rocketchip.system.DefaultRV32Config.fir@176992.4]
  wire [32:0] tlb__T_87; // @[Parameters.scala 137:52:freechips.rocketchip.system.DefaultRV32Config.fir@177001.4]
  wire  tlb__T_88; // @[Parameters.scala 137:67:freechips.rocketchip.system.DefaultRV32Config.fir@177002.4]
  wire  tlb__T_93; // @[TLB.scala 197:19:freechips.rocketchip.system.DefaultRV32Config.fir@177008.4]
  wire [31:0] tlb__T_148; // @[Parameters.scala 137:31:freechips.rocketchip.system.DefaultRV32Config.fir@177065.4]
  wire [32:0] tlb__T_149; // @[Parameters.scala 137:49:freechips.rocketchip.system.DefaultRV32Config.fir@177066.4]
  wire [32:0] tlb__T_151; // @[Parameters.scala 137:52:freechips.rocketchip.system.DefaultRV32Config.fir@177068.4]
  wire  tlb__T_152; // @[Parameters.scala 137:67:freechips.rocketchip.system.DefaultRV32Config.fir@177069.4]
  wire [32:0] tlb__T_165; // @[Parameters.scala 137:52:freechips.rocketchip.system.DefaultRV32Config.fir@177082.4]
  wire  tlb__T_166; // @[Parameters.scala 137:67:freechips.rocketchip.system.DefaultRV32Config.fir@177083.4]
  wire  tlb__T_173; // @[TLBPermissions.scala 82:66:freechips.rocketchip.system.DefaultRV32Config.fir@177090.4]
  wire  tlb__T_186; // @[TLB.scala 200:39:freechips.rocketchip.system.DefaultRV32Config.fir@177103.4]
  wire  tlb_deny_access_to_debug; // @[TLB.scala 200:48:freechips.rocketchip.system.DefaultRV32Config.fir@177109.4]
  wire  tlb__T_198; // @[TLB.scala 201:44:freechips.rocketchip.system.DefaultRV32Config.fir@177116.4]
  wire  tlb__T_199; // @[TLB.scala 201:41:freechips.rocketchip.system.DefaultRV32Config.fir@177117.4]
  wire  tlb_prot_r; // @[TLB.scala 201:66:freechips.rocketchip.system.DefaultRV32Config.fir@177118.4]
  wire [31:0] tlb__T_210; // @[Parameters.scala 137:31:freechips.rocketchip.system.DefaultRV32Config.fir@177129.4]
  wire [32:0] tlb__T_211; // @[Parameters.scala 137:49:freechips.rocketchip.system.DefaultRV32Config.fir@177130.4]
  wire [32:0] tlb__T_213; // @[Parameters.scala 137:52:freechips.rocketchip.system.DefaultRV32Config.fir@177132.4]
  wire  tlb__T_214; // @[Parameters.scala 137:67:freechips.rocketchip.system.DefaultRV32Config.fir@177133.4]
  wire [32:0] tlb__T_218; // @[Parameters.scala 137:52:freechips.rocketchip.system.DefaultRV32Config.fir@177137.4]
  wire  tlb__T_219; // @[Parameters.scala 137:67:freechips.rocketchip.system.DefaultRV32Config.fir@177138.4]
  wire  tlb__T_221; // @[Parameters.scala 528:89:freechips.rocketchip.system.DefaultRV32Config.fir@177140.4]
  wire  tlb__T_222; // @[Parameters.scala 528:89:freechips.rocketchip.system.DefaultRV32Config.fir@177141.4]
  wire  tlb__T_232; // @[TLB.scala 197:19:freechips.rocketchip.system.DefaultRV32Config.fir@177152.4]
  wire  tlb__T_234; // @[TLB.scala 202:45:freechips.rocketchip.system.DefaultRV32Config.fir@177154.4]
  wire  tlb_prot_w; // @[TLB.scala 202:70:freechips.rocketchip.system.DefaultRV32Config.fir@177155.4]
  wire  tlb_prot_al; // @[TLB.scala 197:19:freechips.rocketchip.system.DefaultRV32Config.fir@177223.4]
  wire [32:0] tlb__T_334; // @[Parameters.scala 137:52:freechips.rocketchip.system.DefaultRV32Config.fir@177261.4]
  wire  tlb__T_335; // @[Parameters.scala 137:67:freechips.rocketchip.system.DefaultRV32Config.fir@177262.4]
  wire  tlb__T_346; // @[Parameters.scala 528:89:freechips.rocketchip.system.DefaultRV32Config.fir@177273.4]
  wire  tlb__T_347; // @[Parameters.scala 528:89:freechips.rocketchip.system.DefaultRV32Config.fir@177274.4]
  wire  tlb__T_363; // @[TLB.scala 197:19:freechips.rocketchip.system.DefaultRV32Config.fir@177291.4]
  wire  tlb__T_365; // @[TLB.scala 206:40:freechips.rocketchip.system.DefaultRV32Config.fir@177293.4]
  wire  tlb_prot_x; // @[TLB.scala 206:65:freechips.rocketchip.system.DefaultRV32Config.fir@177294.4]
  wire [32:0] tlb__T_386; // @[Parameters.scala 137:52:freechips.rocketchip.system.DefaultRV32Config.fir@177315.4]
  wire  tlb__T_387; // @[Parameters.scala 137:67:freechips.rocketchip.system.DefaultRV32Config.fir@177316.4]
  wire [32:0] tlb__T_391; // @[Parameters.scala 137:52:freechips.rocketchip.system.DefaultRV32Config.fir@177320.4]
  wire  tlb__T_392; // @[Parameters.scala 137:67:freechips.rocketchip.system.DefaultRV32Config.fir@177321.4]
  wire  tlb__T_403; // @[Parameters.scala 528:89:freechips.rocketchip.system.DefaultRV32Config.fir@177332.4]
  wire  tlb__T_404; // @[Parameters.scala 528:89:freechips.rocketchip.system.DefaultRV32Config.fir@177333.4]
  wire  tlb__T_405; // @[Parameters.scala 528:89:freechips.rocketchip.system.DefaultRV32Config.fir@177334.4]
  wire  tlb_prot_eff; // @[TLB.scala 197:19:freechips.rocketchip.system.DefaultRV32Config.fir@177340.4]
  wire  tlb__T_410; // @[package.scala 64:59:freechips.rocketchip.system.DefaultRV32Config.fir@177341.4]
  wire  tlb__T_411; // @[package.scala 64:59:freechips.rocketchip.system.DefaultRV32Config.fir@177342.4]
  wire  tlb__T_412; // @[package.scala 64:59:freechips.rocketchip.system.DefaultRV32Config.fir@177343.4]
  wire [19:0] tlb__T_413; // @[TLB.scala 88:41:freechips.rocketchip.system.DefaultRV32Config.fir@177344.4]
  wire [17:0] tlb__T_414; // @[TLB.scala 88:48:freechips.rocketchip.system.DefaultRV32Config.fir@177345.4]
  wire  tlb__T_415; // @[TLB.scala 88:66:freechips.rocketchip.system.DefaultRV32Config.fir@177346.4]
  wire  tlb_sector_hits_0; // @[TLB.scala 87:40:freechips.rocketchip.system.DefaultRV32Config.fir@177347.4]
  wire  tlb__T_416; // @[package.scala 64:59:freechips.rocketchip.system.DefaultRV32Config.fir@177348.4]
  wire  tlb__T_417; // @[package.scala 64:59:freechips.rocketchip.system.DefaultRV32Config.fir@177349.4]
  wire  tlb__T_418; // @[package.scala 64:59:freechips.rocketchip.system.DefaultRV32Config.fir@177350.4]
  wire [19:0] tlb__T_419; // @[TLB.scala 88:41:freechips.rocketchip.system.DefaultRV32Config.fir@177351.4]
  wire [17:0] tlb__T_420; // @[TLB.scala 88:48:freechips.rocketchip.system.DefaultRV32Config.fir@177352.4]
  wire  tlb__T_421; // @[TLB.scala 88:66:freechips.rocketchip.system.DefaultRV32Config.fir@177353.4]
  wire  tlb_sector_hits_1; // @[TLB.scala 87:40:freechips.rocketchip.system.DefaultRV32Config.fir@177354.4]
  wire  tlb__T_422; // @[package.scala 64:59:freechips.rocketchip.system.DefaultRV32Config.fir@177355.4]
  wire  tlb__T_423; // @[package.scala 64:59:freechips.rocketchip.system.DefaultRV32Config.fir@177356.4]
  wire  tlb__T_424; // @[package.scala 64:59:freechips.rocketchip.system.DefaultRV32Config.fir@177357.4]
  wire [19:0] tlb__T_425; // @[TLB.scala 88:41:freechips.rocketchip.system.DefaultRV32Config.fir@177358.4]
  wire [17:0] tlb__T_426; // @[TLB.scala 88:48:freechips.rocketchip.system.DefaultRV32Config.fir@177359.4]
  wire  tlb__T_427; // @[TLB.scala 88:66:freechips.rocketchip.system.DefaultRV32Config.fir@177360.4]
  wire  tlb_sector_hits_2; // @[TLB.scala 87:40:freechips.rocketchip.system.DefaultRV32Config.fir@177361.4]
  wire  tlb__T_428; // @[package.scala 64:59:freechips.rocketchip.system.DefaultRV32Config.fir@177362.4]
  wire  tlb__T_429; // @[package.scala 64:59:freechips.rocketchip.system.DefaultRV32Config.fir@177363.4]
  wire  tlb__T_430; // @[package.scala 64:59:freechips.rocketchip.system.DefaultRV32Config.fir@177364.4]
  wire [19:0] tlb__T_431; // @[TLB.scala 88:41:freechips.rocketchip.system.DefaultRV32Config.fir@177365.4]
  wire [17:0] tlb__T_432; // @[TLB.scala 88:48:freechips.rocketchip.system.DefaultRV32Config.fir@177366.4]
  wire  tlb__T_433; // @[TLB.scala 88:66:freechips.rocketchip.system.DefaultRV32Config.fir@177367.4]
  wire  tlb_sector_hits_3; // @[TLB.scala 87:40:freechips.rocketchip.system.DefaultRV32Config.fir@177368.4]
  wire  tlb__T_434; // @[package.scala 64:59:freechips.rocketchip.system.DefaultRV32Config.fir@177369.4]
  wire  tlb__T_435; // @[package.scala 64:59:freechips.rocketchip.system.DefaultRV32Config.fir@177370.4]
  wire  tlb__T_436; // @[package.scala 64:59:freechips.rocketchip.system.DefaultRV32Config.fir@177371.4]
  wire [19:0] tlb__T_437; // @[TLB.scala 88:41:freechips.rocketchip.system.DefaultRV32Config.fir@177372.4]
  wire [17:0] tlb__T_438; // @[TLB.scala 88:48:freechips.rocketchip.system.DefaultRV32Config.fir@177373.4]
  wire  tlb__T_439; // @[TLB.scala 88:66:freechips.rocketchip.system.DefaultRV32Config.fir@177374.4]
  wire  tlb_sector_hits_4; // @[TLB.scala 87:40:freechips.rocketchip.system.DefaultRV32Config.fir@177375.4]
  wire  tlb__T_440; // @[package.scala 64:59:freechips.rocketchip.system.DefaultRV32Config.fir@177376.4]
  wire  tlb__T_441; // @[package.scala 64:59:freechips.rocketchip.system.DefaultRV32Config.fir@177377.4]
  wire  tlb__T_442; // @[package.scala 64:59:freechips.rocketchip.system.DefaultRV32Config.fir@177378.4]
  wire [19:0] tlb__T_443; // @[TLB.scala 88:41:freechips.rocketchip.system.DefaultRV32Config.fir@177379.4]
  wire [17:0] tlb__T_444; // @[TLB.scala 88:48:freechips.rocketchip.system.DefaultRV32Config.fir@177380.4]
  wire  tlb__T_445; // @[TLB.scala 88:66:freechips.rocketchip.system.DefaultRV32Config.fir@177381.4]
  wire  tlb_sector_hits_5; // @[TLB.scala 87:40:freechips.rocketchip.system.DefaultRV32Config.fir@177382.4]
  wire  tlb__T_446; // @[package.scala 64:59:freechips.rocketchip.system.DefaultRV32Config.fir@177383.4]
  wire  tlb__T_447; // @[package.scala 64:59:freechips.rocketchip.system.DefaultRV32Config.fir@177384.4]
  wire  tlb__T_448; // @[package.scala 64:59:freechips.rocketchip.system.DefaultRV32Config.fir@177385.4]
  wire [19:0] tlb__T_449; // @[TLB.scala 88:41:freechips.rocketchip.system.DefaultRV32Config.fir@177386.4]
  wire [17:0] tlb__T_450; // @[TLB.scala 88:48:freechips.rocketchip.system.DefaultRV32Config.fir@177387.4]
  wire  tlb__T_451; // @[TLB.scala 88:66:freechips.rocketchip.system.DefaultRV32Config.fir@177388.4]
  wire  tlb_sector_hits_6; // @[TLB.scala 87:40:freechips.rocketchip.system.DefaultRV32Config.fir@177389.4]
  wire  tlb__T_452; // @[package.scala 64:59:freechips.rocketchip.system.DefaultRV32Config.fir@177390.4]
  wire  tlb__T_453; // @[package.scala 64:59:freechips.rocketchip.system.DefaultRV32Config.fir@177391.4]
  wire  tlb__T_454; // @[package.scala 64:59:freechips.rocketchip.system.DefaultRV32Config.fir@177392.4]
  wire [19:0] tlb__T_455; // @[TLB.scala 88:41:freechips.rocketchip.system.DefaultRV32Config.fir@177393.4]
  wire [17:0] tlb__T_456; // @[TLB.scala 88:48:freechips.rocketchip.system.DefaultRV32Config.fir@177394.4]
  wire  tlb__T_457; // @[TLB.scala 88:66:freechips.rocketchip.system.DefaultRV32Config.fir@177395.4]
  wire  tlb_sector_hits_7; // @[TLB.scala 87:40:freechips.rocketchip.system.DefaultRV32Config.fir@177396.4]
  wire [9:0] tlb__T_460; // @[TLB.scala 95:46:freechips.rocketchip.system.DefaultRV32Config.fir@177399.4]
  wire [9:0] tlb__T_461; // @[TLB.scala 95:84:freechips.rocketchip.system.DefaultRV32Config.fir@177400.4]
  wire  tlb__T_462; // @[TLB.scala 95:77:freechips.rocketchip.system.DefaultRV32Config.fir@177401.4]
  wire  tlb__T_464; // @[TLB.scala 95:29:freechips.rocketchip.system.DefaultRV32Config.fir@177403.4]
  wire [9:0] tlb__T_468; // @[TLB.scala 95:84:freechips.rocketchip.system.DefaultRV32Config.fir@177407.4]
  wire [9:0] tlb__T_473; // @[TLB.scala 95:46:freechips.rocketchip.system.DefaultRV32Config.fir@177413.4]
  wire  tlb__T_475; // @[TLB.scala 95:77:freechips.rocketchip.system.DefaultRV32Config.fir@177415.4]
  wire  tlb__T_477; // @[TLB.scala 95:29:freechips.rocketchip.system.DefaultRV32Config.fir@177417.4]
  wire [9:0] tlb__T_486; // @[TLB.scala 95:46:freechips.rocketchip.system.DefaultRV32Config.fir@177427.4]
  wire  tlb__T_488; // @[TLB.scala 95:77:freechips.rocketchip.system.DefaultRV32Config.fir@177429.4]
  wire  tlb__T_490; // @[TLB.scala 95:29:freechips.rocketchip.system.DefaultRV32Config.fir@177431.4]
  wire [9:0] tlb__T_499; // @[TLB.scala 95:46:freechips.rocketchip.system.DefaultRV32Config.fir@177441.4]
  wire  tlb__T_501; // @[TLB.scala 95:77:freechips.rocketchip.system.DefaultRV32Config.fir@177443.4]
  wire  tlb__T_503; // @[TLB.scala 95:29:freechips.rocketchip.system.DefaultRV32Config.fir@177445.4]
  wire [1:0] tlb__T_510; // @[package.scala 138:13:freechips.rocketchip.system.DefaultRV32Config.fir@177453.4]
  wire  tlb__GEN_1; // @[TLB.scala 100:18:freechips.rocketchip.system.DefaultRV32Config.fir@177457.4]
  wire  tlb__GEN_2; // @[TLB.scala 100:18:freechips.rocketchip.system.DefaultRV32Config.fir@177457.4]
  wire  tlb__GEN_3; // @[TLB.scala 100:18:freechips.rocketchip.system.DefaultRV32Config.fir@177457.4]
  wire  tlb__T_514; // @[TLB.scala 100:18:freechips.rocketchip.system.DefaultRV32Config.fir@177457.4]
  wire  tlb_hitsVec_0; // @[TLB.scala 211:44:freechips.rocketchip.system.DefaultRV32Config.fir@177458.4]
  wire  tlb__GEN_5; // @[TLB.scala 100:18:freechips.rocketchip.system.DefaultRV32Config.fir@177463.4]
  wire  tlb__GEN_6; // @[TLB.scala 100:18:freechips.rocketchip.system.DefaultRV32Config.fir@177463.4]
  wire  tlb__GEN_7; // @[TLB.scala 100:18:freechips.rocketchip.system.DefaultRV32Config.fir@177463.4]
  wire  tlb__T_519; // @[TLB.scala 100:18:freechips.rocketchip.system.DefaultRV32Config.fir@177463.4]
  wire  tlb_hitsVec_1; // @[TLB.scala 211:44:freechips.rocketchip.system.DefaultRV32Config.fir@177464.4]
  wire  tlb__GEN_9; // @[TLB.scala 100:18:freechips.rocketchip.system.DefaultRV32Config.fir@177469.4]
  wire  tlb__GEN_10; // @[TLB.scala 100:18:freechips.rocketchip.system.DefaultRV32Config.fir@177469.4]
  wire  tlb__GEN_11; // @[TLB.scala 100:18:freechips.rocketchip.system.DefaultRV32Config.fir@177469.4]
  wire  tlb__T_524; // @[TLB.scala 100:18:freechips.rocketchip.system.DefaultRV32Config.fir@177469.4]
  wire  tlb_hitsVec_2; // @[TLB.scala 211:44:freechips.rocketchip.system.DefaultRV32Config.fir@177470.4]
  wire  tlb__GEN_13; // @[TLB.scala 100:18:freechips.rocketchip.system.DefaultRV32Config.fir@177475.4]
  wire  tlb__GEN_14; // @[TLB.scala 100:18:freechips.rocketchip.system.DefaultRV32Config.fir@177475.4]
  wire  tlb__GEN_15; // @[TLB.scala 100:18:freechips.rocketchip.system.DefaultRV32Config.fir@177475.4]
  wire  tlb__T_529; // @[TLB.scala 100:18:freechips.rocketchip.system.DefaultRV32Config.fir@177475.4]
  wire  tlb_hitsVec_3; // @[TLB.scala 211:44:freechips.rocketchip.system.DefaultRV32Config.fir@177476.4]
  wire  tlb__GEN_17; // @[TLB.scala 100:18:freechips.rocketchip.system.DefaultRV32Config.fir@177481.4]
  wire  tlb__GEN_18; // @[TLB.scala 100:18:freechips.rocketchip.system.DefaultRV32Config.fir@177481.4]
  wire  tlb__GEN_19; // @[TLB.scala 100:18:freechips.rocketchip.system.DefaultRV32Config.fir@177481.4]
  wire  tlb__T_534; // @[TLB.scala 100:18:freechips.rocketchip.system.DefaultRV32Config.fir@177481.4]
  wire  tlb_hitsVec_4; // @[TLB.scala 211:44:freechips.rocketchip.system.DefaultRV32Config.fir@177482.4]
  wire  tlb__GEN_21; // @[TLB.scala 100:18:freechips.rocketchip.system.DefaultRV32Config.fir@177487.4]
  wire  tlb__GEN_22; // @[TLB.scala 100:18:freechips.rocketchip.system.DefaultRV32Config.fir@177487.4]
  wire  tlb__GEN_23; // @[TLB.scala 100:18:freechips.rocketchip.system.DefaultRV32Config.fir@177487.4]
  wire  tlb__T_539; // @[TLB.scala 100:18:freechips.rocketchip.system.DefaultRV32Config.fir@177487.4]
  wire  tlb_hitsVec_5; // @[TLB.scala 211:44:freechips.rocketchip.system.DefaultRV32Config.fir@177488.4]
  wire  tlb__GEN_25; // @[TLB.scala 100:18:freechips.rocketchip.system.DefaultRV32Config.fir@177493.4]
  wire  tlb__GEN_26; // @[TLB.scala 100:18:freechips.rocketchip.system.DefaultRV32Config.fir@177493.4]
  wire  tlb__GEN_27; // @[TLB.scala 100:18:freechips.rocketchip.system.DefaultRV32Config.fir@177493.4]
  wire  tlb__T_544; // @[TLB.scala 100:18:freechips.rocketchip.system.DefaultRV32Config.fir@177493.4]
  wire  tlb_hitsVec_6; // @[TLB.scala 211:44:freechips.rocketchip.system.DefaultRV32Config.fir@177494.4]
  wire  tlb__GEN_29; // @[TLB.scala 100:18:freechips.rocketchip.system.DefaultRV32Config.fir@177499.4]
  wire  tlb__GEN_30; // @[TLB.scala 100:18:freechips.rocketchip.system.DefaultRV32Config.fir@177499.4]
  wire  tlb__GEN_31; // @[TLB.scala 100:18:freechips.rocketchip.system.DefaultRV32Config.fir@177499.4]
  wire  tlb__T_549; // @[TLB.scala 100:18:freechips.rocketchip.system.DefaultRV32Config.fir@177499.4]
  wire  tlb_hitsVec_7; // @[TLB.scala 211:44:freechips.rocketchip.system.DefaultRV32Config.fir@177500.4]
  wire  tlb_hitsVec_8; // @[TLB.scala 211:44:freechips.rocketchip.system.DefaultRV32Config.fir@177515.4]
  wire  tlb_hitsVec_9; // @[TLB.scala 211:44:freechips.rocketchip.system.DefaultRV32Config.fir@177530.4]
  wire  tlb_hitsVec_10; // @[TLB.scala 211:44:freechips.rocketchip.system.DefaultRV32Config.fir@177545.4]
  wire  tlb_hitsVec_11; // @[TLB.scala 211:44:freechips.rocketchip.system.DefaultRV32Config.fir@177560.4]
  wire [9:0] tlb__T_608; // @[TLB.scala 95:46:freechips.rocketchip.system.DefaultRV32Config.fir@177563.4]
  wire  tlb__T_610; // @[TLB.scala 95:77:freechips.rocketchip.system.DefaultRV32Config.fir@177565.4]
  wire  tlb__T_612; // @[TLB.scala 95:29:freechips.rocketchip.system.DefaultRV32Config.fir@177567.4]
  wire [9:0] tlb__T_615; // @[TLB.scala 95:46:freechips.rocketchip.system.DefaultRV32Config.fir@177570.4]
  wire  tlb__T_617; // @[TLB.scala 95:77:freechips.rocketchip.system.DefaultRV32Config.fir@177572.4]
  wire  tlb__T_618; // @[TLB.scala 95:40:freechips.rocketchip.system.DefaultRV32Config.fir@177573.4]
  wire  tlb__T_619; // @[TLB.scala 95:29:freechips.rocketchip.system.DefaultRV32Config.fir@177574.4]
  wire  tlb_hitsVec_12; // @[TLB.scala 211:44:freechips.rocketchip.system.DefaultRV32Config.fir@177575.4]
  wire [5:0] tlb__T_624; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@177580.4]
  wire [12:0] tlb_real_hits; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@177587.4]
  wire  tlb__T_631; // @[TLB.scala 213:18:freechips.rocketchip.system.DefaultRV32Config.fir@177588.4]
  wire [13:0] tlb_hits; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@177589.4]
  wire [34:0] tlb__GEN_33; // @[:freechips.rocketchip.system.DefaultRV32Config.fir@177596.4]
  wire [34:0] tlb__GEN_34; // @[:freechips.rocketchip.system.DefaultRV32Config.fir@177596.4]
  wire [34:0] tlb__GEN_35; // @[:freechips.rocketchip.system.DefaultRV32Config.fir@177596.4]
  wire [34:0] tlb__GEN_37; // @[:freechips.rocketchip.system.DefaultRV32Config.fir@177639.4]
  wire [34:0] tlb__GEN_38; // @[:freechips.rocketchip.system.DefaultRV32Config.fir@177639.4]
  wire [34:0] tlb__GEN_39; // @[:freechips.rocketchip.system.DefaultRV32Config.fir@177639.4]
  wire [34:0] tlb__GEN_41; // @[:freechips.rocketchip.system.DefaultRV32Config.fir@177682.4]
  wire [34:0] tlb__GEN_42; // @[:freechips.rocketchip.system.DefaultRV32Config.fir@177682.4]
  wire [34:0] tlb__GEN_43; // @[:freechips.rocketchip.system.DefaultRV32Config.fir@177682.4]
  wire [34:0] tlb__GEN_45; // @[:freechips.rocketchip.system.DefaultRV32Config.fir@177725.4]
  wire [34:0] tlb__GEN_46; // @[:freechips.rocketchip.system.DefaultRV32Config.fir@177725.4]
  wire [34:0] tlb__GEN_47; // @[:freechips.rocketchip.system.DefaultRV32Config.fir@177725.4]
  wire [34:0] tlb__GEN_49; // @[:freechips.rocketchip.system.DefaultRV32Config.fir@177768.4]
  wire [34:0] tlb__GEN_50; // @[:freechips.rocketchip.system.DefaultRV32Config.fir@177768.4]
  wire [34:0] tlb__GEN_51; // @[:freechips.rocketchip.system.DefaultRV32Config.fir@177768.4]
  wire [34:0] tlb__GEN_53; // @[:freechips.rocketchip.system.DefaultRV32Config.fir@177811.4]
  wire [34:0] tlb__GEN_54; // @[:freechips.rocketchip.system.DefaultRV32Config.fir@177811.4]
  wire [34:0] tlb__GEN_55; // @[:freechips.rocketchip.system.DefaultRV32Config.fir@177811.4]
  wire [34:0] tlb__GEN_57; // @[:freechips.rocketchip.system.DefaultRV32Config.fir@177854.4]
  wire [34:0] tlb__GEN_58; // @[:freechips.rocketchip.system.DefaultRV32Config.fir@177854.4]
  wire [34:0] tlb__GEN_59; // @[:freechips.rocketchip.system.DefaultRV32Config.fir@177854.4]
  wire [34:0] tlb__GEN_61; // @[:freechips.rocketchip.system.DefaultRV32Config.fir@177897.4]
  wire [34:0] tlb__GEN_62; // @[:freechips.rocketchip.system.DefaultRV32Config.fir@177897.4]
  wire [34:0] tlb__GEN_63; // @[:freechips.rocketchip.system.DefaultRV32Config.fir@177897.4]
  wire  tlb__T_800; // @[TLB.scala 86:77:freechips.rocketchip.system.DefaultRV32Config.fir@177966.4]
  wire [9:0] tlb__T_803; // @[TLB.scala 106:26:freechips.rocketchip.system.DefaultRV32Config.fir@177977.4]
  wire [19:0] tlb__T_807; // @[TLB.scala 109:47:freechips.rocketchip.system.DefaultRV32Config.fir@177981.4]
  wire [9:0] tlb__T_808; // @[TLB.scala 109:58:freechips.rocketchip.system.DefaultRV32Config.fir@177982.4]
  wire [19:0] tlb__T_809; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@177983.4]
  wire  tlb__T_825; // @[TLB.scala 86:77:freechips.rocketchip.system.DefaultRV32Config.fir@178015.4]
  wire [9:0] tlb__T_828; // @[TLB.scala 106:26:freechips.rocketchip.system.DefaultRV32Config.fir@178026.4]
  wire [19:0] tlb__T_832; // @[TLB.scala 109:47:freechips.rocketchip.system.DefaultRV32Config.fir@178030.4]
  wire [9:0] tlb__T_833; // @[TLB.scala 109:58:freechips.rocketchip.system.DefaultRV32Config.fir@178031.4]
  wire [19:0] tlb__T_834; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@178032.4]
  wire  tlb__T_850; // @[TLB.scala 86:77:freechips.rocketchip.system.DefaultRV32Config.fir@178064.4]
  wire [9:0] tlb__T_853; // @[TLB.scala 106:26:freechips.rocketchip.system.DefaultRV32Config.fir@178075.4]
  wire [19:0] tlb__T_857; // @[TLB.scala 109:47:freechips.rocketchip.system.DefaultRV32Config.fir@178079.4]
  wire [9:0] tlb__T_858; // @[TLB.scala 109:58:freechips.rocketchip.system.DefaultRV32Config.fir@178080.4]
  wire [19:0] tlb__T_859; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@178081.4]
  wire  tlb__T_875; // @[TLB.scala 86:77:freechips.rocketchip.system.DefaultRV32Config.fir@178113.4]
  wire [9:0] tlb__T_878; // @[TLB.scala 106:26:freechips.rocketchip.system.DefaultRV32Config.fir@178124.4]
  wire [19:0] tlb__T_882; // @[TLB.scala 109:47:freechips.rocketchip.system.DefaultRV32Config.fir@178128.4]
  wire [9:0] tlb__T_883; // @[TLB.scala 109:58:freechips.rocketchip.system.DefaultRV32Config.fir@178129.4]
  wire [19:0] tlb__T_884; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@178130.4]
  wire [9:0] tlb__T_903; // @[TLB.scala 106:26:freechips.rocketchip.system.DefaultRV32Config.fir@178173.4]
  wire [19:0] tlb__T_907; // @[TLB.scala 109:47:freechips.rocketchip.system.DefaultRV32Config.fir@178177.4]
  wire [9:0] tlb__T_908; // @[TLB.scala 109:58:freechips.rocketchip.system.DefaultRV32Config.fir@178178.4]
  wire [19:0] tlb__T_909; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@178179.4]
  wire [19:0] tlb__T_911; // @[Mux.scala 27:72:freechips.rocketchip.system.DefaultRV32Config.fir@178181.4]
  wire [19:0] tlb__T_912; // @[Mux.scala 27:72:freechips.rocketchip.system.DefaultRV32Config.fir@178182.4]
  wire [19:0] tlb__T_913; // @[Mux.scala 27:72:freechips.rocketchip.system.DefaultRV32Config.fir@178183.4]
  wire [19:0] tlb__T_914; // @[Mux.scala 27:72:freechips.rocketchip.system.DefaultRV32Config.fir@178184.4]
  wire [19:0] tlb__T_915; // @[Mux.scala 27:72:freechips.rocketchip.system.DefaultRV32Config.fir@178185.4]
  wire [19:0] tlb__T_916; // @[Mux.scala 27:72:freechips.rocketchip.system.DefaultRV32Config.fir@178186.4]
  wire [19:0] tlb__T_917; // @[Mux.scala 27:72:freechips.rocketchip.system.DefaultRV32Config.fir@178187.4]
  wire [19:0] tlb__T_918; // @[Mux.scala 27:72:freechips.rocketchip.system.DefaultRV32Config.fir@178188.4]
  wire [19:0] tlb__T_919; // @[Mux.scala 27:72:freechips.rocketchip.system.DefaultRV32Config.fir@178189.4]
  wire [19:0] tlb__T_920; // @[Mux.scala 27:72:freechips.rocketchip.system.DefaultRV32Config.fir@178190.4]
  wire [19:0] tlb__T_921; // @[Mux.scala 27:72:freechips.rocketchip.system.DefaultRV32Config.fir@178191.4]
  wire [19:0] tlb__T_922; // @[Mux.scala 27:72:freechips.rocketchip.system.DefaultRV32Config.fir@178192.4]
  wire [19:0] tlb__T_923; // @[Mux.scala 27:72:freechips.rocketchip.system.DefaultRV32Config.fir@178193.4]
  wire [19:0] tlb__T_924; // @[Mux.scala 27:72:freechips.rocketchip.system.DefaultRV32Config.fir@178194.4]
  wire [19:0] tlb__T_925; // @[Mux.scala 27:72:freechips.rocketchip.system.DefaultRV32Config.fir@178195.4]
  wire [19:0] tlb__T_926; // @[Mux.scala 27:72:freechips.rocketchip.system.DefaultRV32Config.fir@178196.4]
  wire [19:0] tlb__T_927; // @[Mux.scala 27:72:freechips.rocketchip.system.DefaultRV32Config.fir@178197.4]
  wire [19:0] tlb__T_928; // @[Mux.scala 27:72:freechips.rocketchip.system.DefaultRV32Config.fir@178198.4]
  wire [19:0] tlb__T_929; // @[Mux.scala 27:72:freechips.rocketchip.system.DefaultRV32Config.fir@178199.4]
  wire [19:0] tlb__T_930; // @[Mux.scala 27:72:freechips.rocketchip.system.DefaultRV32Config.fir@178200.4]
  wire [19:0] tlb__T_931; // @[Mux.scala 27:72:freechips.rocketchip.system.DefaultRV32Config.fir@178201.4]
  wire [19:0] tlb__T_932; // @[Mux.scala 27:72:freechips.rocketchip.system.DefaultRV32Config.fir@178202.4]
  wire [19:0] tlb__T_933; // @[Mux.scala 27:72:freechips.rocketchip.system.DefaultRV32Config.fir@178203.4]
  wire [19:0] tlb__T_934; // @[Mux.scala 27:72:freechips.rocketchip.system.DefaultRV32Config.fir@178204.4]
  wire [19:0] tlb__T_935; // @[Mux.scala 27:72:freechips.rocketchip.system.DefaultRV32Config.fir@178205.4]
  wire [19:0] tlb__T_936; // @[Mux.scala 27:72:freechips.rocketchip.system.DefaultRV32Config.fir@178206.4]
  wire [19:0] tlb__T_937; // @[Mux.scala 27:72:freechips.rocketchip.system.DefaultRV32Config.fir@178207.4]
  wire  tlb__T_938; // @[TLB.scala 217:22:freechips.rocketchip.system.DefaultRV32Config.fir@178210.4]
  wire  tlb__T_939; // @[TLB.scala 217:19:freechips.rocketchip.system.DefaultRV32Config.fir@178211.4]
  wire  tlb__T_941; // @[TLB.scala 223:25:freechips.rocketchip.system.DefaultRV32Config.fir@178218.6]
  wire  tlb__T_942; // @[PTW.scala 69:47:freechips.rocketchip.system.DefaultRV32Config.fir@178221.6]
  wire  tlb__T_943; // @[PTW.scala 69:44:freechips.rocketchip.system.DefaultRV32Config.fir@178222.6]
  wire  tlb__T_944; // @[PTW.scala 69:38:freechips.rocketchip.system.DefaultRV32Config.fir@178223.6]
  wire  tlb__T_945; // @[PTW.scala 69:32:freechips.rocketchip.system.DefaultRV32Config.fir@178224.6]
  wire  tlb__T_946; // @[PTW.scala 69:52:freechips.rocketchip.system.DefaultRV32Config.fir@178225.6]
  wire  tlb__T_947; // @[PTW.scala 73:35:freechips.rocketchip.system.DefaultRV32Config.fir@178226.6]
  wire  tlb__T_953; // @[PTW.scala 74:35:freechips.rocketchip.system.DefaultRV32Config.fir@178233.6]
  wire  tlb__T_954; // @[PTW.scala 74:40:freechips.rocketchip.system.DefaultRV32Config.fir@178234.6]
  wire  tlb__T_960; // @[PTW.scala 75:35:freechips.rocketchip.system.DefaultRV32Config.fir@178241.6]
  wire  tlb__T_961; // @[TLB.scala 237:37:freechips.rocketchip.system.DefaultRV32Config.fir@178251.6]
  wire [7:0] tlb__T_970; // @[TLB.scala 123:24:freechips.rocketchip.system.DefaultRV32Config.fir@178264.8]
  wire [34:0] tlb__T_978; // @[TLB.scala 123:24:freechips.rocketchip.system.DefaultRV32Config.fir@178272.8]
  wire  tlb__T_979; // @[TLB.scala 239:40:freechips.rocketchip.system.DefaultRV32Config.fir@178276.8]
  wire  tlb__T_980; // @[TLB.scala 240:82:freechips.rocketchip.system.DefaultRV32Config.fir@178278.10]
  wire  tlb__GEN_66; // @[TLB.scala 240:89:freechips.rocketchip.system.DefaultRV32Config.fir@178279.10]
  wire  tlb__T_996; // @[TLB.scala 240:82:freechips.rocketchip.system.DefaultRV32Config.fir@178300.10]
  wire  tlb__GEN_70; // @[TLB.scala 240:89:freechips.rocketchip.system.DefaultRV32Config.fir@178301.10]
  wire  tlb__T_1012; // @[TLB.scala 240:82:freechips.rocketchip.system.DefaultRV32Config.fir@178322.10]
  wire  tlb__GEN_74; // @[TLB.scala 240:89:freechips.rocketchip.system.DefaultRV32Config.fir@178323.10]
  wire  tlb__T_1028; // @[TLB.scala 240:82:freechips.rocketchip.system.DefaultRV32Config.fir@178344.10]
  wire  tlb__GEN_78; // @[TLB.scala 240:89:freechips.rocketchip.system.DefaultRV32Config.fir@178345.10]
  wire [2:0] tlb__T_1044; // @[TLB.scala 244:22:freechips.rocketchip.system.DefaultRV32Config.fir@178368.10]
  wire  tlb__T_1045; // @[TLB.scala 245:65:freechips.rocketchip.system.DefaultRV32Config.fir@178369.10]
  wire  tlb__T_1046; // @[TLB.scala 246:15:freechips.rocketchip.system.DefaultRV32Config.fir@178371.12]
  wire  tlb__GEN_80; // @[TLB.scala 246:32:freechips.rocketchip.system.DefaultRV32Config.fir@178372.12]
  wire  tlb__GEN_81; // @[TLB.scala 246:32:freechips.rocketchip.system.DefaultRV32Config.fir@178372.12]
  wire  tlb__GEN_82; // @[TLB.scala 246:32:freechips.rocketchip.system.DefaultRV32Config.fir@178372.12]
  wire  tlb__GEN_83; // @[TLB.scala 246:32:freechips.rocketchip.system.DefaultRV32Config.fir@178372.12]
  wire [1:0] tlb__T_1047; // @[package.scala 138:13:freechips.rocketchip.system.DefaultRV32Config.fir@178380.12]
  wire  _GEN_343; // @[TLB.scala 122:16:freechips.rocketchip.system.DefaultRV32Config.fir@178381.12]
  wire  tlb__GEN_84; // @[TLB.scala 122:16:freechips.rocketchip.system.DefaultRV32Config.fir@178381.12]
  wire  _GEN_344; // @[TLB.scala 122:16:freechips.rocketchip.system.DefaultRV32Config.fir@178381.12]
  wire  tlb__GEN_85; // @[TLB.scala 122:16:freechips.rocketchip.system.DefaultRV32Config.fir@178381.12]
  wire  _GEN_345; // @[TLB.scala 122:16:freechips.rocketchip.system.DefaultRV32Config.fir@178381.12]
  wire  tlb__GEN_86; // @[TLB.scala 122:16:freechips.rocketchip.system.DefaultRV32Config.fir@178381.12]
  wire  _GEN_346; // @[TLB.scala 122:16:freechips.rocketchip.system.DefaultRV32Config.fir@178381.12]
  wire  tlb__GEN_87; // @[TLB.scala 122:16:freechips.rocketchip.system.DefaultRV32Config.fir@178381.12]
  wire  tlb__GEN_92; // @[TLB.scala 245:72:freechips.rocketchip.system.DefaultRV32Config.fir@178370.10]
  wire  tlb__GEN_93; // @[TLB.scala 245:72:freechips.rocketchip.system.DefaultRV32Config.fir@178370.10]
  wire  tlb__GEN_94; // @[TLB.scala 245:72:freechips.rocketchip.system.DefaultRV32Config.fir@178370.10]
  wire  tlb__GEN_95; // @[TLB.scala 245:72:freechips.rocketchip.system.DefaultRV32Config.fir@178370.10]
  wire  tlb__T_1063; // @[TLB.scala 245:65:freechips.rocketchip.system.DefaultRV32Config.fir@178399.10]
  wire  tlb__GEN_102; // @[TLB.scala 246:32:freechips.rocketchip.system.DefaultRV32Config.fir@178402.12]
  wire  tlb__GEN_103; // @[TLB.scala 246:32:freechips.rocketchip.system.DefaultRV32Config.fir@178402.12]
  wire  tlb__GEN_104; // @[TLB.scala 246:32:freechips.rocketchip.system.DefaultRV32Config.fir@178402.12]
  wire  tlb__GEN_105; // @[TLB.scala 246:32:freechips.rocketchip.system.DefaultRV32Config.fir@178402.12]
  wire  tlb__GEN_106; // @[TLB.scala 122:16:freechips.rocketchip.system.DefaultRV32Config.fir@178411.12]
  wire  tlb__GEN_107; // @[TLB.scala 122:16:freechips.rocketchip.system.DefaultRV32Config.fir@178411.12]
  wire  tlb__GEN_108; // @[TLB.scala 122:16:freechips.rocketchip.system.DefaultRV32Config.fir@178411.12]
  wire  tlb__GEN_109; // @[TLB.scala 122:16:freechips.rocketchip.system.DefaultRV32Config.fir@178411.12]
  wire  tlb__GEN_114; // @[TLB.scala 245:72:freechips.rocketchip.system.DefaultRV32Config.fir@178400.10]
  wire  tlb__GEN_115; // @[TLB.scala 245:72:freechips.rocketchip.system.DefaultRV32Config.fir@178400.10]
  wire  tlb__GEN_116; // @[TLB.scala 245:72:freechips.rocketchip.system.DefaultRV32Config.fir@178400.10]
  wire  tlb__GEN_117; // @[TLB.scala 245:72:freechips.rocketchip.system.DefaultRV32Config.fir@178400.10]
  wire  tlb__T_1081; // @[TLB.scala 245:65:freechips.rocketchip.system.DefaultRV32Config.fir@178429.10]
  wire  tlb__GEN_124; // @[TLB.scala 246:32:freechips.rocketchip.system.DefaultRV32Config.fir@178432.12]
  wire  tlb__GEN_125; // @[TLB.scala 246:32:freechips.rocketchip.system.DefaultRV32Config.fir@178432.12]
  wire  tlb__GEN_126; // @[TLB.scala 246:32:freechips.rocketchip.system.DefaultRV32Config.fir@178432.12]
  wire  tlb__GEN_127; // @[TLB.scala 246:32:freechips.rocketchip.system.DefaultRV32Config.fir@178432.12]
  wire  tlb__GEN_128; // @[TLB.scala 122:16:freechips.rocketchip.system.DefaultRV32Config.fir@178441.12]
  wire  tlb__GEN_129; // @[TLB.scala 122:16:freechips.rocketchip.system.DefaultRV32Config.fir@178441.12]
  wire  tlb__GEN_130; // @[TLB.scala 122:16:freechips.rocketchip.system.DefaultRV32Config.fir@178441.12]
  wire  tlb__GEN_131; // @[TLB.scala 122:16:freechips.rocketchip.system.DefaultRV32Config.fir@178441.12]
  wire  tlb__GEN_136; // @[TLB.scala 245:72:freechips.rocketchip.system.DefaultRV32Config.fir@178430.10]
  wire  tlb__GEN_137; // @[TLB.scala 245:72:freechips.rocketchip.system.DefaultRV32Config.fir@178430.10]
  wire  tlb__GEN_138; // @[TLB.scala 245:72:freechips.rocketchip.system.DefaultRV32Config.fir@178430.10]
  wire  tlb__GEN_139; // @[TLB.scala 245:72:freechips.rocketchip.system.DefaultRV32Config.fir@178430.10]
  wire  tlb__T_1099; // @[TLB.scala 245:65:freechips.rocketchip.system.DefaultRV32Config.fir@178459.10]
  wire  tlb__GEN_146; // @[TLB.scala 246:32:freechips.rocketchip.system.DefaultRV32Config.fir@178462.12]
  wire  tlb__GEN_147; // @[TLB.scala 246:32:freechips.rocketchip.system.DefaultRV32Config.fir@178462.12]
  wire  tlb__GEN_148; // @[TLB.scala 246:32:freechips.rocketchip.system.DefaultRV32Config.fir@178462.12]
  wire  tlb__GEN_149; // @[TLB.scala 246:32:freechips.rocketchip.system.DefaultRV32Config.fir@178462.12]
  wire  tlb__GEN_150; // @[TLB.scala 122:16:freechips.rocketchip.system.DefaultRV32Config.fir@178471.12]
  wire  tlb__GEN_151; // @[TLB.scala 122:16:freechips.rocketchip.system.DefaultRV32Config.fir@178471.12]
  wire  tlb__GEN_152; // @[TLB.scala 122:16:freechips.rocketchip.system.DefaultRV32Config.fir@178471.12]
  wire  tlb__GEN_153; // @[TLB.scala 122:16:freechips.rocketchip.system.DefaultRV32Config.fir@178471.12]
  wire  tlb__GEN_158; // @[TLB.scala 245:72:freechips.rocketchip.system.DefaultRV32Config.fir@178460.10]
  wire  tlb__GEN_159; // @[TLB.scala 245:72:freechips.rocketchip.system.DefaultRV32Config.fir@178460.10]
  wire  tlb__GEN_160; // @[TLB.scala 245:72:freechips.rocketchip.system.DefaultRV32Config.fir@178460.10]
  wire  tlb__GEN_161; // @[TLB.scala 245:72:freechips.rocketchip.system.DefaultRV32Config.fir@178460.10]
  wire  tlb__T_1117; // @[TLB.scala 245:65:freechips.rocketchip.system.DefaultRV32Config.fir@178489.10]
  wire  tlb__GEN_168; // @[TLB.scala 246:32:freechips.rocketchip.system.DefaultRV32Config.fir@178492.12]
  wire  tlb__GEN_169; // @[TLB.scala 246:32:freechips.rocketchip.system.DefaultRV32Config.fir@178492.12]
  wire  tlb__GEN_170; // @[TLB.scala 246:32:freechips.rocketchip.system.DefaultRV32Config.fir@178492.12]
  wire  tlb__GEN_171; // @[TLB.scala 246:32:freechips.rocketchip.system.DefaultRV32Config.fir@178492.12]
  wire  tlb__GEN_172; // @[TLB.scala 122:16:freechips.rocketchip.system.DefaultRV32Config.fir@178501.12]
  wire  tlb__GEN_173; // @[TLB.scala 122:16:freechips.rocketchip.system.DefaultRV32Config.fir@178501.12]
  wire  tlb__GEN_174; // @[TLB.scala 122:16:freechips.rocketchip.system.DefaultRV32Config.fir@178501.12]
  wire  tlb__GEN_175; // @[TLB.scala 122:16:freechips.rocketchip.system.DefaultRV32Config.fir@178501.12]
  wire  tlb__GEN_180; // @[TLB.scala 245:72:freechips.rocketchip.system.DefaultRV32Config.fir@178490.10]
  wire  tlb__GEN_181; // @[TLB.scala 245:72:freechips.rocketchip.system.DefaultRV32Config.fir@178490.10]
  wire  tlb__GEN_182; // @[TLB.scala 245:72:freechips.rocketchip.system.DefaultRV32Config.fir@178490.10]
  wire  tlb__GEN_183; // @[TLB.scala 245:72:freechips.rocketchip.system.DefaultRV32Config.fir@178490.10]
  wire  tlb__T_1135; // @[TLB.scala 245:65:freechips.rocketchip.system.DefaultRV32Config.fir@178519.10]
  wire  tlb__GEN_190; // @[TLB.scala 246:32:freechips.rocketchip.system.DefaultRV32Config.fir@178522.12]
  wire  tlb__GEN_191; // @[TLB.scala 246:32:freechips.rocketchip.system.DefaultRV32Config.fir@178522.12]
  wire  tlb__GEN_192; // @[TLB.scala 246:32:freechips.rocketchip.system.DefaultRV32Config.fir@178522.12]
  wire  tlb__GEN_193; // @[TLB.scala 246:32:freechips.rocketchip.system.DefaultRV32Config.fir@178522.12]
  wire  tlb__GEN_194; // @[TLB.scala 122:16:freechips.rocketchip.system.DefaultRV32Config.fir@178531.12]
  wire  tlb__GEN_195; // @[TLB.scala 122:16:freechips.rocketchip.system.DefaultRV32Config.fir@178531.12]
  wire  tlb__GEN_196; // @[TLB.scala 122:16:freechips.rocketchip.system.DefaultRV32Config.fir@178531.12]
  wire  tlb__GEN_197; // @[TLB.scala 122:16:freechips.rocketchip.system.DefaultRV32Config.fir@178531.12]
  wire  tlb__GEN_202; // @[TLB.scala 245:72:freechips.rocketchip.system.DefaultRV32Config.fir@178520.10]
  wire  tlb__GEN_203; // @[TLB.scala 245:72:freechips.rocketchip.system.DefaultRV32Config.fir@178520.10]
  wire  tlb__GEN_204; // @[TLB.scala 245:72:freechips.rocketchip.system.DefaultRV32Config.fir@178520.10]
  wire  tlb__GEN_205; // @[TLB.scala 245:72:freechips.rocketchip.system.DefaultRV32Config.fir@178520.10]
  wire  tlb__T_1153; // @[TLB.scala 245:65:freechips.rocketchip.system.DefaultRV32Config.fir@178549.10]
  wire  tlb__GEN_212; // @[TLB.scala 246:32:freechips.rocketchip.system.DefaultRV32Config.fir@178552.12]
  wire  tlb__GEN_213; // @[TLB.scala 246:32:freechips.rocketchip.system.DefaultRV32Config.fir@178552.12]
  wire  tlb__GEN_214; // @[TLB.scala 246:32:freechips.rocketchip.system.DefaultRV32Config.fir@178552.12]
  wire  tlb__GEN_215; // @[TLB.scala 246:32:freechips.rocketchip.system.DefaultRV32Config.fir@178552.12]
  wire  tlb__GEN_216; // @[TLB.scala 122:16:freechips.rocketchip.system.DefaultRV32Config.fir@178561.12]
  wire  tlb__GEN_217; // @[TLB.scala 122:16:freechips.rocketchip.system.DefaultRV32Config.fir@178561.12]
  wire  tlb__GEN_218; // @[TLB.scala 122:16:freechips.rocketchip.system.DefaultRV32Config.fir@178561.12]
  wire  tlb__GEN_219; // @[TLB.scala 122:16:freechips.rocketchip.system.DefaultRV32Config.fir@178561.12]
  wire  tlb__GEN_224; // @[TLB.scala 245:72:freechips.rocketchip.system.DefaultRV32Config.fir@178550.10]
  wire  tlb__GEN_225; // @[TLB.scala 245:72:freechips.rocketchip.system.DefaultRV32Config.fir@178550.10]
  wire  tlb__GEN_226; // @[TLB.scala 245:72:freechips.rocketchip.system.DefaultRV32Config.fir@178550.10]
  wire  tlb__GEN_227; // @[TLB.scala 245:72:freechips.rocketchip.system.DefaultRV32Config.fir@178550.10]
  wire  tlb__T_1171; // @[TLB.scala 245:65:freechips.rocketchip.system.DefaultRV32Config.fir@178579.10]
  wire  tlb__GEN_234; // @[TLB.scala 246:32:freechips.rocketchip.system.DefaultRV32Config.fir@178582.12]
  wire  tlb__GEN_235; // @[TLB.scala 246:32:freechips.rocketchip.system.DefaultRV32Config.fir@178582.12]
  wire  tlb__GEN_236; // @[TLB.scala 246:32:freechips.rocketchip.system.DefaultRV32Config.fir@178582.12]
  wire  tlb__GEN_237; // @[TLB.scala 246:32:freechips.rocketchip.system.DefaultRV32Config.fir@178582.12]
  wire  tlb__GEN_238; // @[TLB.scala 122:16:freechips.rocketchip.system.DefaultRV32Config.fir@178591.12]
  wire  tlb__GEN_239; // @[TLB.scala 122:16:freechips.rocketchip.system.DefaultRV32Config.fir@178591.12]
  wire  tlb__GEN_240; // @[TLB.scala 122:16:freechips.rocketchip.system.DefaultRV32Config.fir@178591.12]
  wire  tlb__GEN_241; // @[TLB.scala 122:16:freechips.rocketchip.system.DefaultRV32Config.fir@178591.12]
  wire  tlb__GEN_246; // @[TLB.scala 245:72:freechips.rocketchip.system.DefaultRV32Config.fir@178580.10]
  wire  tlb__GEN_247; // @[TLB.scala 245:72:freechips.rocketchip.system.DefaultRV32Config.fir@178580.10]
  wire  tlb__GEN_248; // @[TLB.scala 245:72:freechips.rocketchip.system.DefaultRV32Config.fir@178580.10]
  wire  tlb__GEN_249; // @[TLB.scala 245:72:freechips.rocketchip.system.DefaultRV32Config.fir@178580.10]
  wire  tlb__GEN_258; // @[TLB.scala 239:54:freechips.rocketchip.system.DefaultRV32Config.fir@178277.8]
  wire  tlb__GEN_262; // @[TLB.scala 239:54:freechips.rocketchip.system.DefaultRV32Config.fir@178277.8]
  wire  tlb__GEN_266; // @[TLB.scala 239:54:freechips.rocketchip.system.DefaultRV32Config.fir@178277.8]
  wire  tlb__GEN_270; // @[TLB.scala 239:54:freechips.rocketchip.system.DefaultRV32Config.fir@178277.8]
  wire  tlb__GEN_272; // @[TLB.scala 239:54:freechips.rocketchip.system.DefaultRV32Config.fir@178277.8]
  wire  tlb__GEN_273; // @[TLB.scala 239:54:freechips.rocketchip.system.DefaultRV32Config.fir@178277.8]
  wire  tlb__GEN_274; // @[TLB.scala 239:54:freechips.rocketchip.system.DefaultRV32Config.fir@178277.8]
  wire  tlb__GEN_275; // @[TLB.scala 239:54:freechips.rocketchip.system.DefaultRV32Config.fir@178277.8]
  wire  tlb__GEN_282; // @[TLB.scala 239:54:freechips.rocketchip.system.DefaultRV32Config.fir@178277.8]
  wire  tlb__GEN_283; // @[TLB.scala 239:54:freechips.rocketchip.system.DefaultRV32Config.fir@178277.8]
  wire  tlb__GEN_284; // @[TLB.scala 239:54:freechips.rocketchip.system.DefaultRV32Config.fir@178277.8]
  wire  tlb__GEN_285; // @[TLB.scala 239:54:freechips.rocketchip.system.DefaultRV32Config.fir@178277.8]
  wire  tlb__GEN_292; // @[TLB.scala 239:54:freechips.rocketchip.system.DefaultRV32Config.fir@178277.8]
  wire  tlb__GEN_293; // @[TLB.scala 239:54:freechips.rocketchip.system.DefaultRV32Config.fir@178277.8]
  wire  tlb__GEN_294; // @[TLB.scala 239:54:freechips.rocketchip.system.DefaultRV32Config.fir@178277.8]
  wire  tlb__GEN_295; // @[TLB.scala 239:54:freechips.rocketchip.system.DefaultRV32Config.fir@178277.8]
  wire  tlb__GEN_302; // @[TLB.scala 239:54:freechips.rocketchip.system.DefaultRV32Config.fir@178277.8]
  wire  tlb__GEN_303; // @[TLB.scala 239:54:freechips.rocketchip.system.DefaultRV32Config.fir@178277.8]
  wire  tlb__GEN_304; // @[TLB.scala 239:54:freechips.rocketchip.system.DefaultRV32Config.fir@178277.8]
  wire  tlb__GEN_305; // @[TLB.scala 239:54:freechips.rocketchip.system.DefaultRV32Config.fir@178277.8]
  wire  tlb__GEN_312; // @[TLB.scala 239:54:freechips.rocketchip.system.DefaultRV32Config.fir@178277.8]
  wire  tlb__GEN_313; // @[TLB.scala 239:54:freechips.rocketchip.system.DefaultRV32Config.fir@178277.8]
  wire  tlb__GEN_314; // @[TLB.scala 239:54:freechips.rocketchip.system.DefaultRV32Config.fir@178277.8]
  wire  tlb__GEN_315; // @[TLB.scala 239:54:freechips.rocketchip.system.DefaultRV32Config.fir@178277.8]
  wire  tlb__GEN_322; // @[TLB.scala 239:54:freechips.rocketchip.system.DefaultRV32Config.fir@178277.8]
  wire  tlb__GEN_323; // @[TLB.scala 239:54:freechips.rocketchip.system.DefaultRV32Config.fir@178277.8]
  wire  tlb__GEN_324; // @[TLB.scala 239:54:freechips.rocketchip.system.DefaultRV32Config.fir@178277.8]
  wire  tlb__GEN_325; // @[TLB.scala 239:54:freechips.rocketchip.system.DefaultRV32Config.fir@178277.8]
  wire  tlb__GEN_332; // @[TLB.scala 239:54:freechips.rocketchip.system.DefaultRV32Config.fir@178277.8]
  wire  tlb__GEN_333; // @[TLB.scala 239:54:freechips.rocketchip.system.DefaultRV32Config.fir@178277.8]
  wire  tlb__GEN_334; // @[TLB.scala 239:54:freechips.rocketchip.system.DefaultRV32Config.fir@178277.8]
  wire  tlb__GEN_335; // @[TLB.scala 239:54:freechips.rocketchip.system.DefaultRV32Config.fir@178277.8]
  wire  tlb__GEN_342; // @[TLB.scala 239:54:freechips.rocketchip.system.DefaultRV32Config.fir@178277.8]
  wire  tlb__GEN_343; // @[TLB.scala 239:54:freechips.rocketchip.system.DefaultRV32Config.fir@178277.8]
  wire  tlb__GEN_344; // @[TLB.scala 239:54:freechips.rocketchip.system.DefaultRV32Config.fir@178277.8]
  wire  tlb__GEN_345; // @[TLB.scala 239:54:freechips.rocketchip.system.DefaultRV32Config.fir@178277.8]
  wire  tlb__GEN_354; // @[TLB.scala 237:68:freechips.rocketchip.system.DefaultRV32Config.fir@178253.6]
  wire  tlb__GEN_358; // @[TLB.scala 237:68:freechips.rocketchip.system.DefaultRV32Config.fir@178253.6]
  wire  tlb__GEN_362; // @[TLB.scala 237:68:freechips.rocketchip.system.DefaultRV32Config.fir@178253.6]
  wire  tlb__GEN_366; // @[TLB.scala 237:68:freechips.rocketchip.system.DefaultRV32Config.fir@178253.6]
  wire  tlb__GEN_370; // @[TLB.scala 237:68:freechips.rocketchip.system.DefaultRV32Config.fir@178253.6]
  wire  tlb__GEN_372; // @[TLB.scala 237:68:freechips.rocketchip.system.DefaultRV32Config.fir@178253.6]
  wire  tlb__GEN_373; // @[TLB.scala 237:68:freechips.rocketchip.system.DefaultRV32Config.fir@178253.6]
  wire  tlb__GEN_374; // @[TLB.scala 237:68:freechips.rocketchip.system.DefaultRV32Config.fir@178253.6]
  wire  tlb__GEN_375; // @[TLB.scala 237:68:freechips.rocketchip.system.DefaultRV32Config.fir@178253.6]
  wire  tlb__GEN_382; // @[TLB.scala 237:68:freechips.rocketchip.system.DefaultRV32Config.fir@178253.6]
  wire  tlb__GEN_383; // @[TLB.scala 237:68:freechips.rocketchip.system.DefaultRV32Config.fir@178253.6]
  wire  tlb__GEN_384; // @[TLB.scala 237:68:freechips.rocketchip.system.DefaultRV32Config.fir@178253.6]
  wire  tlb__GEN_385; // @[TLB.scala 237:68:freechips.rocketchip.system.DefaultRV32Config.fir@178253.6]
  wire  tlb__GEN_392; // @[TLB.scala 237:68:freechips.rocketchip.system.DefaultRV32Config.fir@178253.6]
  wire  tlb__GEN_393; // @[TLB.scala 237:68:freechips.rocketchip.system.DefaultRV32Config.fir@178253.6]
  wire  tlb__GEN_394; // @[TLB.scala 237:68:freechips.rocketchip.system.DefaultRV32Config.fir@178253.6]
  wire  tlb__GEN_395; // @[TLB.scala 237:68:freechips.rocketchip.system.DefaultRV32Config.fir@178253.6]
  wire  tlb__GEN_402; // @[TLB.scala 237:68:freechips.rocketchip.system.DefaultRV32Config.fir@178253.6]
  wire  tlb__GEN_403; // @[TLB.scala 237:68:freechips.rocketchip.system.DefaultRV32Config.fir@178253.6]
  wire  tlb__GEN_404; // @[TLB.scala 237:68:freechips.rocketchip.system.DefaultRV32Config.fir@178253.6]
  wire  tlb__GEN_405; // @[TLB.scala 237:68:freechips.rocketchip.system.DefaultRV32Config.fir@178253.6]
  wire  tlb__GEN_412; // @[TLB.scala 237:68:freechips.rocketchip.system.DefaultRV32Config.fir@178253.6]
  wire  tlb__GEN_413; // @[TLB.scala 237:68:freechips.rocketchip.system.DefaultRV32Config.fir@178253.6]
  wire  tlb__GEN_414; // @[TLB.scala 237:68:freechips.rocketchip.system.DefaultRV32Config.fir@178253.6]
  wire  tlb__GEN_415; // @[TLB.scala 237:68:freechips.rocketchip.system.DefaultRV32Config.fir@178253.6]
  wire  tlb__GEN_422; // @[TLB.scala 237:68:freechips.rocketchip.system.DefaultRV32Config.fir@178253.6]
  wire  tlb__GEN_423; // @[TLB.scala 237:68:freechips.rocketchip.system.DefaultRV32Config.fir@178253.6]
  wire  tlb__GEN_424; // @[TLB.scala 237:68:freechips.rocketchip.system.DefaultRV32Config.fir@178253.6]
  wire  tlb__GEN_425; // @[TLB.scala 237:68:freechips.rocketchip.system.DefaultRV32Config.fir@178253.6]
  wire  tlb__GEN_432; // @[TLB.scala 237:68:freechips.rocketchip.system.DefaultRV32Config.fir@178253.6]
  wire  tlb__GEN_433; // @[TLB.scala 237:68:freechips.rocketchip.system.DefaultRV32Config.fir@178253.6]
  wire  tlb__GEN_434; // @[TLB.scala 237:68:freechips.rocketchip.system.DefaultRV32Config.fir@178253.6]
  wire  tlb__GEN_435; // @[TLB.scala 237:68:freechips.rocketchip.system.DefaultRV32Config.fir@178253.6]
  wire  tlb__GEN_442; // @[TLB.scala 237:68:freechips.rocketchip.system.DefaultRV32Config.fir@178253.6]
  wire  tlb__GEN_443; // @[TLB.scala 237:68:freechips.rocketchip.system.DefaultRV32Config.fir@178253.6]
  wire  tlb__GEN_444; // @[TLB.scala 237:68:freechips.rocketchip.system.DefaultRV32Config.fir@178253.6]
  wire  tlb__GEN_445; // @[TLB.scala 237:68:freechips.rocketchip.system.DefaultRV32Config.fir@178253.6]
  wire  tlb__GEN_454; // @[TLB.scala 217:42:freechips.rocketchip.system.DefaultRV32Config.fir@178212.4]
  wire  tlb__GEN_458; // @[TLB.scala 217:42:freechips.rocketchip.system.DefaultRV32Config.fir@178212.4]
  wire  tlb__GEN_462; // @[TLB.scala 217:42:freechips.rocketchip.system.DefaultRV32Config.fir@178212.4]
  wire  tlb__GEN_466; // @[TLB.scala 217:42:freechips.rocketchip.system.DefaultRV32Config.fir@178212.4]
  wire  tlb__GEN_470; // @[TLB.scala 217:42:freechips.rocketchip.system.DefaultRV32Config.fir@178212.4]
  wire  tlb__GEN_472; // @[TLB.scala 217:42:freechips.rocketchip.system.DefaultRV32Config.fir@178212.4]
  wire  tlb__GEN_473; // @[TLB.scala 217:42:freechips.rocketchip.system.DefaultRV32Config.fir@178212.4]
  wire  tlb__GEN_474; // @[TLB.scala 217:42:freechips.rocketchip.system.DefaultRV32Config.fir@178212.4]
  wire  tlb__GEN_475; // @[TLB.scala 217:42:freechips.rocketchip.system.DefaultRV32Config.fir@178212.4]
  wire  tlb__GEN_482; // @[TLB.scala 217:42:freechips.rocketchip.system.DefaultRV32Config.fir@178212.4]
  wire  tlb__GEN_483; // @[TLB.scala 217:42:freechips.rocketchip.system.DefaultRV32Config.fir@178212.4]
  wire  tlb__GEN_484; // @[TLB.scala 217:42:freechips.rocketchip.system.DefaultRV32Config.fir@178212.4]
  wire  tlb__GEN_485; // @[TLB.scala 217:42:freechips.rocketchip.system.DefaultRV32Config.fir@178212.4]
  wire  tlb__GEN_492; // @[TLB.scala 217:42:freechips.rocketchip.system.DefaultRV32Config.fir@178212.4]
  wire  tlb__GEN_493; // @[TLB.scala 217:42:freechips.rocketchip.system.DefaultRV32Config.fir@178212.4]
  wire  tlb__GEN_494; // @[TLB.scala 217:42:freechips.rocketchip.system.DefaultRV32Config.fir@178212.4]
  wire  tlb__GEN_495; // @[TLB.scala 217:42:freechips.rocketchip.system.DefaultRV32Config.fir@178212.4]
  wire  tlb__GEN_502; // @[TLB.scala 217:42:freechips.rocketchip.system.DefaultRV32Config.fir@178212.4]
  wire  tlb__GEN_503; // @[TLB.scala 217:42:freechips.rocketchip.system.DefaultRV32Config.fir@178212.4]
  wire  tlb__GEN_504; // @[TLB.scala 217:42:freechips.rocketchip.system.DefaultRV32Config.fir@178212.4]
  wire  tlb__GEN_505; // @[TLB.scala 217:42:freechips.rocketchip.system.DefaultRV32Config.fir@178212.4]
  wire  tlb__GEN_512; // @[TLB.scala 217:42:freechips.rocketchip.system.DefaultRV32Config.fir@178212.4]
  wire  tlb__GEN_513; // @[TLB.scala 217:42:freechips.rocketchip.system.DefaultRV32Config.fir@178212.4]
  wire  tlb__GEN_514; // @[TLB.scala 217:42:freechips.rocketchip.system.DefaultRV32Config.fir@178212.4]
  wire  tlb__GEN_515; // @[TLB.scala 217:42:freechips.rocketchip.system.DefaultRV32Config.fir@178212.4]
  wire  tlb__GEN_522; // @[TLB.scala 217:42:freechips.rocketchip.system.DefaultRV32Config.fir@178212.4]
  wire  tlb__GEN_523; // @[TLB.scala 217:42:freechips.rocketchip.system.DefaultRV32Config.fir@178212.4]
  wire  tlb__GEN_524; // @[TLB.scala 217:42:freechips.rocketchip.system.DefaultRV32Config.fir@178212.4]
  wire  tlb__GEN_525; // @[TLB.scala 217:42:freechips.rocketchip.system.DefaultRV32Config.fir@178212.4]
  wire  tlb__GEN_532; // @[TLB.scala 217:42:freechips.rocketchip.system.DefaultRV32Config.fir@178212.4]
  wire  tlb__GEN_533; // @[TLB.scala 217:42:freechips.rocketchip.system.DefaultRV32Config.fir@178212.4]
  wire  tlb__GEN_534; // @[TLB.scala 217:42:freechips.rocketchip.system.DefaultRV32Config.fir@178212.4]
  wire  tlb__GEN_535; // @[TLB.scala 217:42:freechips.rocketchip.system.DefaultRV32Config.fir@178212.4]
  wire  tlb__GEN_542; // @[TLB.scala 217:42:freechips.rocketchip.system.DefaultRV32Config.fir@178212.4]
  wire  tlb__GEN_543; // @[TLB.scala 217:42:freechips.rocketchip.system.DefaultRV32Config.fir@178212.4]
  wire  tlb__GEN_544; // @[TLB.scala 217:42:freechips.rocketchip.system.DefaultRV32Config.fir@178212.4]
  wire  tlb__GEN_545; // @[TLB.scala 217:42:freechips.rocketchip.system.DefaultRV32Config.fir@178212.4]
  wire [5:0] tlb__T_1659; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@179681.4]
  wire [13:0] tlb_ptw_ae_array; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@179689.4]
  wire  tlb__T_1667; // @[TLB.scala 256:24:freechips.rocketchip.system.DefaultRV32Config.fir@179690.4]
  wire  tlb__T_1668; // @[TLB.scala 256:32:freechips.rocketchip.system.DefaultRV32Config.fir@179691.4]
  wire [5:0] tlb__T_1673; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@179696.4]
  wire [12:0] tlb__T_1680; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@179703.4]
  wire [12:0] tlb__T_1681; // @[TLB.scala 256:23:freechips.rocketchip.system.DefaultRV32Config.fir@179704.4]
  wire [12:0] tlb__T_1694; // @[TLB.scala 256:98:freechips.rocketchip.system.DefaultRV32Config.fir@179717.4]
  wire [12:0] tlb__T_1695; // @[TLB.scala 256:89:freechips.rocketchip.system.DefaultRV32Config.fir@179718.4]
  wire [12:0] tlb_priv_rw_ok; // @[TLB.scala 256:84:freechips.rocketchip.system.DefaultRV32Config.fir@179719.4]
  wire [5:0] tlb__T_1725; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@179750.4]
  wire [12:0] tlb__T_1732; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@179757.4]
  wire [5:0] tlb__T_1737; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@179762.4]
  wire [12:0] tlb__T_1744; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@179769.4]
  wire [12:0] tlb__T_1745; // @[TLB.scala 258:73:freechips.rocketchip.system.DefaultRV32Config.fir@179770.4]
  wire [12:0] tlb__T_1746; // @[TLB.scala 258:68:freechips.rocketchip.system.DefaultRV32Config.fir@179771.4]
  wire [12:0] tlb__T_1747; // @[TLB.scala 258:40:freechips.rocketchip.system.DefaultRV32Config.fir@179772.4]
  wire [13:0] tlb_r_array; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@179773.4]
  wire [5:0] tlb__T_1752; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@179778.4]
  wire [12:0] tlb__T_1759; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@179785.4]
  wire [12:0] tlb__T_1760; // @[TLB.scala 259:40:freechips.rocketchip.system.DefaultRV32Config.fir@179786.4]
  wire [13:0] tlb_w_array; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@179787.4]
  wire [1:0] tlb__T_1775; // @[Bitwise.scala 72:12:freechips.rocketchip.system.DefaultRV32Config.fir@179803.4]
  wire [5:0] tlb__T_1780; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@179808.4]
  wire [13:0] tlb__T_1787; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@179815.4]
  wire [13:0] tlb__T_1788; // @[TLB.scala 261:89:freechips.rocketchip.system.DefaultRV32Config.fir@179816.4]
  wire [13:0] tlb_pr_array; // @[TLB.scala 261:87:freechips.rocketchip.system.DefaultRV32Config.fir@179817.4]
  wire [1:0] tlb__T_1790; // @[Bitwise.scala 72:12:freechips.rocketchip.system.DefaultRV32Config.fir@179819.4]
  wire [5:0] tlb__T_1795; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@179824.4]
  wire [13:0] tlb__T_1802; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@179831.4]
  wire [13:0] tlb_pw_array; // @[TLB.scala 262:87:freechips.rocketchip.system.DefaultRV32Config.fir@179833.4]
  wire [1:0] tlb__T_1820; // @[Bitwise.scala 72:12:freechips.rocketchip.system.DefaultRV32Config.fir@179851.4]
  wire [5:0] tlb__T_1825; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@179856.4]
  wire [13:0] tlb_eff_array; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@179863.4]
  wire [1:0] tlb__T_1833; // @[Bitwise.scala 72:12:freechips.rocketchip.system.DefaultRV32Config.fir@179865.4]
  wire [5:0] tlb__T_1838; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@179870.4]
  wire [13:0] tlb_c_array; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@179877.4]
  wire [1:0] tlb__T_1846; // @[Bitwise.scala 72:12:freechips.rocketchip.system.DefaultRV32Config.fir@179879.4]
  wire [5:0] tlb__T_1851; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@179884.4]
  wire [13:0] tlb_ppp_array; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@179891.4]
  wire [1:0] tlb__T_1859; // @[Bitwise.scala 72:12:freechips.rocketchip.system.DefaultRV32Config.fir@179893.4]
  wire [5:0] tlb__T_1864; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@179898.4]
  wire [13:0] tlb_paa_array; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@179905.4]
  wire [5:0] tlb__T_1877; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@179912.4]
  wire [13:0] tlb_pal_array; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@179919.4]
  wire [13:0] tlb_ppp_array_if_cached; // @[TLB.scala 269:39:freechips.rocketchip.system.DefaultRV32Config.fir@179920.4]
  wire [13:0] tlb_paa_array_if_cached; // @[TLB.scala 270:39:freechips.rocketchip.system.DefaultRV32Config.fir@179922.4]
  wire [13:0] tlb_pal_array_if_cached; // @[TLB.scala 271:39:freechips.rocketchip.system.DefaultRV32Config.fir@179924.4]
  wire [3:0] tlb__T_1899; // @[OneHot.scala 58:35:freechips.rocketchip.system.DefaultRV32Config.fir@179939.4]
  wire [3:0] tlb__T_1901; // @[TLB.scala 274:69:freechips.rocketchip.system.DefaultRV32Config.fir@179941.4]
  wire [31:0] _GEN_375; // @[TLB.scala 274:39:freechips.rocketchip.system.DefaultRV32Config.fir@179942.4]
  wire [31:0] tlb__T_1902; // @[TLB.scala 274:39:freechips.rocketchip.system.DefaultRV32Config.fir@179942.4]
  wire  tlb_misaligned; // @[TLB.scala 274:75:freechips.rocketchip.system.DefaultRV32Config.fir@179943.4]
  wire  tlb__T_1903; // @[package.scala 15:47:freechips.rocketchip.system.DefaultRV32Config.fir@179944.4]
  wire  tlb__T_1904; // @[package.scala 15:47:freechips.rocketchip.system.DefaultRV32Config.fir@179945.4]
  wire  tlb__T_1905; // @[package.scala 64:59:freechips.rocketchip.system.DefaultRV32Config.fir@179946.4]
  wire  tlb__T_1906; // @[package.scala 15:47:freechips.rocketchip.system.DefaultRV32Config.fir@179948.4]
  wire  tlb__T_1907; // @[package.scala 15:47:freechips.rocketchip.system.DefaultRV32Config.fir@179949.4]
  wire  tlb__T_1908; // @[package.scala 15:47:freechips.rocketchip.system.DefaultRV32Config.fir@179950.4]
  wire  tlb__T_1909; // @[package.scala 15:47:freechips.rocketchip.system.DefaultRV32Config.fir@179951.4]
  wire  tlb__T_1910; // @[package.scala 64:59:freechips.rocketchip.system.DefaultRV32Config.fir@179952.4]
  wire  tlb__T_1911; // @[package.scala 64:59:freechips.rocketchip.system.DefaultRV32Config.fir@179953.4]
  wire  tlb__T_1912; // @[package.scala 64:59:freechips.rocketchip.system.DefaultRV32Config.fir@179954.4]
  wire  tlb__T_1913; // @[package.scala 15:47:freechips.rocketchip.system.DefaultRV32Config.fir@179956.4]
  wire  tlb__T_1914; // @[package.scala 15:47:freechips.rocketchip.system.DefaultRV32Config.fir@179957.4]
  wire  tlb__T_1915; // @[package.scala 15:47:freechips.rocketchip.system.DefaultRV32Config.fir@179958.4]
  wire  tlb__T_1916; // @[package.scala 15:47:freechips.rocketchip.system.DefaultRV32Config.fir@179959.4]
  wire  tlb__T_1917; // @[package.scala 15:47:freechips.rocketchip.system.DefaultRV32Config.fir@179960.4]
  wire  tlb__T_1918; // @[package.scala 64:59:freechips.rocketchip.system.DefaultRV32Config.fir@179961.4]
  wire  tlb__T_1919; // @[package.scala 64:59:freechips.rocketchip.system.DefaultRV32Config.fir@179962.4]
  wire  tlb__T_1920; // @[package.scala 64:59:freechips.rocketchip.system.DefaultRV32Config.fir@179963.4]
  wire  tlb__T_1921; // @[package.scala 64:59:freechips.rocketchip.system.DefaultRV32Config.fir@179964.4]
  wire  tlb_cmd_put_partial; // @[TLB.scala 288:41:freechips.rocketchip.system.DefaultRV32Config.fir@179966.4]
  wire  tlb__T_1922; // @[Consts.scala 82:31:freechips.rocketchip.system.DefaultRV32Config.fir@179967.4]
  wire  tlb__T_1924; // @[Consts.scala 82:41:freechips.rocketchip.system.DefaultRV32Config.fir@179969.4]
  wire  tlb__T_1926; // @[Consts.scala 82:58:freechips.rocketchip.system.DefaultRV32Config.fir@179971.4]
  wire  tlb__T_1943; // @[Consts.scala 80:44:freechips.rocketchip.system.DefaultRV32Config.fir@179988.4]
  wire  tlb_cmd_read; // @[Consts.scala 82:75:freechips.rocketchip.system.DefaultRV32Config.fir@179989.4]
  wire  tlb__T_1944; // @[Consts.scala 83:32:freechips.rocketchip.system.DefaultRV32Config.fir@179990.4]
  wire  tlb__T_1946; // @[Consts.scala 83:42:freechips.rocketchip.system.DefaultRV32Config.fir@179992.4]
  wire  tlb__T_1948; // @[Consts.scala 83:59:freechips.rocketchip.system.DefaultRV32Config.fir@179994.4]
  wire  tlb_cmd_write; // @[Consts.scala 83:76:freechips.rocketchip.system.DefaultRV32Config.fir@180012.4]
  wire  tlb__T_1966; // @[package.scala 15:47:freechips.rocketchip.system.DefaultRV32Config.fir@180013.4]
  wire  tlb__T_1967; // @[package.scala 15:47:freechips.rocketchip.system.DefaultRV32Config.fir@180014.4]
  wire  tlb__T_1968; // @[package.scala 64:59:freechips.rocketchip.system.DefaultRV32Config.fir@180015.4]
  wire  tlb_cmd_write_perms; // @[TLB.scala 291:35:freechips.rocketchip.system.DefaultRV32Config.fir@180016.4]
  wire [13:0] tlb__T_1969; // @[TLB.scala 296:8:freechips.rocketchip.system.DefaultRV32Config.fir@180018.4]
  wire [13:0] tlb__T_1970; // @[TLB.scala 297:19:freechips.rocketchip.system.DefaultRV32Config.fir@180019.4]
  wire [13:0] tlb__T_1971; // @[TLB.scala 297:8:freechips.rocketchip.system.DefaultRV32Config.fir@180020.4]
  wire [13:0] tlb_ae_array; // @[TLB.scala 296:37:freechips.rocketchip.system.DefaultRV32Config.fir@180021.4]
  wire [13:0] tlb__T_1972; // @[TLB.scala 298:46:freechips.rocketchip.system.DefaultRV32Config.fir@180022.4]
  wire [13:0] tlb__T_1973; // @[TLB.scala 298:44:freechips.rocketchip.system.DefaultRV32Config.fir@180023.4]
  wire [13:0] tlb_ae_ld_array; // @[TLB.scala 298:24:freechips.rocketchip.system.DefaultRV32Config.fir@180024.4]
  wire [13:0] tlb__T_1974; // @[TLB.scala 300:37:freechips.rocketchip.system.DefaultRV32Config.fir@180025.4]
  wire [13:0] tlb__T_1975; // @[TLB.scala 300:35:freechips.rocketchip.system.DefaultRV32Config.fir@180026.4]
  wire [13:0] tlb__T_1976; // @[TLB.scala 300:8:freechips.rocketchip.system.DefaultRV32Config.fir@180027.4]
  wire [13:0] tlb__T_1977; // @[TLB.scala 301:26:freechips.rocketchip.system.DefaultRV32Config.fir@180028.4]
  wire [13:0] tlb__T_1978; // @[TLB.scala 301:8:freechips.rocketchip.system.DefaultRV32Config.fir@180029.4]
  wire [13:0] tlb__T_1979; // @[TLB.scala 300:53:freechips.rocketchip.system.DefaultRV32Config.fir@180030.4]
  wire [13:0] tlb__T_1980; // @[TLB.scala 302:26:freechips.rocketchip.system.DefaultRV32Config.fir@180031.4]
  wire [13:0] tlb__T_1981; // @[TLB.scala 302:8:freechips.rocketchip.system.DefaultRV32Config.fir@180032.4]
  wire [13:0] tlb__T_1982; // @[TLB.scala 301:53:freechips.rocketchip.system.DefaultRV32Config.fir@180033.4]
  wire [13:0] tlb__T_1983; // @[TLB.scala 303:29:freechips.rocketchip.system.DefaultRV32Config.fir@180034.4]
  wire [13:0] tlb__T_1984; // @[TLB.scala 303:8:freechips.rocketchip.system.DefaultRV32Config.fir@180035.4]
  wire [13:0] tlb_ae_st_array; // @[TLB.scala 302:53:freechips.rocketchip.system.DefaultRV32Config.fir@180036.4]
  wire  tlb__T_1995; // @[TLB.scala 309:36:freechips.rocketchip.system.DefaultRV32Config.fir@180048.4]
  wire [13:0] tlb__T_1996; // @[TLB.scala 309:49:freechips.rocketchip.system.DefaultRV32Config.fir@180049.4]
  wire [13:0] tlb_ma_ld_array; // @[TLB.scala 309:24:freechips.rocketchip.system.DefaultRV32Config.fir@180050.4]
  wire  tlb__T_1997; // @[TLB.scala 310:36:freechips.rocketchip.system.DefaultRV32Config.fir@180051.4]
  wire [13:0] tlb_ma_st_array; // @[TLB.scala 310:24:freechips.rocketchip.system.DefaultRV32Config.fir@180053.4]
  wire [13:0] tlb__T_1999; // @[TLB.scala 311:45:freechips.rocketchip.system.DefaultRV32Config.fir@180054.4]
  wire [13:0] tlb__T_2000; // @[TLB.scala 311:35:freechips.rocketchip.system.DefaultRV32Config.fir@180055.4]
  wire [13:0] tlb_pf_ld_array; // @[TLB.scala 311:24:freechips.rocketchip.system.DefaultRV32Config.fir@180056.4]
  wire [13:0] tlb__T_2001; // @[TLB.scala 312:52:freechips.rocketchip.system.DefaultRV32Config.fir@180057.4]
  wire [13:0] tlb__T_2002; // @[TLB.scala 312:42:freechips.rocketchip.system.DefaultRV32Config.fir@180058.4]
  wire [13:0] tlb_pf_st_array; // @[TLB.scala 312:24:freechips.rocketchip.system.DefaultRV32Config.fir@180059.4]
  wire  tlb_tlb_hit; // @[TLB.scala 315:27:freechips.rocketchip.system.DefaultRV32Config.fir@180062.4]
  wire  tlb__T_2006; // @[TLB.scala 316:43:freechips.rocketchip.system.DefaultRV32Config.fir@180065.4]
  wire  tlb_tlb_miss; // @[TLB.scala 316:40:freechips.rocketchip.system.DefaultRV32Config.fir@180066.4]
  reg [6:0] tlb__T_2007; // @[Replacement.scala 158:30:freechips.rocketchip.system.DefaultRV32Config.fir@180067.4]
  reg [2:0] tlb__T_2008; // @[Replacement.scala 158:30:freechips.rocketchip.system.DefaultRV32Config.fir@180068.4]
  wire  tlb__T_2009; // @[TLB.scala 320:22:freechips.rocketchip.system.DefaultRV32Config.fir@180069.4]
  wire  tlb__T_2010; // @[package.scala 64:59:freechips.rocketchip.system.DefaultRV32Config.fir@180071.6]
  wire  tlb__T_2011; // @[package.scala 64:59:freechips.rocketchip.system.DefaultRV32Config.fir@180072.6]
  wire  tlb__T_2012; // @[package.scala 64:59:freechips.rocketchip.system.DefaultRV32Config.fir@180073.6]
  wire  tlb__T_2013; // @[package.scala 64:59:freechips.rocketchip.system.DefaultRV32Config.fir@180074.6]
  wire  tlb__T_2014; // @[package.scala 64:59:freechips.rocketchip.system.DefaultRV32Config.fir@180075.6]
  wire  tlb__T_2015; // @[package.scala 64:59:freechips.rocketchip.system.DefaultRV32Config.fir@180076.6]
  wire  tlb__T_2016; // @[package.scala 64:59:freechips.rocketchip.system.DefaultRV32Config.fir@180077.6]
  wire [7:0] tlb__T_2023; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@180085.8]
  wire [3:0] tlb__T_2024; // @[OneHot.scala 30:18:freechips.rocketchip.system.DefaultRV32Config.fir@180086.8]
  wire [3:0] tlb__T_2025; // @[OneHot.scala 31:18:freechips.rocketchip.system.DefaultRV32Config.fir@180087.8]
  wire  tlb__T_2026; // @[OneHot.scala 32:14:freechips.rocketchip.system.DefaultRV32Config.fir@180088.8]
  wire [3:0] tlb__T_2027; // @[OneHot.scala 32:28:freechips.rocketchip.system.DefaultRV32Config.fir@180089.8]
  wire [1:0] tlb__T_2028; // @[OneHot.scala 30:18:freechips.rocketchip.system.DefaultRV32Config.fir@180090.8]
  wire [1:0] tlb__T_2029; // @[OneHot.scala 31:18:freechips.rocketchip.system.DefaultRV32Config.fir@180091.8]
  wire  tlb__T_2030; // @[OneHot.scala 32:14:freechips.rocketchip.system.DefaultRV32Config.fir@180092.8]
  wire [1:0] tlb__T_2031; // @[OneHot.scala 32:28:freechips.rocketchip.system.DefaultRV32Config.fir@180093.8]
  wire  tlb__T_2032; // @[CircuitMath.scala 30:8:freechips.rocketchip.system.DefaultRV32Config.fir@180094.8]
  wire [2:0] tlb__T_2034; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@180096.8]
  wire  tlb__T_2036; // @[Replacement.scala 186:43:freechips.rocketchip.system.DefaultRV32Config.fir@180098.8]
  wire  tlb__T_2037; // @[Replacement.scala 186:33:freechips.rocketchip.system.DefaultRV32Config.fir@180099.8]
  wire [2:0] tlb__T_2038; // @[package.scala 138:13:freechips.rocketchip.system.DefaultRV32Config.fir@180100.8]
  wire [2:0] tlb__T_2039; // @[Replacement.scala 188:38:freechips.rocketchip.system.DefaultRV32Config.fir@180101.8]
  wire [1:0] tlb__T_2040; // @[package.scala 138:13:freechips.rocketchip.system.DefaultRV32Config.fir@180102.8]
  wire  tlb__T_2041; // @[Replacement.scala 186:43:freechips.rocketchip.system.DefaultRV32Config.fir@180103.8]
  wire  tlb__T_2042; // @[Replacement.scala 186:33:freechips.rocketchip.system.DefaultRV32Config.fir@180104.8]
  wire  tlb__T_2043; // @[package.scala 138:13:freechips.rocketchip.system.DefaultRV32Config.fir@180105.8]
  wire  tlb__T_2044; // @[Replacement.scala 188:38:freechips.rocketchip.system.DefaultRV32Config.fir@180106.8]
  wire  tlb__T_2045; // @[package.scala 138:13:freechips.rocketchip.system.DefaultRV32Config.fir@180107.8]
  wire  tlb__T_2047; // @[Replacement.scala 208:7:freechips.rocketchip.system.DefaultRV32Config.fir@180109.8]
  wire  tlb__T_2048; // @[Replacement.scala 193:16:freechips.rocketchip.system.DefaultRV32Config.fir@180110.8]
  wire  tlb__T_2052; // @[Replacement.scala 196:16:freechips.rocketchip.system.DefaultRV32Config.fir@180114.8]
  wire [2:0] tlb__T_2054; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@180116.8]
  wire [2:0] tlb__T_2055; // @[Replacement.scala 193:16:freechips.rocketchip.system.DefaultRV32Config.fir@180117.8]
  wire  tlb__T_2059; // @[package.scala 138:13:freechips.rocketchip.system.DefaultRV32Config.fir@180121.8]
  wire  tlb__T_2060; // @[Replacement.scala 188:38:freechips.rocketchip.system.DefaultRV32Config.fir@180122.8]
  wire  tlb__T_2064; // @[Replacement.scala 193:16:freechips.rocketchip.system.DefaultRV32Config.fir@180126.8]
  wire  tlb__T_2068; // @[Replacement.scala 196:16:freechips.rocketchip.system.DefaultRV32Config.fir@180130.8]
  wire [2:0] tlb__T_2070; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@180132.8]
  wire [2:0] tlb__T_2071; // @[Replacement.scala 196:16:freechips.rocketchip.system.DefaultRV32Config.fir@180133.8]
  wire [6:0] tlb__T_2073; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@180135.8]
  wire  tlb__T_2074; // @[package.scala 64:59:freechips.rocketchip.system.DefaultRV32Config.fir@180138.6]
  wire  tlb__T_2075; // @[package.scala 64:59:freechips.rocketchip.system.DefaultRV32Config.fir@180139.6]
  wire  tlb__T_2076; // @[package.scala 64:59:freechips.rocketchip.system.DefaultRV32Config.fir@180140.6]
  wire [3:0] tlb__T_2079; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@180144.8]
  wire [1:0] tlb__T_2080; // @[OneHot.scala 30:18:freechips.rocketchip.system.DefaultRV32Config.fir@180145.8]
  wire [1:0] tlb__T_2081; // @[OneHot.scala 31:18:freechips.rocketchip.system.DefaultRV32Config.fir@180146.8]
  wire  tlb__T_2082; // @[OneHot.scala 32:14:freechips.rocketchip.system.DefaultRV32Config.fir@180147.8]
  wire [1:0] tlb__T_2083; // @[OneHot.scala 32:28:freechips.rocketchip.system.DefaultRV32Config.fir@180148.8]
  wire  tlb__T_2084; // @[CircuitMath.scala 30:8:freechips.rocketchip.system.DefaultRV32Config.fir@180149.8]
  wire [1:0] tlb__T_2085; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@180150.8]
  wire  tlb__T_2087; // @[Replacement.scala 186:43:freechips.rocketchip.system.DefaultRV32Config.fir@180152.8]
  wire  tlb__T_2088; // @[Replacement.scala 186:33:freechips.rocketchip.system.DefaultRV32Config.fir@180153.8]
  wire  tlb__T_2089; // @[package.scala 138:13:freechips.rocketchip.system.DefaultRV32Config.fir@180154.8]
  wire  tlb__T_2090; // @[Replacement.scala 188:38:freechips.rocketchip.system.DefaultRV32Config.fir@180155.8]
  wire  tlb__T_2091; // @[package.scala 138:13:freechips.rocketchip.system.DefaultRV32Config.fir@180156.8]
  wire  tlb__T_2093; // @[Replacement.scala 208:7:freechips.rocketchip.system.DefaultRV32Config.fir@180158.8]
  wire  tlb__T_2094; // @[Replacement.scala 193:16:freechips.rocketchip.system.DefaultRV32Config.fir@180159.8]
  wire  tlb__T_2098; // @[Replacement.scala 196:16:freechips.rocketchip.system.DefaultRV32Config.fir@180163.8]
  wire [2:0] tlb__T_2100; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@180165.8]
  wire [5:0] tlb__T_2101; // @[Misc.scala 180:37:freechips.rocketchip.system.DefaultRV32Config.fir@180169.4]
  wire [2:0] tlb__T_2102; // @[Misc.scala 180:37:freechips.rocketchip.system.DefaultRV32Config.fir@180170.4]
  wire  tlb__T_2103; // @[Misc.scala 180:37:freechips.rocketchip.system.DefaultRV32Config.fir@180171.4]
  wire [1:0] tlb__T_2105; // @[Misc.scala 181:39:freechips.rocketchip.system.DefaultRV32Config.fir@180173.4]
  wire  tlb__T_2106; // @[Misc.scala 180:37:freechips.rocketchip.system.DefaultRV32Config.fir@180174.4]
  wire  tlb__T_2108; // @[Misc.scala 181:39:freechips.rocketchip.system.DefaultRV32Config.fir@180176.4]
  wire  tlb__T_2110; // @[Misc.scala 182:16:freechips.rocketchip.system.DefaultRV32Config.fir@180178.4]
  wire  tlb__T_2112; // @[Misc.scala 182:61:freechips.rocketchip.system.DefaultRV32Config.fir@180180.4]
  wire  tlb__T_2114; // @[Misc.scala 182:16:freechips.rocketchip.system.DefaultRV32Config.fir@180182.4]
  wire  tlb__T_2116; // @[Misc.scala 182:61:freechips.rocketchip.system.DefaultRV32Config.fir@180184.4]
  wire  tlb__T_2117; // @[Misc.scala 182:49:freechips.rocketchip.system.DefaultRV32Config.fir@180185.4]
  wire [2:0] tlb__T_2118; // @[Misc.scala 181:39:freechips.rocketchip.system.DefaultRV32Config.fir@180186.4]
  wire  tlb__T_2119; // @[Misc.scala 180:37:freechips.rocketchip.system.DefaultRV32Config.fir@180187.4]
  wire [1:0] tlb__T_2121; // @[Misc.scala 181:39:freechips.rocketchip.system.DefaultRV32Config.fir@180189.4]
  wire  tlb__T_2122; // @[Misc.scala 180:37:freechips.rocketchip.system.DefaultRV32Config.fir@180190.4]
  wire  tlb__T_2124; // @[Misc.scala 181:39:freechips.rocketchip.system.DefaultRV32Config.fir@180192.4]
  wire  tlb__T_2126; // @[Misc.scala 182:16:freechips.rocketchip.system.DefaultRV32Config.fir@180194.4]
  wire  tlb__T_2128; // @[Misc.scala 182:61:freechips.rocketchip.system.DefaultRV32Config.fir@180196.4]
  wire  tlb__T_2130; // @[Misc.scala 182:16:freechips.rocketchip.system.DefaultRV32Config.fir@180198.4]
  wire  tlb__T_2132; // @[Misc.scala 182:61:freechips.rocketchip.system.DefaultRV32Config.fir@180200.4]
  wire  tlb__T_2133; // @[Misc.scala 182:49:freechips.rocketchip.system.DefaultRV32Config.fir@180201.4]
  wire  tlb__T_2134; // @[Misc.scala 182:16:freechips.rocketchip.system.DefaultRV32Config.fir@180202.4]
  wire  tlb__T_2135; // @[Misc.scala 182:37:freechips.rocketchip.system.DefaultRV32Config.fir@180203.4]
  wire  tlb__T_2136; // @[Misc.scala 182:61:freechips.rocketchip.system.DefaultRV32Config.fir@180204.4]
  wire  tlb__T_2137; // @[Misc.scala 182:49:freechips.rocketchip.system.DefaultRV32Config.fir@180205.4]
  wire [6:0] tlb__T_2138; // @[Misc.scala 181:39:freechips.rocketchip.system.DefaultRV32Config.fir@180206.4]
  wire [2:0] tlb__T_2139; // @[Misc.scala 180:37:freechips.rocketchip.system.DefaultRV32Config.fir@180207.4]
  wire  tlb__T_2140; // @[Misc.scala 180:37:freechips.rocketchip.system.DefaultRV32Config.fir@180208.4]
  wire [1:0] tlb__T_2142; // @[Misc.scala 181:39:freechips.rocketchip.system.DefaultRV32Config.fir@180210.4]
  wire  tlb__T_2143; // @[Misc.scala 180:37:freechips.rocketchip.system.DefaultRV32Config.fir@180211.4]
  wire  tlb__T_2145; // @[Misc.scala 181:39:freechips.rocketchip.system.DefaultRV32Config.fir@180213.4]
  wire  tlb__T_2147; // @[Misc.scala 182:16:freechips.rocketchip.system.DefaultRV32Config.fir@180215.4]
  wire  tlb__T_2149; // @[Misc.scala 182:61:freechips.rocketchip.system.DefaultRV32Config.fir@180217.4]
  wire  tlb__T_2151; // @[Misc.scala 182:16:freechips.rocketchip.system.DefaultRV32Config.fir@180219.4]
  wire  tlb__T_2153; // @[Misc.scala 182:61:freechips.rocketchip.system.DefaultRV32Config.fir@180221.4]
  wire  tlb__T_2154; // @[Misc.scala 182:49:freechips.rocketchip.system.DefaultRV32Config.fir@180222.4]
  wire [3:0] tlb__T_2155; // @[Misc.scala 181:39:freechips.rocketchip.system.DefaultRV32Config.fir@180223.4]
  wire [1:0] tlb__T_2156; // @[Misc.scala 180:37:freechips.rocketchip.system.DefaultRV32Config.fir@180224.4]
  wire  tlb__T_2157; // @[Misc.scala 180:37:freechips.rocketchip.system.DefaultRV32Config.fir@180225.4]
  wire  tlb__T_2159; // @[Misc.scala 181:39:freechips.rocketchip.system.DefaultRV32Config.fir@180227.4]
  wire  tlb__T_2161; // @[Misc.scala 182:16:freechips.rocketchip.system.DefaultRV32Config.fir@180229.4]
  wire  tlb__T_2163; // @[Misc.scala 182:61:freechips.rocketchip.system.DefaultRV32Config.fir@180231.4]
  wire [1:0] tlb__T_2165; // @[Misc.scala 181:39:freechips.rocketchip.system.DefaultRV32Config.fir@180233.4]
  wire  tlb__T_2166; // @[Misc.scala 180:37:freechips.rocketchip.system.DefaultRV32Config.fir@180234.4]
  wire  tlb__T_2168; // @[Misc.scala 181:39:freechips.rocketchip.system.DefaultRV32Config.fir@180236.4]
  wire  tlb__T_2170; // @[Misc.scala 182:16:freechips.rocketchip.system.DefaultRV32Config.fir@180238.4]
  wire  tlb__T_2172; // @[Misc.scala 182:61:freechips.rocketchip.system.DefaultRV32Config.fir@180240.4]
  wire  tlb__T_2174; // @[Misc.scala 182:16:freechips.rocketchip.system.DefaultRV32Config.fir@180242.4]
  wire  tlb__T_2175; // @[Misc.scala 182:37:freechips.rocketchip.system.DefaultRV32Config.fir@180243.4]
  wire  tlb__T_2176; // @[Misc.scala 182:61:freechips.rocketchip.system.DefaultRV32Config.fir@180244.4]
  wire  tlb__T_2177; // @[Misc.scala 182:49:freechips.rocketchip.system.DefaultRV32Config.fir@180245.4]
  wire  tlb__T_2178; // @[Misc.scala 182:16:freechips.rocketchip.system.DefaultRV32Config.fir@180246.4]
  wire  tlb__T_2179; // @[Misc.scala 182:37:freechips.rocketchip.system.DefaultRV32Config.fir@180247.4]
  wire  tlb__T_2180; // @[Misc.scala 182:61:freechips.rocketchip.system.DefaultRV32Config.fir@180248.4]
  wire  tlb__T_2181; // @[Misc.scala 182:49:freechips.rocketchip.system.DefaultRV32Config.fir@180249.4]
  wire  tlb__T_2183; // @[Misc.scala 182:37:freechips.rocketchip.system.DefaultRV32Config.fir@180251.4]
  wire  tlb__T_2184; // @[Misc.scala 182:61:freechips.rocketchip.system.DefaultRV32Config.fir@180252.4]
  wire  tlb_multipleHits; // @[Misc.scala 182:49:freechips.rocketchip.system.DefaultRV32Config.fir@180253.4]
  wire [13:0] tlb__T_2187; // @[TLB.scala 333:57:freechips.rocketchip.system.DefaultRV32Config.fir@180257.4]
  wire [13:0] tlb__T_2191; // @[TLB.scala 334:64:freechips.rocketchip.system.DefaultRV32Config.fir@180262.4]
  wire [13:0] tlb__T_2197; // @[TLB.scala 336:33:freechips.rocketchip.system.DefaultRV32Config.fir@180270.4]
  wire [13:0] tlb__T_2199; // @[TLB.scala 337:33:freechips.rocketchip.system.DefaultRV32Config.fir@180273.4]
  wire [13:0] tlb__T_2204; // @[TLB.scala 339:33:freechips.rocketchip.system.DefaultRV32Config.fir@180280.4]
  wire [13:0] tlb__T_2206; // @[TLB.scala 340:33:freechips.rocketchip.system.DefaultRV32Config.fir@180283.4]
  wire [13:0] tlb__T_2208; // @[TLB.scala 342:33:freechips.rocketchip.system.DefaultRV32Config.fir@180287.4]
  wire  tlb__T_2215; // @[TLB.scala 345:29:freechips.rocketchip.system.DefaultRV32Config.fir@180297.4]
  wire  tlb__T_2221; // @[Decoupled.scala 40:37:freechips.rocketchip.system.DefaultRV32Config.fir@180308.4]
  wire  tlb__T_2222; // @[TLB.scala 354:25:freechips.rocketchip.system.DefaultRV32Config.fir@180309.4]
  wire  tlb__T_2223; // @[Replacement.scala 233:38:freechips.rocketchip.system.DefaultRV32Config.fir@180313.6]
  wire  tlb__T_2228; // @[Replacement.scala 240:16:freechips.rocketchip.system.DefaultRV32Config.fir@180318.6]
  wire [1:0] tlb__T_2229; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@180319.6]
  wire [3:0] tlb__T_2232; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@180322.6]
  wire  tlb__T_2233; // @[TLB.scala 402:16:freechips.rocketchip.system.DefaultRV32Config.fir@180323.6]
  wire [3:0] tlb__T_2234; // @[TLB.scala 402:43:freechips.rocketchip.system.DefaultRV32Config.fir@180324.6]
  wire  tlb__T_2235; // @[OneHot.scala 47:40:freechips.rocketchip.system.DefaultRV32Config.fir@180325.6]
  wire  tlb__T_2236; // @[OneHot.scala 47:40:freechips.rocketchip.system.DefaultRV32Config.fir@180326.6]
  wire  tlb__T_2237; // @[OneHot.scala 47:40:freechips.rocketchip.system.DefaultRV32Config.fir@180327.6]
  wire  tlb__T_2243; // @[Replacement.scala 233:38:freechips.rocketchip.system.DefaultRV32Config.fir@180334.6]
  wire  tlb__T_2246; // @[Replacement.scala 233:38:freechips.rocketchip.system.DefaultRV32Config.fir@180337.6]
  wire  tlb__T_2251; // @[Replacement.scala 240:16:freechips.rocketchip.system.DefaultRV32Config.fir@180342.6]
  wire [1:0] tlb__T_2252; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@180343.6]
  wire  tlb__T_2253; // @[Replacement.scala 233:38:freechips.rocketchip.system.DefaultRV32Config.fir@180344.6]
  wire  tlb__T_2258; // @[Replacement.scala 240:16:freechips.rocketchip.system.DefaultRV32Config.fir@180349.6]
  wire [1:0] tlb__T_2259; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@180350.6]
  wire [1:0] tlb__T_2260; // @[Replacement.scala 240:16:freechips.rocketchip.system.DefaultRV32Config.fir@180351.6]
  wire [2:0] tlb__T_2261; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@180352.6]
  wire [7:0] tlb__T_2292; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@180383.6]
  wire  tlb__T_2293; // @[TLB.scala 402:16:freechips.rocketchip.system.DefaultRV32Config.fir@180384.6]
  wire [7:0] tlb__T_2294; // @[TLB.scala 402:43:freechips.rocketchip.system.DefaultRV32Config.fir@180385.6]
  wire  tlb__T_2295; // @[OneHot.scala 47:40:freechips.rocketchip.system.DefaultRV32Config.fir@180386.6]
  wire  tlb__T_2296; // @[OneHot.scala 47:40:freechips.rocketchip.system.DefaultRV32Config.fir@180387.6]
  wire  tlb__T_2297; // @[OneHot.scala 47:40:freechips.rocketchip.system.DefaultRV32Config.fir@180388.6]
  wire  tlb__T_2298; // @[OneHot.scala 47:40:freechips.rocketchip.system.DefaultRV32Config.fir@180389.6]
  wire  tlb__T_2299; // @[OneHot.scala 47:40:freechips.rocketchip.system.DefaultRV32Config.fir@180390.6]
  wire  tlb__T_2300; // @[OneHot.scala 47:40:freechips.rocketchip.system.DefaultRV32Config.fir@180391.6]
  wire  tlb__T_2301; // @[OneHot.scala 47:40:freechips.rocketchip.system.DefaultRV32Config.fir@180392.6]
  wire  tlb__T_2338; // @[TLB.scala 368:17:freechips.rocketchip.system.DefaultRV32Config.fir@180444.4]
  wire  tlb__T_2339; // @[TLB.scala 368:28:freechips.rocketchip.system.DefaultRV32Config.fir@180445.4]
  wire  tlb__T_2340; // @[TLB.scala 376:14:freechips.rocketchip.system.DefaultRV32Config.fir@180453.6]
  wire [19:0] tlb__T_2341; // @[TLB.scala 376:58:freechips.rocketchip.system.DefaultRV32Config.fir@180454.6]
  wire  tlb__T_2342; // @[TLB.scala 376:72:freechips.rocketchip.system.DefaultRV32Config.fir@180455.6]
  wire  tlb__T_2343; // @[TLB.scala 376:34:freechips.rocketchip.system.DefaultRV32Config.fir@180456.6]
  wire  tlb__T_2345; // @[TLB.scala 376:13:freechips.rocketchip.system.DefaultRV32Config.fir@180458.6]
  wire  tlb__T_2346; // @[TLB.scala 376:13:freechips.rocketchip.system.DefaultRV32Config.fir@180459.6]
  wire [9:0] tlb__T_2352; // @[TLB.scala 135:26:freechips.rocketchip.system.DefaultRV32Config.fir@180473.8]
  wire  tlb__T_2353; // @[TLB.scala 135:61:freechips.rocketchip.system.DefaultRV32Config.fir@180474.8]
  wire  tlb__T_2356; // @[TLB.scala 83:39:freechips.rocketchip.system.DefaultRV32Config.fir@180481.10]
  wire  tlb__T_2369; // @[TLB.scala 83:39:freechips.rocketchip.system.DefaultRV32Config.fir@180507.10]
  wire  tlb__T_2374; // @[TLB.scala 83:39:freechips.rocketchip.system.DefaultRV32Config.fir@180518.10]
  wire  tlb__T_2387; // @[TLB.scala 83:39:freechips.rocketchip.system.DefaultRV32Config.fir@180544.10]
  wire  tlb__T_2392; // @[TLB.scala 83:39:freechips.rocketchip.system.DefaultRV32Config.fir@180555.10]
  wire  tlb__T_2405; // @[TLB.scala 83:39:freechips.rocketchip.system.DefaultRV32Config.fir@180581.10]
  wire  tlb__T_2410; // @[TLB.scala 83:39:freechips.rocketchip.system.DefaultRV32Config.fir@180592.10]
  wire  tlb__T_2423; // @[TLB.scala 83:39:freechips.rocketchip.system.DefaultRV32Config.fir@180618.10]
  wire  tlb__T_2498; // @[TLB.scala 143:13:freechips.rocketchip.system.DefaultRV32Config.fir@180788.10]
  wire  tlb__GEN_648; // @[TLB.scala 143:19:freechips.rocketchip.system.DefaultRV32Config.fir@180789.10]
  wire  tlb__T_2499; // @[TLB.scala 143:13:freechips.rocketchip.system.DefaultRV32Config.fir@180792.10]
  wire  tlb__GEN_649; // @[TLB.scala 143:19:freechips.rocketchip.system.DefaultRV32Config.fir@180793.10]
  wire  tlb__T_2500; // @[TLB.scala 143:13:freechips.rocketchip.system.DefaultRV32Config.fir@180796.10]
  wire  tlb__GEN_650; // @[TLB.scala 143:19:freechips.rocketchip.system.DefaultRV32Config.fir@180797.10]
  wire  tlb__T_2501; // @[TLB.scala 143:13:freechips.rocketchip.system.DefaultRV32Config.fir@180800.10]
  wire  tlb__GEN_651; // @[TLB.scala 143:19:freechips.rocketchip.system.DefaultRV32Config.fir@180801.10]
  wire  tlb__GEN_652; // @[TLB.scala 379:40:freechips.rocketchip.system.DefaultRV32Config.fir@180639.8]
  wire  tlb__GEN_653; // @[TLB.scala 379:40:freechips.rocketchip.system.DefaultRV32Config.fir@180639.8]
  wire  tlb__GEN_654; // @[TLB.scala 379:40:freechips.rocketchip.system.DefaultRV32Config.fir@180639.8]
  wire  tlb__GEN_655; // @[TLB.scala 379:40:freechips.rocketchip.system.DefaultRV32Config.fir@180639.8]
  wire [9:0] tlb__T_2507; // @[TLB.scala 135:26:freechips.rocketchip.system.DefaultRV32Config.fir@180820.8]
  wire  tlb__T_2508; // @[TLB.scala 135:61:freechips.rocketchip.system.DefaultRV32Config.fir@180821.8]
  wire  tlb__T_2511; // @[TLB.scala 83:39:freechips.rocketchip.system.DefaultRV32Config.fir@180828.10]
  wire  tlb__T_2524; // @[TLB.scala 83:39:freechips.rocketchip.system.DefaultRV32Config.fir@180854.10]
  wire  tlb__T_2529; // @[TLB.scala 83:39:freechips.rocketchip.system.DefaultRV32Config.fir@180865.10]
  wire  tlb__T_2542; // @[TLB.scala 83:39:freechips.rocketchip.system.DefaultRV32Config.fir@180891.10]
  wire  tlb__T_2547; // @[TLB.scala 83:39:freechips.rocketchip.system.DefaultRV32Config.fir@180902.10]
  wire  tlb__T_2560; // @[TLB.scala 83:39:freechips.rocketchip.system.DefaultRV32Config.fir@180928.10]
  wire  tlb__T_2565; // @[TLB.scala 83:39:freechips.rocketchip.system.DefaultRV32Config.fir@180939.10]
  wire  tlb__T_2578; // @[TLB.scala 83:39:freechips.rocketchip.system.DefaultRV32Config.fir@180965.10]
  wire  tlb__T_2653; // @[TLB.scala 143:13:freechips.rocketchip.system.DefaultRV32Config.fir@181135.10]
  wire  tlb__GEN_676; // @[TLB.scala 143:19:freechips.rocketchip.system.DefaultRV32Config.fir@181136.10]
  wire  tlb__T_2654; // @[TLB.scala 143:13:freechips.rocketchip.system.DefaultRV32Config.fir@181139.10]
  wire  tlb__GEN_677; // @[TLB.scala 143:19:freechips.rocketchip.system.DefaultRV32Config.fir@181140.10]
  wire  tlb__T_2655; // @[TLB.scala 143:13:freechips.rocketchip.system.DefaultRV32Config.fir@181143.10]
  wire  tlb__GEN_678; // @[TLB.scala 143:19:freechips.rocketchip.system.DefaultRV32Config.fir@181144.10]
  wire  tlb__T_2656; // @[TLB.scala 143:13:freechips.rocketchip.system.DefaultRV32Config.fir@181147.10]
  wire  tlb__GEN_679; // @[TLB.scala 143:19:freechips.rocketchip.system.DefaultRV32Config.fir@181148.10]
  wire  tlb__GEN_680; // @[TLB.scala 379:40:freechips.rocketchip.system.DefaultRV32Config.fir@180986.8]
  wire  tlb__GEN_681; // @[TLB.scala 379:40:freechips.rocketchip.system.DefaultRV32Config.fir@180986.8]
  wire  tlb__GEN_682; // @[TLB.scala 379:40:freechips.rocketchip.system.DefaultRV32Config.fir@180986.8]
  wire  tlb__GEN_683; // @[TLB.scala 379:40:freechips.rocketchip.system.DefaultRV32Config.fir@180986.8]
  wire [9:0] tlb__T_2662; // @[TLB.scala 135:26:freechips.rocketchip.system.DefaultRV32Config.fir@181167.8]
  wire  tlb__T_2663; // @[TLB.scala 135:61:freechips.rocketchip.system.DefaultRV32Config.fir@181168.8]
  wire  tlb__T_2666; // @[TLB.scala 83:39:freechips.rocketchip.system.DefaultRV32Config.fir@181175.10]
  wire  tlb__T_2679; // @[TLB.scala 83:39:freechips.rocketchip.system.DefaultRV32Config.fir@181201.10]
  wire  tlb__T_2684; // @[TLB.scala 83:39:freechips.rocketchip.system.DefaultRV32Config.fir@181212.10]
  wire  tlb__T_2697; // @[TLB.scala 83:39:freechips.rocketchip.system.DefaultRV32Config.fir@181238.10]
  wire  tlb__T_2702; // @[TLB.scala 83:39:freechips.rocketchip.system.DefaultRV32Config.fir@181249.10]
  wire  tlb__T_2715; // @[TLB.scala 83:39:freechips.rocketchip.system.DefaultRV32Config.fir@181275.10]
  wire  tlb__T_2720; // @[TLB.scala 83:39:freechips.rocketchip.system.DefaultRV32Config.fir@181286.10]
  wire  tlb__T_2733; // @[TLB.scala 83:39:freechips.rocketchip.system.DefaultRV32Config.fir@181312.10]
  wire  tlb__T_2808; // @[TLB.scala 143:13:freechips.rocketchip.system.DefaultRV32Config.fir@181482.10]
  wire  tlb__GEN_704; // @[TLB.scala 143:19:freechips.rocketchip.system.DefaultRV32Config.fir@181483.10]
  wire  tlb__T_2809; // @[TLB.scala 143:13:freechips.rocketchip.system.DefaultRV32Config.fir@181486.10]
  wire  tlb__GEN_705; // @[TLB.scala 143:19:freechips.rocketchip.system.DefaultRV32Config.fir@181487.10]
  wire  tlb__T_2810; // @[TLB.scala 143:13:freechips.rocketchip.system.DefaultRV32Config.fir@181490.10]
  wire  tlb__GEN_706; // @[TLB.scala 143:19:freechips.rocketchip.system.DefaultRV32Config.fir@181491.10]
  wire  tlb__T_2811; // @[TLB.scala 143:13:freechips.rocketchip.system.DefaultRV32Config.fir@181494.10]
  wire  tlb__GEN_707; // @[TLB.scala 143:19:freechips.rocketchip.system.DefaultRV32Config.fir@181495.10]
  wire  tlb__GEN_708; // @[TLB.scala 379:40:freechips.rocketchip.system.DefaultRV32Config.fir@181333.8]
  wire  tlb__GEN_709; // @[TLB.scala 379:40:freechips.rocketchip.system.DefaultRV32Config.fir@181333.8]
  wire  tlb__GEN_710; // @[TLB.scala 379:40:freechips.rocketchip.system.DefaultRV32Config.fir@181333.8]
  wire  tlb__GEN_711; // @[TLB.scala 379:40:freechips.rocketchip.system.DefaultRV32Config.fir@181333.8]
  wire [9:0] tlb__T_2817; // @[TLB.scala 135:26:freechips.rocketchip.system.DefaultRV32Config.fir@181514.8]
  wire  tlb__T_2818; // @[TLB.scala 135:61:freechips.rocketchip.system.DefaultRV32Config.fir@181515.8]
  wire  tlb__T_2821; // @[TLB.scala 83:39:freechips.rocketchip.system.DefaultRV32Config.fir@181522.10]
  wire  tlb__T_2834; // @[TLB.scala 83:39:freechips.rocketchip.system.DefaultRV32Config.fir@181548.10]
  wire  tlb__T_2839; // @[TLB.scala 83:39:freechips.rocketchip.system.DefaultRV32Config.fir@181559.10]
  wire  tlb__T_2852; // @[TLB.scala 83:39:freechips.rocketchip.system.DefaultRV32Config.fir@181585.10]
  wire  tlb__T_2857; // @[TLB.scala 83:39:freechips.rocketchip.system.DefaultRV32Config.fir@181596.10]
  wire  tlb__T_2870; // @[TLB.scala 83:39:freechips.rocketchip.system.DefaultRV32Config.fir@181622.10]
  wire  tlb__T_2875; // @[TLB.scala 83:39:freechips.rocketchip.system.DefaultRV32Config.fir@181633.10]
  wire  tlb__T_2888; // @[TLB.scala 83:39:freechips.rocketchip.system.DefaultRV32Config.fir@181659.10]
  wire  tlb__T_2963; // @[TLB.scala 143:13:freechips.rocketchip.system.DefaultRV32Config.fir@181829.10]
  wire  tlb__GEN_732; // @[TLB.scala 143:19:freechips.rocketchip.system.DefaultRV32Config.fir@181830.10]
  wire  tlb__T_2964; // @[TLB.scala 143:13:freechips.rocketchip.system.DefaultRV32Config.fir@181833.10]
  wire  tlb__GEN_733; // @[TLB.scala 143:19:freechips.rocketchip.system.DefaultRV32Config.fir@181834.10]
  wire  tlb__T_2965; // @[TLB.scala 143:13:freechips.rocketchip.system.DefaultRV32Config.fir@181837.10]
  wire  tlb__GEN_734; // @[TLB.scala 143:19:freechips.rocketchip.system.DefaultRV32Config.fir@181838.10]
  wire  tlb__T_2966; // @[TLB.scala 143:13:freechips.rocketchip.system.DefaultRV32Config.fir@181841.10]
  wire  tlb__GEN_735; // @[TLB.scala 143:19:freechips.rocketchip.system.DefaultRV32Config.fir@181842.10]
  wire  tlb__GEN_736; // @[TLB.scala 379:40:freechips.rocketchip.system.DefaultRV32Config.fir@181680.8]
  wire  tlb__GEN_737; // @[TLB.scala 379:40:freechips.rocketchip.system.DefaultRV32Config.fir@181680.8]
  wire  tlb__GEN_738; // @[TLB.scala 379:40:freechips.rocketchip.system.DefaultRV32Config.fir@181680.8]
  wire  tlb__GEN_739; // @[TLB.scala 379:40:freechips.rocketchip.system.DefaultRV32Config.fir@181680.8]
  wire [9:0] tlb__T_2972; // @[TLB.scala 135:26:freechips.rocketchip.system.DefaultRV32Config.fir@181861.8]
  wire  tlb__T_2973; // @[TLB.scala 135:61:freechips.rocketchip.system.DefaultRV32Config.fir@181862.8]
  wire  tlb__T_2976; // @[TLB.scala 83:39:freechips.rocketchip.system.DefaultRV32Config.fir@181869.10]
  wire  tlb__T_2989; // @[TLB.scala 83:39:freechips.rocketchip.system.DefaultRV32Config.fir@181895.10]
  wire  tlb__T_2994; // @[TLB.scala 83:39:freechips.rocketchip.system.DefaultRV32Config.fir@181906.10]
  wire  tlb__T_3007; // @[TLB.scala 83:39:freechips.rocketchip.system.DefaultRV32Config.fir@181932.10]
  wire  tlb__T_3012; // @[TLB.scala 83:39:freechips.rocketchip.system.DefaultRV32Config.fir@181943.10]
  wire  tlb__T_3025; // @[TLB.scala 83:39:freechips.rocketchip.system.DefaultRV32Config.fir@181969.10]
  wire  tlb__T_3030; // @[TLB.scala 83:39:freechips.rocketchip.system.DefaultRV32Config.fir@181980.10]
  wire  tlb__T_3043; // @[TLB.scala 83:39:freechips.rocketchip.system.DefaultRV32Config.fir@182006.10]
  wire  tlb__T_3118; // @[TLB.scala 143:13:freechips.rocketchip.system.DefaultRV32Config.fir@182176.10]
  wire  tlb__GEN_760; // @[TLB.scala 143:19:freechips.rocketchip.system.DefaultRV32Config.fir@182177.10]
  wire  tlb__T_3119; // @[TLB.scala 143:13:freechips.rocketchip.system.DefaultRV32Config.fir@182180.10]
  wire  tlb__GEN_761; // @[TLB.scala 143:19:freechips.rocketchip.system.DefaultRV32Config.fir@182181.10]
  wire  tlb__T_3120; // @[TLB.scala 143:13:freechips.rocketchip.system.DefaultRV32Config.fir@182184.10]
  wire  tlb__GEN_762; // @[TLB.scala 143:19:freechips.rocketchip.system.DefaultRV32Config.fir@182185.10]
  wire  tlb__T_3121; // @[TLB.scala 143:13:freechips.rocketchip.system.DefaultRV32Config.fir@182188.10]
  wire  tlb__GEN_763; // @[TLB.scala 143:19:freechips.rocketchip.system.DefaultRV32Config.fir@182189.10]
  wire  tlb__GEN_764; // @[TLB.scala 379:40:freechips.rocketchip.system.DefaultRV32Config.fir@182027.8]
  wire  tlb__GEN_765; // @[TLB.scala 379:40:freechips.rocketchip.system.DefaultRV32Config.fir@182027.8]
  wire  tlb__GEN_766; // @[TLB.scala 379:40:freechips.rocketchip.system.DefaultRV32Config.fir@182027.8]
  wire  tlb__GEN_767; // @[TLB.scala 379:40:freechips.rocketchip.system.DefaultRV32Config.fir@182027.8]
  wire [9:0] tlb__T_3127; // @[TLB.scala 135:26:freechips.rocketchip.system.DefaultRV32Config.fir@182208.8]
  wire  tlb__T_3128; // @[TLB.scala 135:61:freechips.rocketchip.system.DefaultRV32Config.fir@182209.8]
  wire  tlb__T_3131; // @[TLB.scala 83:39:freechips.rocketchip.system.DefaultRV32Config.fir@182216.10]
  wire  tlb__T_3144; // @[TLB.scala 83:39:freechips.rocketchip.system.DefaultRV32Config.fir@182242.10]
  wire  tlb__T_3149; // @[TLB.scala 83:39:freechips.rocketchip.system.DefaultRV32Config.fir@182253.10]
  wire  tlb__T_3162; // @[TLB.scala 83:39:freechips.rocketchip.system.DefaultRV32Config.fir@182279.10]
  wire  tlb__T_3167; // @[TLB.scala 83:39:freechips.rocketchip.system.DefaultRV32Config.fir@182290.10]
  wire  tlb__T_3180; // @[TLB.scala 83:39:freechips.rocketchip.system.DefaultRV32Config.fir@182316.10]
  wire  tlb__T_3185; // @[TLB.scala 83:39:freechips.rocketchip.system.DefaultRV32Config.fir@182327.10]
  wire  tlb__T_3198; // @[TLB.scala 83:39:freechips.rocketchip.system.DefaultRV32Config.fir@182353.10]
  wire  tlb__T_3273; // @[TLB.scala 143:13:freechips.rocketchip.system.DefaultRV32Config.fir@182523.10]
  wire  tlb__GEN_788; // @[TLB.scala 143:19:freechips.rocketchip.system.DefaultRV32Config.fir@182524.10]
  wire  tlb__T_3274; // @[TLB.scala 143:13:freechips.rocketchip.system.DefaultRV32Config.fir@182527.10]
  wire  tlb__GEN_789; // @[TLB.scala 143:19:freechips.rocketchip.system.DefaultRV32Config.fir@182528.10]
  wire  tlb__T_3275; // @[TLB.scala 143:13:freechips.rocketchip.system.DefaultRV32Config.fir@182531.10]
  wire  tlb__GEN_790; // @[TLB.scala 143:19:freechips.rocketchip.system.DefaultRV32Config.fir@182532.10]
  wire  tlb__T_3276; // @[TLB.scala 143:13:freechips.rocketchip.system.DefaultRV32Config.fir@182535.10]
  wire  tlb__GEN_791; // @[TLB.scala 143:19:freechips.rocketchip.system.DefaultRV32Config.fir@182536.10]
  wire  tlb__GEN_792; // @[TLB.scala 379:40:freechips.rocketchip.system.DefaultRV32Config.fir@182374.8]
  wire  tlb__GEN_793; // @[TLB.scala 379:40:freechips.rocketchip.system.DefaultRV32Config.fir@182374.8]
  wire  tlb__GEN_794; // @[TLB.scala 379:40:freechips.rocketchip.system.DefaultRV32Config.fir@182374.8]
  wire  tlb__GEN_795; // @[TLB.scala 379:40:freechips.rocketchip.system.DefaultRV32Config.fir@182374.8]
  wire [9:0] tlb__T_3282; // @[TLB.scala 135:26:freechips.rocketchip.system.DefaultRV32Config.fir@182555.8]
  wire  tlb__T_3283; // @[TLB.scala 135:61:freechips.rocketchip.system.DefaultRV32Config.fir@182556.8]
  wire  tlb__T_3286; // @[TLB.scala 83:39:freechips.rocketchip.system.DefaultRV32Config.fir@182563.10]
  wire  tlb__T_3299; // @[TLB.scala 83:39:freechips.rocketchip.system.DefaultRV32Config.fir@182589.10]
  wire  tlb__T_3304; // @[TLB.scala 83:39:freechips.rocketchip.system.DefaultRV32Config.fir@182600.10]
  wire  tlb__T_3317; // @[TLB.scala 83:39:freechips.rocketchip.system.DefaultRV32Config.fir@182626.10]
  wire  tlb__T_3322; // @[TLB.scala 83:39:freechips.rocketchip.system.DefaultRV32Config.fir@182637.10]
  wire  tlb__T_3335; // @[TLB.scala 83:39:freechips.rocketchip.system.DefaultRV32Config.fir@182663.10]
  wire  tlb__T_3340; // @[TLB.scala 83:39:freechips.rocketchip.system.DefaultRV32Config.fir@182674.10]
  wire  tlb__T_3353; // @[TLB.scala 83:39:freechips.rocketchip.system.DefaultRV32Config.fir@182700.10]
  wire  tlb__T_3428; // @[TLB.scala 143:13:freechips.rocketchip.system.DefaultRV32Config.fir@182870.10]
  wire  tlb__GEN_816; // @[TLB.scala 143:19:freechips.rocketchip.system.DefaultRV32Config.fir@182871.10]
  wire  tlb__T_3429; // @[TLB.scala 143:13:freechips.rocketchip.system.DefaultRV32Config.fir@182874.10]
  wire  tlb__GEN_817; // @[TLB.scala 143:19:freechips.rocketchip.system.DefaultRV32Config.fir@182875.10]
  wire  tlb__T_3430; // @[TLB.scala 143:13:freechips.rocketchip.system.DefaultRV32Config.fir@182878.10]
  wire  tlb__GEN_818; // @[TLB.scala 143:19:freechips.rocketchip.system.DefaultRV32Config.fir@182879.10]
  wire  tlb__T_3431; // @[TLB.scala 143:13:freechips.rocketchip.system.DefaultRV32Config.fir@182882.10]
  wire  tlb__GEN_819; // @[TLB.scala 143:19:freechips.rocketchip.system.DefaultRV32Config.fir@182883.10]
  wire  tlb__GEN_820; // @[TLB.scala 379:40:freechips.rocketchip.system.DefaultRV32Config.fir@182721.8]
  wire  tlb__GEN_821; // @[TLB.scala 379:40:freechips.rocketchip.system.DefaultRV32Config.fir@182721.8]
  wire  tlb__GEN_822; // @[TLB.scala 379:40:freechips.rocketchip.system.DefaultRV32Config.fir@182721.8]
  wire  tlb__GEN_823; // @[TLB.scala 379:40:freechips.rocketchip.system.DefaultRV32Config.fir@182721.8]
  wire [9:0] tlb__T_3437; // @[TLB.scala 135:26:freechips.rocketchip.system.DefaultRV32Config.fir@182902.8]
  wire  tlb__T_3438; // @[TLB.scala 135:61:freechips.rocketchip.system.DefaultRV32Config.fir@182903.8]
  wire  tlb__T_3441; // @[TLB.scala 83:39:freechips.rocketchip.system.DefaultRV32Config.fir@182910.10]
  wire  tlb__T_3454; // @[TLB.scala 83:39:freechips.rocketchip.system.DefaultRV32Config.fir@182936.10]
  wire  tlb__T_3459; // @[TLB.scala 83:39:freechips.rocketchip.system.DefaultRV32Config.fir@182947.10]
  wire  tlb__T_3472; // @[TLB.scala 83:39:freechips.rocketchip.system.DefaultRV32Config.fir@182973.10]
  wire  tlb__T_3477; // @[TLB.scala 83:39:freechips.rocketchip.system.DefaultRV32Config.fir@182984.10]
  wire  tlb__T_3490; // @[TLB.scala 83:39:freechips.rocketchip.system.DefaultRV32Config.fir@183010.10]
  wire  tlb__T_3495; // @[TLB.scala 83:39:freechips.rocketchip.system.DefaultRV32Config.fir@183021.10]
  wire  tlb__T_3508; // @[TLB.scala 83:39:freechips.rocketchip.system.DefaultRV32Config.fir@183047.10]
  wire  tlb__T_3583; // @[TLB.scala 143:13:freechips.rocketchip.system.DefaultRV32Config.fir@183217.10]
  wire  tlb__GEN_844; // @[TLB.scala 143:19:freechips.rocketchip.system.DefaultRV32Config.fir@183218.10]
  wire  tlb__T_3584; // @[TLB.scala 143:13:freechips.rocketchip.system.DefaultRV32Config.fir@183221.10]
  wire  tlb__GEN_845; // @[TLB.scala 143:19:freechips.rocketchip.system.DefaultRV32Config.fir@183222.10]
  wire  tlb__T_3585; // @[TLB.scala 143:13:freechips.rocketchip.system.DefaultRV32Config.fir@183225.10]
  wire  tlb__GEN_846; // @[TLB.scala 143:19:freechips.rocketchip.system.DefaultRV32Config.fir@183226.10]
  wire  tlb__T_3586; // @[TLB.scala 143:13:freechips.rocketchip.system.DefaultRV32Config.fir@183229.10]
  wire  tlb__GEN_847; // @[TLB.scala 143:19:freechips.rocketchip.system.DefaultRV32Config.fir@183230.10]
  wire  tlb__GEN_848; // @[TLB.scala 379:40:freechips.rocketchip.system.DefaultRV32Config.fir@183068.8]
  wire  tlb__GEN_849; // @[TLB.scala 379:40:freechips.rocketchip.system.DefaultRV32Config.fir@183068.8]
  wire  tlb__GEN_850; // @[TLB.scala 379:40:freechips.rocketchip.system.DefaultRV32Config.fir@183068.8]
  wire  tlb__GEN_851; // @[TLB.scala 379:40:freechips.rocketchip.system.DefaultRV32Config.fir@183068.8]
  wire  tlb__T_3619; // @[TLB.scala 143:13:freechips.rocketchip.system.DefaultRV32Config.fir@183298.10]
  wire  tlb__GEN_857; // @[TLB.scala 143:19:freechips.rocketchip.system.DefaultRV32Config.fir@183299.10]
  wire  tlb__GEN_858; // @[TLB.scala 379:40:freechips.rocketchip.system.DefaultRV32Config.fir@183260.8]
  wire  tlb__T_3652; // @[TLB.scala 143:13:freechips.rocketchip.system.DefaultRV32Config.fir@183364.10]
  wire  tlb__GEN_861; // @[TLB.scala 143:19:freechips.rocketchip.system.DefaultRV32Config.fir@183365.10]
  wire  tlb__GEN_862; // @[TLB.scala 379:40:freechips.rocketchip.system.DefaultRV32Config.fir@183326.8]
  wire  tlb__T_3685; // @[TLB.scala 143:13:freechips.rocketchip.system.DefaultRV32Config.fir@183430.10]
  wire  tlb__GEN_865; // @[TLB.scala 143:19:freechips.rocketchip.system.DefaultRV32Config.fir@183431.10]
  wire  tlb__GEN_866; // @[TLB.scala 379:40:freechips.rocketchip.system.DefaultRV32Config.fir@183392.8]
  wire  tlb__T_3718; // @[TLB.scala 143:13:freechips.rocketchip.system.DefaultRV32Config.fir@183496.10]
  wire  tlb__GEN_869; // @[TLB.scala 143:19:freechips.rocketchip.system.DefaultRV32Config.fir@183497.10]
  wire  tlb__GEN_870; // @[TLB.scala 379:40:freechips.rocketchip.system.DefaultRV32Config.fir@183458.8]
  wire  tlb__T_3751; // @[TLB.scala 143:13:freechips.rocketchip.system.DefaultRV32Config.fir@183562.10]
  wire  tlb__GEN_873; // @[TLB.scala 143:19:freechips.rocketchip.system.DefaultRV32Config.fir@183563.10]
  wire  tlb__GEN_874; // @[TLB.scala 379:40:freechips.rocketchip.system.DefaultRV32Config.fir@183524.8]
  wire  tlb__T_3753; // @[TLB.scala 383:24:freechips.rocketchip.system.DefaultRV32Config.fir@183572.4]
  wire [19:0] pma_checker_OptimizationBarrier_io_x_ppn; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@176907.4]
  wire  pma_checker_OptimizationBarrier_io_x_u; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@176907.4]
  wire  pma_checker_OptimizationBarrier_io_x_ae; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@176907.4]
  wire  pma_checker_OptimizationBarrier_io_x_sw; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@176907.4]
  wire  pma_checker_OptimizationBarrier_io_x_sx; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@176907.4]
  wire  pma_checker_OptimizationBarrier_io_x_sr; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@176907.4]
  wire  pma_checker_OptimizationBarrier_io_x_pw; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@176907.4]
  wire  pma_checker_OptimizationBarrier_io_x_px; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@176907.4]
  wire  pma_checker_OptimizationBarrier_io_x_pr; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@176907.4]
  wire  pma_checker_OptimizationBarrier_io_x_ppp; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@176907.4]
  wire  pma_checker_OptimizationBarrier_io_x_pal; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@176907.4]
  wire  pma_checker_OptimizationBarrier_io_x_paa; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@176907.4]
  wire  pma_checker_OptimizationBarrier_io_x_eff; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@176907.4]
  wire  pma_checker_OptimizationBarrier_io_x_c; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@176907.4]
  wire [19:0] pma_checker_OptimizationBarrier_io_y_ppn; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@176907.4]
  wire  pma_checker_OptimizationBarrier_io_y_u; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@176907.4]
  wire  pma_checker_OptimizationBarrier_io_y_ae; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@176907.4]
  wire  pma_checker_OptimizationBarrier_io_y_sw; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@176907.4]
  wire  pma_checker_OptimizationBarrier_io_y_sx; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@176907.4]
  wire  pma_checker_OptimizationBarrier_io_y_sr; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@176907.4]
  wire  pma_checker_OptimizationBarrier_io_y_pw; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@176907.4]
  wire  pma_checker_OptimizationBarrier_io_y_px; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@176907.4]
  wire  pma_checker_OptimizationBarrier_io_y_pr; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@176907.4]
  wire  pma_checker_OptimizationBarrier_io_y_ppp; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@176907.4]
  wire  pma_checker_OptimizationBarrier_io_y_pal; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@176907.4]
  wire  pma_checker_OptimizationBarrier_io_y_paa; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@176907.4]
  wire  pma_checker_OptimizationBarrier_io_y_eff; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@176907.4]
  wire  pma_checker_OptimizationBarrier_io_y_c; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@176907.4]
  wire [1:0] pma_checker_pmp_io_prv; // @[TLB.scala 190:19:freechips.rocketchip.system.DefaultRV32Config.fir@176928.4]
  wire  pma_checker_pmp_io_pmp_0_cfg_l; // @[TLB.scala 190:19:freechips.rocketchip.system.DefaultRV32Config.fir@176928.4]
  wire [1:0] pma_checker_pmp_io_pmp_0_cfg_a; // @[TLB.scala 190:19:freechips.rocketchip.system.DefaultRV32Config.fir@176928.4]
  wire  pma_checker_pmp_io_pmp_0_cfg_x; // @[TLB.scala 190:19:freechips.rocketchip.system.DefaultRV32Config.fir@176928.4]
  wire  pma_checker_pmp_io_pmp_0_cfg_w; // @[TLB.scala 190:19:freechips.rocketchip.system.DefaultRV32Config.fir@176928.4]
  wire  pma_checker_pmp_io_pmp_0_cfg_r; // @[TLB.scala 190:19:freechips.rocketchip.system.DefaultRV32Config.fir@176928.4]
  wire [29:0] pma_checker_pmp_io_pmp_0_addr; // @[TLB.scala 190:19:freechips.rocketchip.system.DefaultRV32Config.fir@176928.4]
  wire [31:0] pma_checker_pmp_io_pmp_0_mask; // @[TLB.scala 190:19:freechips.rocketchip.system.DefaultRV32Config.fir@176928.4]
  wire  pma_checker_pmp_io_pmp_1_cfg_l; // @[TLB.scala 190:19:freechips.rocketchip.system.DefaultRV32Config.fir@176928.4]
  wire [1:0] pma_checker_pmp_io_pmp_1_cfg_a; // @[TLB.scala 190:19:freechips.rocketchip.system.DefaultRV32Config.fir@176928.4]
  wire  pma_checker_pmp_io_pmp_1_cfg_x; // @[TLB.scala 190:19:freechips.rocketchip.system.DefaultRV32Config.fir@176928.4]
  wire  pma_checker_pmp_io_pmp_1_cfg_w; // @[TLB.scala 190:19:freechips.rocketchip.system.DefaultRV32Config.fir@176928.4]
  wire  pma_checker_pmp_io_pmp_1_cfg_r; // @[TLB.scala 190:19:freechips.rocketchip.system.DefaultRV32Config.fir@176928.4]
  wire [29:0] pma_checker_pmp_io_pmp_1_addr; // @[TLB.scala 190:19:freechips.rocketchip.system.DefaultRV32Config.fir@176928.4]
  wire [31:0] pma_checker_pmp_io_pmp_1_mask; // @[TLB.scala 190:19:freechips.rocketchip.system.DefaultRV32Config.fir@176928.4]
  wire  pma_checker_pmp_io_pmp_2_cfg_l; // @[TLB.scala 190:19:freechips.rocketchip.system.DefaultRV32Config.fir@176928.4]
  wire [1:0] pma_checker_pmp_io_pmp_2_cfg_a; // @[TLB.scala 190:19:freechips.rocketchip.system.DefaultRV32Config.fir@176928.4]
  wire  pma_checker_pmp_io_pmp_2_cfg_x; // @[TLB.scala 190:19:freechips.rocketchip.system.DefaultRV32Config.fir@176928.4]
  wire  pma_checker_pmp_io_pmp_2_cfg_w; // @[TLB.scala 190:19:freechips.rocketchip.system.DefaultRV32Config.fir@176928.4]
  wire  pma_checker_pmp_io_pmp_2_cfg_r; // @[TLB.scala 190:19:freechips.rocketchip.system.DefaultRV32Config.fir@176928.4]
  wire [29:0] pma_checker_pmp_io_pmp_2_addr; // @[TLB.scala 190:19:freechips.rocketchip.system.DefaultRV32Config.fir@176928.4]
  wire [31:0] pma_checker_pmp_io_pmp_2_mask; // @[TLB.scala 190:19:freechips.rocketchip.system.DefaultRV32Config.fir@176928.4]
  wire  pma_checker_pmp_io_pmp_3_cfg_l; // @[TLB.scala 190:19:freechips.rocketchip.system.DefaultRV32Config.fir@176928.4]
  wire [1:0] pma_checker_pmp_io_pmp_3_cfg_a; // @[TLB.scala 190:19:freechips.rocketchip.system.DefaultRV32Config.fir@176928.4]
  wire  pma_checker_pmp_io_pmp_3_cfg_x; // @[TLB.scala 190:19:freechips.rocketchip.system.DefaultRV32Config.fir@176928.4]
  wire  pma_checker_pmp_io_pmp_3_cfg_w; // @[TLB.scala 190:19:freechips.rocketchip.system.DefaultRV32Config.fir@176928.4]
  wire  pma_checker_pmp_io_pmp_3_cfg_r; // @[TLB.scala 190:19:freechips.rocketchip.system.DefaultRV32Config.fir@176928.4]
  wire [29:0] pma_checker_pmp_io_pmp_3_addr; // @[TLB.scala 190:19:freechips.rocketchip.system.DefaultRV32Config.fir@176928.4]
  wire [31:0] pma_checker_pmp_io_pmp_3_mask; // @[TLB.scala 190:19:freechips.rocketchip.system.DefaultRV32Config.fir@176928.4]
  wire  pma_checker_pmp_io_pmp_4_cfg_l; // @[TLB.scala 190:19:freechips.rocketchip.system.DefaultRV32Config.fir@176928.4]
  wire [1:0] pma_checker_pmp_io_pmp_4_cfg_a; // @[TLB.scala 190:19:freechips.rocketchip.system.DefaultRV32Config.fir@176928.4]
  wire  pma_checker_pmp_io_pmp_4_cfg_x; // @[TLB.scala 190:19:freechips.rocketchip.system.DefaultRV32Config.fir@176928.4]
  wire  pma_checker_pmp_io_pmp_4_cfg_w; // @[TLB.scala 190:19:freechips.rocketchip.system.DefaultRV32Config.fir@176928.4]
  wire  pma_checker_pmp_io_pmp_4_cfg_r; // @[TLB.scala 190:19:freechips.rocketchip.system.DefaultRV32Config.fir@176928.4]
  wire [29:0] pma_checker_pmp_io_pmp_4_addr; // @[TLB.scala 190:19:freechips.rocketchip.system.DefaultRV32Config.fir@176928.4]
  wire [31:0] pma_checker_pmp_io_pmp_4_mask; // @[TLB.scala 190:19:freechips.rocketchip.system.DefaultRV32Config.fir@176928.4]
  wire  pma_checker_pmp_io_pmp_5_cfg_l; // @[TLB.scala 190:19:freechips.rocketchip.system.DefaultRV32Config.fir@176928.4]
  wire [1:0] pma_checker_pmp_io_pmp_5_cfg_a; // @[TLB.scala 190:19:freechips.rocketchip.system.DefaultRV32Config.fir@176928.4]
  wire  pma_checker_pmp_io_pmp_5_cfg_x; // @[TLB.scala 190:19:freechips.rocketchip.system.DefaultRV32Config.fir@176928.4]
  wire  pma_checker_pmp_io_pmp_5_cfg_w; // @[TLB.scala 190:19:freechips.rocketchip.system.DefaultRV32Config.fir@176928.4]
  wire  pma_checker_pmp_io_pmp_5_cfg_r; // @[TLB.scala 190:19:freechips.rocketchip.system.DefaultRV32Config.fir@176928.4]
  wire [29:0] pma_checker_pmp_io_pmp_5_addr; // @[TLB.scala 190:19:freechips.rocketchip.system.DefaultRV32Config.fir@176928.4]
  wire [31:0] pma_checker_pmp_io_pmp_5_mask; // @[TLB.scala 190:19:freechips.rocketchip.system.DefaultRV32Config.fir@176928.4]
  wire  pma_checker_pmp_io_pmp_6_cfg_l; // @[TLB.scala 190:19:freechips.rocketchip.system.DefaultRV32Config.fir@176928.4]
  wire [1:0] pma_checker_pmp_io_pmp_6_cfg_a; // @[TLB.scala 190:19:freechips.rocketchip.system.DefaultRV32Config.fir@176928.4]
  wire  pma_checker_pmp_io_pmp_6_cfg_x; // @[TLB.scala 190:19:freechips.rocketchip.system.DefaultRV32Config.fir@176928.4]
  wire  pma_checker_pmp_io_pmp_6_cfg_w; // @[TLB.scala 190:19:freechips.rocketchip.system.DefaultRV32Config.fir@176928.4]
  wire  pma_checker_pmp_io_pmp_6_cfg_r; // @[TLB.scala 190:19:freechips.rocketchip.system.DefaultRV32Config.fir@176928.4]
  wire [29:0] pma_checker_pmp_io_pmp_6_addr; // @[TLB.scala 190:19:freechips.rocketchip.system.DefaultRV32Config.fir@176928.4]
  wire [31:0] pma_checker_pmp_io_pmp_6_mask; // @[TLB.scala 190:19:freechips.rocketchip.system.DefaultRV32Config.fir@176928.4]
  wire  pma_checker_pmp_io_pmp_7_cfg_l; // @[TLB.scala 190:19:freechips.rocketchip.system.DefaultRV32Config.fir@176928.4]
  wire [1:0] pma_checker_pmp_io_pmp_7_cfg_a; // @[TLB.scala 190:19:freechips.rocketchip.system.DefaultRV32Config.fir@176928.4]
  wire  pma_checker_pmp_io_pmp_7_cfg_x; // @[TLB.scala 190:19:freechips.rocketchip.system.DefaultRV32Config.fir@176928.4]
  wire  pma_checker_pmp_io_pmp_7_cfg_w; // @[TLB.scala 190:19:freechips.rocketchip.system.DefaultRV32Config.fir@176928.4]
  wire  pma_checker_pmp_io_pmp_7_cfg_r; // @[TLB.scala 190:19:freechips.rocketchip.system.DefaultRV32Config.fir@176928.4]
  wire [29:0] pma_checker_pmp_io_pmp_7_addr; // @[TLB.scala 190:19:freechips.rocketchip.system.DefaultRV32Config.fir@176928.4]
  wire [31:0] pma_checker_pmp_io_pmp_7_mask; // @[TLB.scala 190:19:freechips.rocketchip.system.DefaultRV32Config.fir@176928.4]
  wire [31:0] pma_checker_pmp_io_addr; // @[TLB.scala 190:19:freechips.rocketchip.system.DefaultRV32Config.fir@176928.4]
  wire  pma_checker_pmp_io_r; // @[TLB.scala 190:19:freechips.rocketchip.system.DefaultRV32Config.fir@176928.4]
  wire  pma_checker_pmp_io_w; // @[TLB.scala 190:19:freechips.rocketchip.system.DefaultRV32Config.fir@176928.4]
  wire  pma_checker_pmp_io_x; // @[TLB.scala 190:19:freechips.rocketchip.system.DefaultRV32Config.fir@176928.4]
  wire [19:0] pma_checker_OptimizationBarrier_1_io_x_ppn; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@177629.4]
  wire  pma_checker_OptimizationBarrier_1_io_x_u; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@177629.4]
  wire  pma_checker_OptimizationBarrier_1_io_x_ae; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@177629.4]
  wire  pma_checker_OptimizationBarrier_1_io_x_sw; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@177629.4]
  wire  pma_checker_OptimizationBarrier_1_io_x_sx; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@177629.4]
  wire  pma_checker_OptimizationBarrier_1_io_x_sr; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@177629.4]
  wire  pma_checker_OptimizationBarrier_1_io_x_pw; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@177629.4]
  wire  pma_checker_OptimizationBarrier_1_io_x_px; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@177629.4]
  wire  pma_checker_OptimizationBarrier_1_io_x_pr; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@177629.4]
  wire  pma_checker_OptimizationBarrier_1_io_x_ppp; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@177629.4]
  wire  pma_checker_OptimizationBarrier_1_io_x_pal; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@177629.4]
  wire  pma_checker_OptimizationBarrier_1_io_x_paa; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@177629.4]
  wire  pma_checker_OptimizationBarrier_1_io_x_eff; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@177629.4]
  wire  pma_checker_OptimizationBarrier_1_io_x_c; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@177629.4]
  wire [19:0] pma_checker_OptimizationBarrier_1_io_y_ppn; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@177629.4]
  wire  pma_checker_OptimizationBarrier_1_io_y_u; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@177629.4]
  wire  pma_checker_OptimizationBarrier_1_io_y_ae; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@177629.4]
  wire  pma_checker_OptimizationBarrier_1_io_y_sw; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@177629.4]
  wire  pma_checker_OptimizationBarrier_1_io_y_sx; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@177629.4]
  wire  pma_checker_OptimizationBarrier_1_io_y_sr; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@177629.4]
  wire  pma_checker_OptimizationBarrier_1_io_y_pw; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@177629.4]
  wire  pma_checker_OptimizationBarrier_1_io_y_px; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@177629.4]
  wire  pma_checker_OptimizationBarrier_1_io_y_pr; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@177629.4]
  wire  pma_checker_OptimizationBarrier_1_io_y_ppp; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@177629.4]
  wire  pma_checker_OptimizationBarrier_1_io_y_pal; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@177629.4]
  wire  pma_checker_OptimizationBarrier_1_io_y_paa; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@177629.4]
  wire  pma_checker_OptimizationBarrier_1_io_y_eff; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@177629.4]
  wire  pma_checker_OptimizationBarrier_1_io_y_c; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@177629.4]
  wire [19:0] pma_checker_OptimizationBarrier_2_io_x_ppn; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@177672.4]
  wire  pma_checker_OptimizationBarrier_2_io_x_u; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@177672.4]
  wire  pma_checker_OptimizationBarrier_2_io_x_ae; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@177672.4]
  wire  pma_checker_OptimizationBarrier_2_io_x_sw; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@177672.4]
  wire  pma_checker_OptimizationBarrier_2_io_x_sx; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@177672.4]
  wire  pma_checker_OptimizationBarrier_2_io_x_sr; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@177672.4]
  wire  pma_checker_OptimizationBarrier_2_io_x_pw; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@177672.4]
  wire  pma_checker_OptimizationBarrier_2_io_x_px; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@177672.4]
  wire  pma_checker_OptimizationBarrier_2_io_x_pr; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@177672.4]
  wire  pma_checker_OptimizationBarrier_2_io_x_ppp; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@177672.4]
  wire  pma_checker_OptimizationBarrier_2_io_x_pal; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@177672.4]
  wire  pma_checker_OptimizationBarrier_2_io_x_paa; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@177672.4]
  wire  pma_checker_OptimizationBarrier_2_io_x_eff; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@177672.4]
  wire  pma_checker_OptimizationBarrier_2_io_x_c; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@177672.4]
  wire [19:0] pma_checker_OptimizationBarrier_2_io_y_ppn; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@177672.4]
  wire  pma_checker_OptimizationBarrier_2_io_y_u; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@177672.4]
  wire  pma_checker_OptimizationBarrier_2_io_y_ae; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@177672.4]
  wire  pma_checker_OptimizationBarrier_2_io_y_sw; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@177672.4]
  wire  pma_checker_OptimizationBarrier_2_io_y_sx; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@177672.4]
  wire  pma_checker_OptimizationBarrier_2_io_y_sr; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@177672.4]
  wire  pma_checker_OptimizationBarrier_2_io_y_pw; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@177672.4]
  wire  pma_checker_OptimizationBarrier_2_io_y_px; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@177672.4]
  wire  pma_checker_OptimizationBarrier_2_io_y_pr; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@177672.4]
  wire  pma_checker_OptimizationBarrier_2_io_y_ppp; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@177672.4]
  wire  pma_checker_OptimizationBarrier_2_io_y_pal; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@177672.4]
  wire  pma_checker_OptimizationBarrier_2_io_y_paa; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@177672.4]
  wire  pma_checker_OptimizationBarrier_2_io_y_eff; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@177672.4]
  wire  pma_checker_OptimizationBarrier_2_io_y_c; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@177672.4]
  wire [19:0] pma_checker_OptimizationBarrier_3_io_x_ppn; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@177715.4]
  wire  pma_checker_OptimizationBarrier_3_io_x_u; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@177715.4]
  wire  pma_checker_OptimizationBarrier_3_io_x_ae; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@177715.4]
  wire  pma_checker_OptimizationBarrier_3_io_x_sw; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@177715.4]
  wire  pma_checker_OptimizationBarrier_3_io_x_sx; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@177715.4]
  wire  pma_checker_OptimizationBarrier_3_io_x_sr; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@177715.4]
  wire  pma_checker_OptimizationBarrier_3_io_x_pw; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@177715.4]
  wire  pma_checker_OptimizationBarrier_3_io_x_px; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@177715.4]
  wire  pma_checker_OptimizationBarrier_3_io_x_pr; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@177715.4]
  wire  pma_checker_OptimizationBarrier_3_io_x_ppp; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@177715.4]
  wire  pma_checker_OptimizationBarrier_3_io_x_pal; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@177715.4]
  wire  pma_checker_OptimizationBarrier_3_io_x_paa; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@177715.4]
  wire  pma_checker_OptimizationBarrier_3_io_x_eff; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@177715.4]
  wire  pma_checker_OptimizationBarrier_3_io_x_c; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@177715.4]
  wire [19:0] pma_checker_OptimizationBarrier_3_io_y_ppn; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@177715.4]
  wire  pma_checker_OptimizationBarrier_3_io_y_u; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@177715.4]
  wire  pma_checker_OptimizationBarrier_3_io_y_ae; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@177715.4]
  wire  pma_checker_OptimizationBarrier_3_io_y_sw; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@177715.4]
  wire  pma_checker_OptimizationBarrier_3_io_y_sx; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@177715.4]
  wire  pma_checker_OptimizationBarrier_3_io_y_sr; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@177715.4]
  wire  pma_checker_OptimizationBarrier_3_io_y_pw; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@177715.4]
  wire  pma_checker_OptimizationBarrier_3_io_y_px; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@177715.4]
  wire  pma_checker_OptimizationBarrier_3_io_y_pr; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@177715.4]
  wire  pma_checker_OptimizationBarrier_3_io_y_ppp; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@177715.4]
  wire  pma_checker_OptimizationBarrier_3_io_y_pal; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@177715.4]
  wire  pma_checker_OptimizationBarrier_3_io_y_paa; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@177715.4]
  wire  pma_checker_OptimizationBarrier_3_io_y_eff; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@177715.4]
  wire  pma_checker_OptimizationBarrier_3_io_y_c; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@177715.4]
  wire [19:0] pma_checker_OptimizationBarrier_4_io_x_ppn; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@177758.4]
  wire  pma_checker_OptimizationBarrier_4_io_x_u; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@177758.4]
  wire  pma_checker_OptimizationBarrier_4_io_x_ae; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@177758.4]
  wire  pma_checker_OptimizationBarrier_4_io_x_sw; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@177758.4]
  wire  pma_checker_OptimizationBarrier_4_io_x_sx; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@177758.4]
  wire  pma_checker_OptimizationBarrier_4_io_x_sr; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@177758.4]
  wire  pma_checker_OptimizationBarrier_4_io_x_pw; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@177758.4]
  wire  pma_checker_OptimizationBarrier_4_io_x_px; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@177758.4]
  wire  pma_checker_OptimizationBarrier_4_io_x_pr; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@177758.4]
  wire  pma_checker_OptimizationBarrier_4_io_x_ppp; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@177758.4]
  wire  pma_checker_OptimizationBarrier_4_io_x_pal; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@177758.4]
  wire  pma_checker_OptimizationBarrier_4_io_x_paa; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@177758.4]
  wire  pma_checker_OptimizationBarrier_4_io_x_eff; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@177758.4]
  wire  pma_checker_OptimizationBarrier_4_io_x_c; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@177758.4]
  wire [19:0] pma_checker_OptimizationBarrier_4_io_y_ppn; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@177758.4]
  wire  pma_checker_OptimizationBarrier_4_io_y_u; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@177758.4]
  wire  pma_checker_OptimizationBarrier_4_io_y_ae; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@177758.4]
  wire  pma_checker_OptimizationBarrier_4_io_y_sw; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@177758.4]
  wire  pma_checker_OptimizationBarrier_4_io_y_sx; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@177758.4]
  wire  pma_checker_OptimizationBarrier_4_io_y_sr; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@177758.4]
  wire  pma_checker_OptimizationBarrier_4_io_y_pw; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@177758.4]
  wire  pma_checker_OptimizationBarrier_4_io_y_px; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@177758.4]
  wire  pma_checker_OptimizationBarrier_4_io_y_pr; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@177758.4]
  wire  pma_checker_OptimizationBarrier_4_io_y_ppp; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@177758.4]
  wire  pma_checker_OptimizationBarrier_4_io_y_pal; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@177758.4]
  wire  pma_checker_OptimizationBarrier_4_io_y_paa; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@177758.4]
  wire  pma_checker_OptimizationBarrier_4_io_y_eff; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@177758.4]
  wire  pma_checker_OptimizationBarrier_4_io_y_c; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@177758.4]
  wire [19:0] pma_checker_OptimizationBarrier_5_io_x_ppn; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@177801.4]
  wire  pma_checker_OptimizationBarrier_5_io_x_u; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@177801.4]
  wire  pma_checker_OptimizationBarrier_5_io_x_ae; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@177801.4]
  wire  pma_checker_OptimizationBarrier_5_io_x_sw; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@177801.4]
  wire  pma_checker_OptimizationBarrier_5_io_x_sx; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@177801.4]
  wire  pma_checker_OptimizationBarrier_5_io_x_sr; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@177801.4]
  wire  pma_checker_OptimizationBarrier_5_io_x_pw; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@177801.4]
  wire  pma_checker_OptimizationBarrier_5_io_x_px; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@177801.4]
  wire  pma_checker_OptimizationBarrier_5_io_x_pr; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@177801.4]
  wire  pma_checker_OptimizationBarrier_5_io_x_ppp; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@177801.4]
  wire  pma_checker_OptimizationBarrier_5_io_x_pal; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@177801.4]
  wire  pma_checker_OptimizationBarrier_5_io_x_paa; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@177801.4]
  wire  pma_checker_OptimizationBarrier_5_io_x_eff; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@177801.4]
  wire  pma_checker_OptimizationBarrier_5_io_x_c; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@177801.4]
  wire [19:0] pma_checker_OptimizationBarrier_5_io_y_ppn; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@177801.4]
  wire  pma_checker_OptimizationBarrier_5_io_y_u; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@177801.4]
  wire  pma_checker_OptimizationBarrier_5_io_y_ae; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@177801.4]
  wire  pma_checker_OptimizationBarrier_5_io_y_sw; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@177801.4]
  wire  pma_checker_OptimizationBarrier_5_io_y_sx; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@177801.4]
  wire  pma_checker_OptimizationBarrier_5_io_y_sr; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@177801.4]
  wire  pma_checker_OptimizationBarrier_5_io_y_pw; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@177801.4]
  wire  pma_checker_OptimizationBarrier_5_io_y_px; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@177801.4]
  wire  pma_checker_OptimizationBarrier_5_io_y_pr; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@177801.4]
  wire  pma_checker_OptimizationBarrier_5_io_y_ppp; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@177801.4]
  wire  pma_checker_OptimizationBarrier_5_io_y_pal; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@177801.4]
  wire  pma_checker_OptimizationBarrier_5_io_y_paa; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@177801.4]
  wire  pma_checker_OptimizationBarrier_5_io_y_eff; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@177801.4]
  wire  pma_checker_OptimizationBarrier_5_io_y_c; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@177801.4]
  wire [19:0] pma_checker_OptimizationBarrier_6_io_x_ppn; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@177844.4]
  wire  pma_checker_OptimizationBarrier_6_io_x_u; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@177844.4]
  wire  pma_checker_OptimizationBarrier_6_io_x_ae; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@177844.4]
  wire  pma_checker_OptimizationBarrier_6_io_x_sw; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@177844.4]
  wire  pma_checker_OptimizationBarrier_6_io_x_sx; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@177844.4]
  wire  pma_checker_OptimizationBarrier_6_io_x_sr; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@177844.4]
  wire  pma_checker_OptimizationBarrier_6_io_x_pw; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@177844.4]
  wire  pma_checker_OptimizationBarrier_6_io_x_px; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@177844.4]
  wire  pma_checker_OptimizationBarrier_6_io_x_pr; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@177844.4]
  wire  pma_checker_OptimizationBarrier_6_io_x_ppp; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@177844.4]
  wire  pma_checker_OptimizationBarrier_6_io_x_pal; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@177844.4]
  wire  pma_checker_OptimizationBarrier_6_io_x_paa; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@177844.4]
  wire  pma_checker_OptimizationBarrier_6_io_x_eff; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@177844.4]
  wire  pma_checker_OptimizationBarrier_6_io_x_c; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@177844.4]
  wire [19:0] pma_checker_OptimizationBarrier_6_io_y_ppn; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@177844.4]
  wire  pma_checker_OptimizationBarrier_6_io_y_u; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@177844.4]
  wire  pma_checker_OptimizationBarrier_6_io_y_ae; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@177844.4]
  wire  pma_checker_OptimizationBarrier_6_io_y_sw; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@177844.4]
  wire  pma_checker_OptimizationBarrier_6_io_y_sx; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@177844.4]
  wire  pma_checker_OptimizationBarrier_6_io_y_sr; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@177844.4]
  wire  pma_checker_OptimizationBarrier_6_io_y_pw; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@177844.4]
  wire  pma_checker_OptimizationBarrier_6_io_y_px; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@177844.4]
  wire  pma_checker_OptimizationBarrier_6_io_y_pr; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@177844.4]
  wire  pma_checker_OptimizationBarrier_6_io_y_ppp; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@177844.4]
  wire  pma_checker_OptimizationBarrier_6_io_y_pal; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@177844.4]
  wire  pma_checker_OptimizationBarrier_6_io_y_paa; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@177844.4]
  wire  pma_checker_OptimizationBarrier_6_io_y_eff; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@177844.4]
  wire  pma_checker_OptimizationBarrier_6_io_y_c; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@177844.4]
  wire [19:0] pma_checker_OptimizationBarrier_7_io_x_ppn; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@177887.4]
  wire  pma_checker_OptimizationBarrier_7_io_x_u; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@177887.4]
  wire  pma_checker_OptimizationBarrier_7_io_x_ae; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@177887.4]
  wire  pma_checker_OptimizationBarrier_7_io_x_sw; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@177887.4]
  wire  pma_checker_OptimizationBarrier_7_io_x_sx; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@177887.4]
  wire  pma_checker_OptimizationBarrier_7_io_x_sr; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@177887.4]
  wire  pma_checker_OptimizationBarrier_7_io_x_pw; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@177887.4]
  wire  pma_checker_OptimizationBarrier_7_io_x_px; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@177887.4]
  wire  pma_checker_OptimizationBarrier_7_io_x_pr; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@177887.4]
  wire  pma_checker_OptimizationBarrier_7_io_x_ppp; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@177887.4]
  wire  pma_checker_OptimizationBarrier_7_io_x_pal; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@177887.4]
  wire  pma_checker_OptimizationBarrier_7_io_x_paa; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@177887.4]
  wire  pma_checker_OptimizationBarrier_7_io_x_eff; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@177887.4]
  wire  pma_checker_OptimizationBarrier_7_io_x_c; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@177887.4]
  wire [19:0] pma_checker_OptimizationBarrier_7_io_y_ppn; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@177887.4]
  wire  pma_checker_OptimizationBarrier_7_io_y_u; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@177887.4]
  wire  pma_checker_OptimizationBarrier_7_io_y_ae; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@177887.4]
  wire  pma_checker_OptimizationBarrier_7_io_y_sw; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@177887.4]
  wire  pma_checker_OptimizationBarrier_7_io_y_sx; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@177887.4]
  wire  pma_checker_OptimizationBarrier_7_io_y_sr; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@177887.4]
  wire  pma_checker_OptimizationBarrier_7_io_y_pw; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@177887.4]
  wire  pma_checker_OptimizationBarrier_7_io_y_px; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@177887.4]
  wire  pma_checker_OptimizationBarrier_7_io_y_pr; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@177887.4]
  wire  pma_checker_OptimizationBarrier_7_io_y_ppp; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@177887.4]
  wire  pma_checker_OptimizationBarrier_7_io_y_pal; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@177887.4]
  wire  pma_checker_OptimizationBarrier_7_io_y_paa; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@177887.4]
  wire  pma_checker_OptimizationBarrier_7_io_y_eff; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@177887.4]
  wire  pma_checker_OptimizationBarrier_7_io_y_c; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@177887.4]
  wire [19:0] pma_checker_OptimizationBarrier_8_io_x_ppn; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@177930.4]
  wire  pma_checker_OptimizationBarrier_8_io_x_u; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@177930.4]
  wire  pma_checker_OptimizationBarrier_8_io_x_ae; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@177930.4]
  wire  pma_checker_OptimizationBarrier_8_io_x_sw; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@177930.4]
  wire  pma_checker_OptimizationBarrier_8_io_x_sx; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@177930.4]
  wire  pma_checker_OptimizationBarrier_8_io_x_sr; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@177930.4]
  wire  pma_checker_OptimizationBarrier_8_io_x_pw; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@177930.4]
  wire  pma_checker_OptimizationBarrier_8_io_x_px; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@177930.4]
  wire  pma_checker_OptimizationBarrier_8_io_x_pr; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@177930.4]
  wire  pma_checker_OptimizationBarrier_8_io_x_ppp; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@177930.4]
  wire  pma_checker_OptimizationBarrier_8_io_x_pal; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@177930.4]
  wire  pma_checker_OptimizationBarrier_8_io_x_paa; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@177930.4]
  wire  pma_checker_OptimizationBarrier_8_io_x_eff; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@177930.4]
  wire  pma_checker_OptimizationBarrier_8_io_x_c; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@177930.4]
  wire [19:0] pma_checker_OptimizationBarrier_8_io_y_ppn; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@177930.4]
  wire  pma_checker_OptimizationBarrier_8_io_y_u; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@177930.4]
  wire  pma_checker_OptimizationBarrier_8_io_y_ae; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@177930.4]
  wire  pma_checker_OptimizationBarrier_8_io_y_sw; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@177930.4]
  wire  pma_checker_OptimizationBarrier_8_io_y_sx; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@177930.4]
  wire  pma_checker_OptimizationBarrier_8_io_y_sr; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@177930.4]
  wire  pma_checker_OptimizationBarrier_8_io_y_pw; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@177930.4]
  wire  pma_checker_OptimizationBarrier_8_io_y_px; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@177930.4]
  wire  pma_checker_OptimizationBarrier_8_io_y_pr; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@177930.4]
  wire  pma_checker_OptimizationBarrier_8_io_y_ppp; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@177930.4]
  wire  pma_checker_OptimizationBarrier_8_io_y_pal; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@177930.4]
  wire  pma_checker_OptimizationBarrier_8_io_y_paa; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@177930.4]
  wire  pma_checker_OptimizationBarrier_8_io_y_eff; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@177930.4]
  wire  pma_checker_OptimizationBarrier_8_io_y_c; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@177930.4]
  wire [19:0] pma_checker_OptimizationBarrier_9_io_x_ppn; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@177972.4]
  wire  pma_checker_OptimizationBarrier_9_io_x_u; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@177972.4]
  wire  pma_checker_OptimizationBarrier_9_io_x_ae; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@177972.4]
  wire  pma_checker_OptimizationBarrier_9_io_x_sw; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@177972.4]
  wire  pma_checker_OptimizationBarrier_9_io_x_sx; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@177972.4]
  wire  pma_checker_OptimizationBarrier_9_io_x_sr; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@177972.4]
  wire  pma_checker_OptimizationBarrier_9_io_x_pw; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@177972.4]
  wire  pma_checker_OptimizationBarrier_9_io_x_px; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@177972.4]
  wire  pma_checker_OptimizationBarrier_9_io_x_pr; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@177972.4]
  wire  pma_checker_OptimizationBarrier_9_io_x_ppp; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@177972.4]
  wire  pma_checker_OptimizationBarrier_9_io_x_pal; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@177972.4]
  wire  pma_checker_OptimizationBarrier_9_io_x_paa; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@177972.4]
  wire  pma_checker_OptimizationBarrier_9_io_x_eff; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@177972.4]
  wire  pma_checker_OptimizationBarrier_9_io_x_c; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@177972.4]
  wire [19:0] pma_checker_OptimizationBarrier_9_io_y_ppn; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@177972.4]
  wire  pma_checker_OptimizationBarrier_9_io_y_u; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@177972.4]
  wire  pma_checker_OptimizationBarrier_9_io_y_ae; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@177972.4]
  wire  pma_checker_OptimizationBarrier_9_io_y_sw; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@177972.4]
  wire  pma_checker_OptimizationBarrier_9_io_y_sx; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@177972.4]
  wire  pma_checker_OptimizationBarrier_9_io_y_sr; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@177972.4]
  wire  pma_checker_OptimizationBarrier_9_io_y_pw; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@177972.4]
  wire  pma_checker_OptimizationBarrier_9_io_y_px; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@177972.4]
  wire  pma_checker_OptimizationBarrier_9_io_y_pr; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@177972.4]
  wire  pma_checker_OptimizationBarrier_9_io_y_ppp; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@177972.4]
  wire  pma_checker_OptimizationBarrier_9_io_y_pal; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@177972.4]
  wire  pma_checker_OptimizationBarrier_9_io_y_paa; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@177972.4]
  wire  pma_checker_OptimizationBarrier_9_io_y_eff; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@177972.4]
  wire  pma_checker_OptimizationBarrier_9_io_y_c; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@177972.4]
  wire [19:0] pma_checker_OptimizationBarrier_10_io_x_ppn; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178021.4]
  wire  pma_checker_OptimizationBarrier_10_io_x_u; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178021.4]
  wire  pma_checker_OptimizationBarrier_10_io_x_ae; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178021.4]
  wire  pma_checker_OptimizationBarrier_10_io_x_sw; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178021.4]
  wire  pma_checker_OptimizationBarrier_10_io_x_sx; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178021.4]
  wire  pma_checker_OptimizationBarrier_10_io_x_sr; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178021.4]
  wire  pma_checker_OptimizationBarrier_10_io_x_pw; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178021.4]
  wire  pma_checker_OptimizationBarrier_10_io_x_px; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178021.4]
  wire  pma_checker_OptimizationBarrier_10_io_x_pr; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178021.4]
  wire  pma_checker_OptimizationBarrier_10_io_x_ppp; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178021.4]
  wire  pma_checker_OptimizationBarrier_10_io_x_pal; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178021.4]
  wire  pma_checker_OptimizationBarrier_10_io_x_paa; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178021.4]
  wire  pma_checker_OptimizationBarrier_10_io_x_eff; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178021.4]
  wire  pma_checker_OptimizationBarrier_10_io_x_c; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178021.4]
  wire [19:0] pma_checker_OptimizationBarrier_10_io_y_ppn; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178021.4]
  wire  pma_checker_OptimizationBarrier_10_io_y_u; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178021.4]
  wire  pma_checker_OptimizationBarrier_10_io_y_ae; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178021.4]
  wire  pma_checker_OptimizationBarrier_10_io_y_sw; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178021.4]
  wire  pma_checker_OptimizationBarrier_10_io_y_sx; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178021.4]
  wire  pma_checker_OptimizationBarrier_10_io_y_sr; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178021.4]
  wire  pma_checker_OptimizationBarrier_10_io_y_pw; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178021.4]
  wire  pma_checker_OptimizationBarrier_10_io_y_px; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178021.4]
  wire  pma_checker_OptimizationBarrier_10_io_y_pr; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178021.4]
  wire  pma_checker_OptimizationBarrier_10_io_y_ppp; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178021.4]
  wire  pma_checker_OptimizationBarrier_10_io_y_pal; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178021.4]
  wire  pma_checker_OptimizationBarrier_10_io_y_paa; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178021.4]
  wire  pma_checker_OptimizationBarrier_10_io_y_eff; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178021.4]
  wire  pma_checker_OptimizationBarrier_10_io_y_c; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178021.4]
  wire [19:0] pma_checker_OptimizationBarrier_11_io_x_ppn; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178070.4]
  wire  pma_checker_OptimizationBarrier_11_io_x_u; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178070.4]
  wire  pma_checker_OptimizationBarrier_11_io_x_ae; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178070.4]
  wire  pma_checker_OptimizationBarrier_11_io_x_sw; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178070.4]
  wire  pma_checker_OptimizationBarrier_11_io_x_sx; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178070.4]
  wire  pma_checker_OptimizationBarrier_11_io_x_sr; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178070.4]
  wire  pma_checker_OptimizationBarrier_11_io_x_pw; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178070.4]
  wire  pma_checker_OptimizationBarrier_11_io_x_px; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178070.4]
  wire  pma_checker_OptimizationBarrier_11_io_x_pr; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178070.4]
  wire  pma_checker_OptimizationBarrier_11_io_x_ppp; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178070.4]
  wire  pma_checker_OptimizationBarrier_11_io_x_pal; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178070.4]
  wire  pma_checker_OptimizationBarrier_11_io_x_paa; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178070.4]
  wire  pma_checker_OptimizationBarrier_11_io_x_eff; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178070.4]
  wire  pma_checker_OptimizationBarrier_11_io_x_c; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178070.4]
  wire [19:0] pma_checker_OptimizationBarrier_11_io_y_ppn; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178070.4]
  wire  pma_checker_OptimizationBarrier_11_io_y_u; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178070.4]
  wire  pma_checker_OptimizationBarrier_11_io_y_ae; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178070.4]
  wire  pma_checker_OptimizationBarrier_11_io_y_sw; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178070.4]
  wire  pma_checker_OptimizationBarrier_11_io_y_sx; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178070.4]
  wire  pma_checker_OptimizationBarrier_11_io_y_sr; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178070.4]
  wire  pma_checker_OptimizationBarrier_11_io_y_pw; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178070.4]
  wire  pma_checker_OptimizationBarrier_11_io_y_px; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178070.4]
  wire  pma_checker_OptimizationBarrier_11_io_y_pr; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178070.4]
  wire  pma_checker_OptimizationBarrier_11_io_y_ppp; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178070.4]
  wire  pma_checker_OptimizationBarrier_11_io_y_pal; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178070.4]
  wire  pma_checker_OptimizationBarrier_11_io_y_paa; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178070.4]
  wire  pma_checker_OptimizationBarrier_11_io_y_eff; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178070.4]
  wire  pma_checker_OptimizationBarrier_11_io_y_c; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178070.4]
  wire [19:0] pma_checker_OptimizationBarrier_12_io_x_ppn; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178119.4]
  wire  pma_checker_OptimizationBarrier_12_io_x_u; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178119.4]
  wire  pma_checker_OptimizationBarrier_12_io_x_ae; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178119.4]
  wire  pma_checker_OptimizationBarrier_12_io_x_sw; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178119.4]
  wire  pma_checker_OptimizationBarrier_12_io_x_sx; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178119.4]
  wire  pma_checker_OptimizationBarrier_12_io_x_sr; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178119.4]
  wire  pma_checker_OptimizationBarrier_12_io_x_pw; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178119.4]
  wire  pma_checker_OptimizationBarrier_12_io_x_px; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178119.4]
  wire  pma_checker_OptimizationBarrier_12_io_x_pr; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178119.4]
  wire  pma_checker_OptimizationBarrier_12_io_x_ppp; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178119.4]
  wire  pma_checker_OptimizationBarrier_12_io_x_pal; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178119.4]
  wire  pma_checker_OptimizationBarrier_12_io_x_paa; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178119.4]
  wire  pma_checker_OptimizationBarrier_12_io_x_eff; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178119.4]
  wire  pma_checker_OptimizationBarrier_12_io_x_c; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178119.4]
  wire [19:0] pma_checker_OptimizationBarrier_12_io_y_ppn; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178119.4]
  wire  pma_checker_OptimizationBarrier_12_io_y_u; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178119.4]
  wire  pma_checker_OptimizationBarrier_12_io_y_ae; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178119.4]
  wire  pma_checker_OptimizationBarrier_12_io_y_sw; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178119.4]
  wire  pma_checker_OptimizationBarrier_12_io_y_sx; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178119.4]
  wire  pma_checker_OptimizationBarrier_12_io_y_sr; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178119.4]
  wire  pma_checker_OptimizationBarrier_12_io_y_pw; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178119.4]
  wire  pma_checker_OptimizationBarrier_12_io_y_px; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178119.4]
  wire  pma_checker_OptimizationBarrier_12_io_y_pr; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178119.4]
  wire  pma_checker_OptimizationBarrier_12_io_y_ppp; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178119.4]
  wire  pma_checker_OptimizationBarrier_12_io_y_pal; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178119.4]
  wire  pma_checker_OptimizationBarrier_12_io_y_paa; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178119.4]
  wire  pma_checker_OptimizationBarrier_12_io_y_eff; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178119.4]
  wire  pma_checker_OptimizationBarrier_12_io_y_c; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178119.4]
  wire [19:0] pma_checker_OptimizationBarrier_13_io_x_ppn; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178168.4]
  wire  pma_checker_OptimizationBarrier_13_io_x_u; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178168.4]
  wire  pma_checker_OptimizationBarrier_13_io_x_ae; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178168.4]
  wire  pma_checker_OptimizationBarrier_13_io_x_sw; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178168.4]
  wire  pma_checker_OptimizationBarrier_13_io_x_sx; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178168.4]
  wire  pma_checker_OptimizationBarrier_13_io_x_sr; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178168.4]
  wire  pma_checker_OptimizationBarrier_13_io_x_pw; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178168.4]
  wire  pma_checker_OptimizationBarrier_13_io_x_px; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178168.4]
  wire  pma_checker_OptimizationBarrier_13_io_x_pr; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178168.4]
  wire  pma_checker_OptimizationBarrier_13_io_x_ppp; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178168.4]
  wire  pma_checker_OptimizationBarrier_13_io_x_pal; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178168.4]
  wire  pma_checker_OptimizationBarrier_13_io_x_paa; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178168.4]
  wire  pma_checker_OptimizationBarrier_13_io_x_eff; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178168.4]
  wire  pma_checker_OptimizationBarrier_13_io_x_c; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178168.4]
  wire [19:0] pma_checker_OptimizationBarrier_13_io_y_ppn; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178168.4]
  wire  pma_checker_OptimizationBarrier_13_io_y_u; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178168.4]
  wire  pma_checker_OptimizationBarrier_13_io_y_ae; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178168.4]
  wire  pma_checker_OptimizationBarrier_13_io_y_sw; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178168.4]
  wire  pma_checker_OptimizationBarrier_13_io_y_sx; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178168.4]
  wire  pma_checker_OptimizationBarrier_13_io_y_sr; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178168.4]
  wire  pma_checker_OptimizationBarrier_13_io_y_pw; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178168.4]
  wire  pma_checker_OptimizationBarrier_13_io_y_px; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178168.4]
  wire  pma_checker_OptimizationBarrier_13_io_y_pr; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178168.4]
  wire  pma_checker_OptimizationBarrier_13_io_y_ppp; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178168.4]
  wire  pma_checker_OptimizationBarrier_13_io_y_pal; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178168.4]
  wire  pma_checker_OptimizationBarrier_13_io_y_paa; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178168.4]
  wire  pma_checker_OptimizationBarrier_13_io_y_eff; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178168.4]
  wire  pma_checker_OptimizationBarrier_13_io_y_c; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178168.4]
  wire [19:0] pma_checker_OptimizationBarrier_14_io_x_ppn; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178649.4]
  wire  pma_checker_OptimizationBarrier_14_io_x_u; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178649.4]
  wire  pma_checker_OptimizationBarrier_14_io_x_ae; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178649.4]
  wire  pma_checker_OptimizationBarrier_14_io_x_sw; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178649.4]
  wire  pma_checker_OptimizationBarrier_14_io_x_sx; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178649.4]
  wire  pma_checker_OptimizationBarrier_14_io_x_sr; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178649.4]
  wire  pma_checker_OptimizationBarrier_14_io_x_pw; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178649.4]
  wire  pma_checker_OptimizationBarrier_14_io_x_px; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178649.4]
  wire  pma_checker_OptimizationBarrier_14_io_x_pr; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178649.4]
  wire  pma_checker_OptimizationBarrier_14_io_x_ppp; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178649.4]
  wire  pma_checker_OptimizationBarrier_14_io_x_pal; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178649.4]
  wire  pma_checker_OptimizationBarrier_14_io_x_paa; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178649.4]
  wire  pma_checker_OptimizationBarrier_14_io_x_eff; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178649.4]
  wire  pma_checker_OptimizationBarrier_14_io_x_c; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178649.4]
  wire [19:0] pma_checker_OptimizationBarrier_14_io_y_ppn; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178649.4]
  wire  pma_checker_OptimizationBarrier_14_io_y_u; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178649.4]
  wire  pma_checker_OptimizationBarrier_14_io_y_ae; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178649.4]
  wire  pma_checker_OptimizationBarrier_14_io_y_sw; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178649.4]
  wire  pma_checker_OptimizationBarrier_14_io_y_sx; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178649.4]
  wire  pma_checker_OptimizationBarrier_14_io_y_sr; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178649.4]
  wire  pma_checker_OptimizationBarrier_14_io_y_pw; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178649.4]
  wire  pma_checker_OptimizationBarrier_14_io_y_px; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178649.4]
  wire  pma_checker_OptimizationBarrier_14_io_y_pr; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178649.4]
  wire  pma_checker_OptimizationBarrier_14_io_y_ppp; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178649.4]
  wire  pma_checker_OptimizationBarrier_14_io_y_pal; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178649.4]
  wire  pma_checker_OptimizationBarrier_14_io_y_paa; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178649.4]
  wire  pma_checker_OptimizationBarrier_14_io_y_eff; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178649.4]
  wire  pma_checker_OptimizationBarrier_14_io_y_c; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178649.4]
  wire [19:0] pma_checker_OptimizationBarrier_15_io_x_ppn; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178692.4]
  wire  pma_checker_OptimizationBarrier_15_io_x_u; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178692.4]
  wire  pma_checker_OptimizationBarrier_15_io_x_ae; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178692.4]
  wire  pma_checker_OptimizationBarrier_15_io_x_sw; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178692.4]
  wire  pma_checker_OptimizationBarrier_15_io_x_sx; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178692.4]
  wire  pma_checker_OptimizationBarrier_15_io_x_sr; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178692.4]
  wire  pma_checker_OptimizationBarrier_15_io_x_pw; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178692.4]
  wire  pma_checker_OptimizationBarrier_15_io_x_px; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178692.4]
  wire  pma_checker_OptimizationBarrier_15_io_x_pr; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178692.4]
  wire  pma_checker_OptimizationBarrier_15_io_x_ppp; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178692.4]
  wire  pma_checker_OptimizationBarrier_15_io_x_pal; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178692.4]
  wire  pma_checker_OptimizationBarrier_15_io_x_paa; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178692.4]
  wire  pma_checker_OptimizationBarrier_15_io_x_eff; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178692.4]
  wire  pma_checker_OptimizationBarrier_15_io_x_c; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178692.4]
  wire [19:0] pma_checker_OptimizationBarrier_15_io_y_ppn; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178692.4]
  wire  pma_checker_OptimizationBarrier_15_io_y_u; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178692.4]
  wire  pma_checker_OptimizationBarrier_15_io_y_ae; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178692.4]
  wire  pma_checker_OptimizationBarrier_15_io_y_sw; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178692.4]
  wire  pma_checker_OptimizationBarrier_15_io_y_sx; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178692.4]
  wire  pma_checker_OptimizationBarrier_15_io_y_sr; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178692.4]
  wire  pma_checker_OptimizationBarrier_15_io_y_pw; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178692.4]
  wire  pma_checker_OptimizationBarrier_15_io_y_px; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178692.4]
  wire  pma_checker_OptimizationBarrier_15_io_y_pr; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178692.4]
  wire  pma_checker_OptimizationBarrier_15_io_y_ppp; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178692.4]
  wire  pma_checker_OptimizationBarrier_15_io_y_pal; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178692.4]
  wire  pma_checker_OptimizationBarrier_15_io_y_paa; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178692.4]
  wire  pma_checker_OptimizationBarrier_15_io_y_eff; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178692.4]
  wire  pma_checker_OptimizationBarrier_15_io_y_c; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178692.4]
  wire [19:0] pma_checker_OptimizationBarrier_16_io_x_ppn; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178735.4]
  wire  pma_checker_OptimizationBarrier_16_io_x_u; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178735.4]
  wire  pma_checker_OptimizationBarrier_16_io_x_ae; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178735.4]
  wire  pma_checker_OptimizationBarrier_16_io_x_sw; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178735.4]
  wire  pma_checker_OptimizationBarrier_16_io_x_sx; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178735.4]
  wire  pma_checker_OptimizationBarrier_16_io_x_sr; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178735.4]
  wire  pma_checker_OptimizationBarrier_16_io_x_pw; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178735.4]
  wire  pma_checker_OptimizationBarrier_16_io_x_px; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178735.4]
  wire  pma_checker_OptimizationBarrier_16_io_x_pr; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178735.4]
  wire  pma_checker_OptimizationBarrier_16_io_x_ppp; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178735.4]
  wire  pma_checker_OptimizationBarrier_16_io_x_pal; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178735.4]
  wire  pma_checker_OptimizationBarrier_16_io_x_paa; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178735.4]
  wire  pma_checker_OptimizationBarrier_16_io_x_eff; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178735.4]
  wire  pma_checker_OptimizationBarrier_16_io_x_c; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178735.4]
  wire [19:0] pma_checker_OptimizationBarrier_16_io_y_ppn; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178735.4]
  wire  pma_checker_OptimizationBarrier_16_io_y_u; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178735.4]
  wire  pma_checker_OptimizationBarrier_16_io_y_ae; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178735.4]
  wire  pma_checker_OptimizationBarrier_16_io_y_sw; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178735.4]
  wire  pma_checker_OptimizationBarrier_16_io_y_sx; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178735.4]
  wire  pma_checker_OptimizationBarrier_16_io_y_sr; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178735.4]
  wire  pma_checker_OptimizationBarrier_16_io_y_pw; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178735.4]
  wire  pma_checker_OptimizationBarrier_16_io_y_px; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178735.4]
  wire  pma_checker_OptimizationBarrier_16_io_y_pr; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178735.4]
  wire  pma_checker_OptimizationBarrier_16_io_y_ppp; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178735.4]
  wire  pma_checker_OptimizationBarrier_16_io_y_pal; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178735.4]
  wire  pma_checker_OptimizationBarrier_16_io_y_paa; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178735.4]
  wire  pma_checker_OptimizationBarrier_16_io_y_eff; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178735.4]
  wire  pma_checker_OptimizationBarrier_16_io_y_c; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178735.4]
  wire [19:0] pma_checker_OptimizationBarrier_17_io_x_ppn; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178778.4]
  wire  pma_checker_OptimizationBarrier_17_io_x_u; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178778.4]
  wire  pma_checker_OptimizationBarrier_17_io_x_ae; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178778.4]
  wire  pma_checker_OptimizationBarrier_17_io_x_sw; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178778.4]
  wire  pma_checker_OptimizationBarrier_17_io_x_sx; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178778.4]
  wire  pma_checker_OptimizationBarrier_17_io_x_sr; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178778.4]
  wire  pma_checker_OptimizationBarrier_17_io_x_pw; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178778.4]
  wire  pma_checker_OptimizationBarrier_17_io_x_px; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178778.4]
  wire  pma_checker_OptimizationBarrier_17_io_x_pr; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178778.4]
  wire  pma_checker_OptimizationBarrier_17_io_x_ppp; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178778.4]
  wire  pma_checker_OptimizationBarrier_17_io_x_pal; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178778.4]
  wire  pma_checker_OptimizationBarrier_17_io_x_paa; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178778.4]
  wire  pma_checker_OptimizationBarrier_17_io_x_eff; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178778.4]
  wire  pma_checker_OptimizationBarrier_17_io_x_c; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178778.4]
  wire [19:0] pma_checker_OptimizationBarrier_17_io_y_ppn; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178778.4]
  wire  pma_checker_OptimizationBarrier_17_io_y_u; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178778.4]
  wire  pma_checker_OptimizationBarrier_17_io_y_ae; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178778.4]
  wire  pma_checker_OptimizationBarrier_17_io_y_sw; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178778.4]
  wire  pma_checker_OptimizationBarrier_17_io_y_sx; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178778.4]
  wire  pma_checker_OptimizationBarrier_17_io_y_sr; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178778.4]
  wire  pma_checker_OptimizationBarrier_17_io_y_pw; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178778.4]
  wire  pma_checker_OptimizationBarrier_17_io_y_px; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178778.4]
  wire  pma_checker_OptimizationBarrier_17_io_y_pr; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178778.4]
  wire  pma_checker_OptimizationBarrier_17_io_y_ppp; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178778.4]
  wire  pma_checker_OptimizationBarrier_17_io_y_pal; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178778.4]
  wire  pma_checker_OptimizationBarrier_17_io_y_paa; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178778.4]
  wire  pma_checker_OptimizationBarrier_17_io_y_eff; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178778.4]
  wire  pma_checker_OptimizationBarrier_17_io_y_c; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178778.4]
  wire [19:0] pma_checker_OptimizationBarrier_18_io_x_ppn; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178821.4]
  wire  pma_checker_OptimizationBarrier_18_io_x_u; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178821.4]
  wire  pma_checker_OptimizationBarrier_18_io_x_ae; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178821.4]
  wire  pma_checker_OptimizationBarrier_18_io_x_sw; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178821.4]
  wire  pma_checker_OptimizationBarrier_18_io_x_sx; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178821.4]
  wire  pma_checker_OptimizationBarrier_18_io_x_sr; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178821.4]
  wire  pma_checker_OptimizationBarrier_18_io_x_pw; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178821.4]
  wire  pma_checker_OptimizationBarrier_18_io_x_px; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178821.4]
  wire  pma_checker_OptimizationBarrier_18_io_x_pr; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178821.4]
  wire  pma_checker_OptimizationBarrier_18_io_x_ppp; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178821.4]
  wire  pma_checker_OptimizationBarrier_18_io_x_pal; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178821.4]
  wire  pma_checker_OptimizationBarrier_18_io_x_paa; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178821.4]
  wire  pma_checker_OptimizationBarrier_18_io_x_eff; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178821.4]
  wire  pma_checker_OptimizationBarrier_18_io_x_c; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178821.4]
  wire [19:0] pma_checker_OptimizationBarrier_18_io_y_ppn; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178821.4]
  wire  pma_checker_OptimizationBarrier_18_io_y_u; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178821.4]
  wire  pma_checker_OptimizationBarrier_18_io_y_ae; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178821.4]
  wire  pma_checker_OptimizationBarrier_18_io_y_sw; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178821.4]
  wire  pma_checker_OptimizationBarrier_18_io_y_sx; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178821.4]
  wire  pma_checker_OptimizationBarrier_18_io_y_sr; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178821.4]
  wire  pma_checker_OptimizationBarrier_18_io_y_pw; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178821.4]
  wire  pma_checker_OptimizationBarrier_18_io_y_px; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178821.4]
  wire  pma_checker_OptimizationBarrier_18_io_y_pr; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178821.4]
  wire  pma_checker_OptimizationBarrier_18_io_y_ppp; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178821.4]
  wire  pma_checker_OptimizationBarrier_18_io_y_pal; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178821.4]
  wire  pma_checker_OptimizationBarrier_18_io_y_paa; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178821.4]
  wire  pma_checker_OptimizationBarrier_18_io_y_eff; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178821.4]
  wire  pma_checker_OptimizationBarrier_18_io_y_c; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178821.4]
  wire [19:0] pma_checker_OptimizationBarrier_19_io_x_ppn; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178864.4]
  wire  pma_checker_OptimizationBarrier_19_io_x_u; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178864.4]
  wire  pma_checker_OptimizationBarrier_19_io_x_ae; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178864.4]
  wire  pma_checker_OptimizationBarrier_19_io_x_sw; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178864.4]
  wire  pma_checker_OptimizationBarrier_19_io_x_sx; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178864.4]
  wire  pma_checker_OptimizationBarrier_19_io_x_sr; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178864.4]
  wire  pma_checker_OptimizationBarrier_19_io_x_pw; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178864.4]
  wire  pma_checker_OptimizationBarrier_19_io_x_px; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178864.4]
  wire  pma_checker_OptimizationBarrier_19_io_x_pr; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178864.4]
  wire  pma_checker_OptimizationBarrier_19_io_x_ppp; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178864.4]
  wire  pma_checker_OptimizationBarrier_19_io_x_pal; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178864.4]
  wire  pma_checker_OptimizationBarrier_19_io_x_paa; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178864.4]
  wire  pma_checker_OptimizationBarrier_19_io_x_eff; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178864.4]
  wire  pma_checker_OptimizationBarrier_19_io_x_c; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178864.4]
  wire [19:0] pma_checker_OptimizationBarrier_19_io_y_ppn; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178864.4]
  wire  pma_checker_OptimizationBarrier_19_io_y_u; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178864.4]
  wire  pma_checker_OptimizationBarrier_19_io_y_ae; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178864.4]
  wire  pma_checker_OptimizationBarrier_19_io_y_sw; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178864.4]
  wire  pma_checker_OptimizationBarrier_19_io_y_sx; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178864.4]
  wire  pma_checker_OptimizationBarrier_19_io_y_sr; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178864.4]
  wire  pma_checker_OptimizationBarrier_19_io_y_pw; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178864.4]
  wire  pma_checker_OptimizationBarrier_19_io_y_px; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178864.4]
  wire  pma_checker_OptimizationBarrier_19_io_y_pr; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178864.4]
  wire  pma_checker_OptimizationBarrier_19_io_y_ppp; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178864.4]
  wire  pma_checker_OptimizationBarrier_19_io_y_pal; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178864.4]
  wire  pma_checker_OptimizationBarrier_19_io_y_paa; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178864.4]
  wire  pma_checker_OptimizationBarrier_19_io_y_eff; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178864.4]
  wire  pma_checker_OptimizationBarrier_19_io_y_c; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178864.4]
  wire [19:0] pma_checker_OptimizationBarrier_20_io_x_ppn; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178907.4]
  wire  pma_checker_OptimizationBarrier_20_io_x_u; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178907.4]
  wire  pma_checker_OptimizationBarrier_20_io_x_ae; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178907.4]
  wire  pma_checker_OptimizationBarrier_20_io_x_sw; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178907.4]
  wire  pma_checker_OptimizationBarrier_20_io_x_sx; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178907.4]
  wire  pma_checker_OptimizationBarrier_20_io_x_sr; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178907.4]
  wire  pma_checker_OptimizationBarrier_20_io_x_pw; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178907.4]
  wire  pma_checker_OptimizationBarrier_20_io_x_px; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178907.4]
  wire  pma_checker_OptimizationBarrier_20_io_x_pr; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178907.4]
  wire  pma_checker_OptimizationBarrier_20_io_x_ppp; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178907.4]
  wire  pma_checker_OptimizationBarrier_20_io_x_pal; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178907.4]
  wire  pma_checker_OptimizationBarrier_20_io_x_paa; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178907.4]
  wire  pma_checker_OptimizationBarrier_20_io_x_eff; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178907.4]
  wire  pma_checker_OptimizationBarrier_20_io_x_c; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178907.4]
  wire [19:0] pma_checker_OptimizationBarrier_20_io_y_ppn; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178907.4]
  wire  pma_checker_OptimizationBarrier_20_io_y_u; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178907.4]
  wire  pma_checker_OptimizationBarrier_20_io_y_ae; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178907.4]
  wire  pma_checker_OptimizationBarrier_20_io_y_sw; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178907.4]
  wire  pma_checker_OptimizationBarrier_20_io_y_sx; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178907.4]
  wire  pma_checker_OptimizationBarrier_20_io_y_sr; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178907.4]
  wire  pma_checker_OptimizationBarrier_20_io_y_pw; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178907.4]
  wire  pma_checker_OptimizationBarrier_20_io_y_px; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178907.4]
  wire  pma_checker_OptimizationBarrier_20_io_y_pr; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178907.4]
  wire  pma_checker_OptimizationBarrier_20_io_y_ppp; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178907.4]
  wire  pma_checker_OptimizationBarrier_20_io_y_pal; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178907.4]
  wire  pma_checker_OptimizationBarrier_20_io_y_paa; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178907.4]
  wire  pma_checker_OptimizationBarrier_20_io_y_eff; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178907.4]
  wire  pma_checker_OptimizationBarrier_20_io_y_c; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178907.4]
  wire [19:0] pma_checker_OptimizationBarrier_21_io_x_ppn; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178950.4]
  wire  pma_checker_OptimizationBarrier_21_io_x_u; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178950.4]
  wire  pma_checker_OptimizationBarrier_21_io_x_ae; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178950.4]
  wire  pma_checker_OptimizationBarrier_21_io_x_sw; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178950.4]
  wire  pma_checker_OptimizationBarrier_21_io_x_sx; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178950.4]
  wire  pma_checker_OptimizationBarrier_21_io_x_sr; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178950.4]
  wire  pma_checker_OptimizationBarrier_21_io_x_pw; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178950.4]
  wire  pma_checker_OptimizationBarrier_21_io_x_px; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178950.4]
  wire  pma_checker_OptimizationBarrier_21_io_x_pr; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178950.4]
  wire  pma_checker_OptimizationBarrier_21_io_x_ppp; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178950.4]
  wire  pma_checker_OptimizationBarrier_21_io_x_pal; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178950.4]
  wire  pma_checker_OptimizationBarrier_21_io_x_paa; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178950.4]
  wire  pma_checker_OptimizationBarrier_21_io_x_eff; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178950.4]
  wire  pma_checker_OptimizationBarrier_21_io_x_c; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178950.4]
  wire [19:0] pma_checker_OptimizationBarrier_21_io_y_ppn; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178950.4]
  wire  pma_checker_OptimizationBarrier_21_io_y_u; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178950.4]
  wire  pma_checker_OptimizationBarrier_21_io_y_ae; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178950.4]
  wire  pma_checker_OptimizationBarrier_21_io_y_sw; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178950.4]
  wire  pma_checker_OptimizationBarrier_21_io_y_sx; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178950.4]
  wire  pma_checker_OptimizationBarrier_21_io_y_sr; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178950.4]
  wire  pma_checker_OptimizationBarrier_21_io_y_pw; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178950.4]
  wire  pma_checker_OptimizationBarrier_21_io_y_px; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178950.4]
  wire  pma_checker_OptimizationBarrier_21_io_y_pr; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178950.4]
  wire  pma_checker_OptimizationBarrier_21_io_y_ppp; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178950.4]
  wire  pma_checker_OptimizationBarrier_21_io_y_pal; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178950.4]
  wire  pma_checker_OptimizationBarrier_21_io_y_paa; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178950.4]
  wire  pma_checker_OptimizationBarrier_21_io_y_eff; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178950.4]
  wire  pma_checker_OptimizationBarrier_21_io_y_c; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178950.4]
  wire [19:0] pma_checker_OptimizationBarrier_22_io_x_ppn; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178992.4]
  wire  pma_checker_OptimizationBarrier_22_io_x_u; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178992.4]
  wire  pma_checker_OptimizationBarrier_22_io_x_ae; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178992.4]
  wire  pma_checker_OptimizationBarrier_22_io_x_sw; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178992.4]
  wire  pma_checker_OptimizationBarrier_22_io_x_sx; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178992.4]
  wire  pma_checker_OptimizationBarrier_22_io_x_sr; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178992.4]
  wire  pma_checker_OptimizationBarrier_22_io_x_pw; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178992.4]
  wire  pma_checker_OptimizationBarrier_22_io_x_px; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178992.4]
  wire  pma_checker_OptimizationBarrier_22_io_x_pr; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178992.4]
  wire  pma_checker_OptimizationBarrier_22_io_x_ppp; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178992.4]
  wire  pma_checker_OptimizationBarrier_22_io_x_pal; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178992.4]
  wire  pma_checker_OptimizationBarrier_22_io_x_paa; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178992.4]
  wire  pma_checker_OptimizationBarrier_22_io_x_eff; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178992.4]
  wire  pma_checker_OptimizationBarrier_22_io_x_c; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178992.4]
  wire [19:0] pma_checker_OptimizationBarrier_22_io_y_ppn; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178992.4]
  wire  pma_checker_OptimizationBarrier_22_io_y_u; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178992.4]
  wire  pma_checker_OptimizationBarrier_22_io_y_ae; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178992.4]
  wire  pma_checker_OptimizationBarrier_22_io_y_sw; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178992.4]
  wire  pma_checker_OptimizationBarrier_22_io_y_sx; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178992.4]
  wire  pma_checker_OptimizationBarrier_22_io_y_sr; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178992.4]
  wire  pma_checker_OptimizationBarrier_22_io_y_pw; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178992.4]
  wire  pma_checker_OptimizationBarrier_22_io_y_px; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178992.4]
  wire  pma_checker_OptimizationBarrier_22_io_y_pr; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178992.4]
  wire  pma_checker_OptimizationBarrier_22_io_y_ppp; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178992.4]
  wire  pma_checker_OptimizationBarrier_22_io_y_pal; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178992.4]
  wire  pma_checker_OptimizationBarrier_22_io_y_paa; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178992.4]
  wire  pma_checker_OptimizationBarrier_22_io_y_eff; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178992.4]
  wire  pma_checker_OptimizationBarrier_22_io_y_c; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178992.4]
  wire [19:0] pma_checker_OptimizationBarrier_23_io_x_ppn; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179034.4]
  wire  pma_checker_OptimizationBarrier_23_io_x_u; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179034.4]
  wire  pma_checker_OptimizationBarrier_23_io_x_ae; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179034.4]
  wire  pma_checker_OptimizationBarrier_23_io_x_sw; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179034.4]
  wire  pma_checker_OptimizationBarrier_23_io_x_sx; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179034.4]
  wire  pma_checker_OptimizationBarrier_23_io_x_sr; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179034.4]
  wire  pma_checker_OptimizationBarrier_23_io_x_pw; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179034.4]
  wire  pma_checker_OptimizationBarrier_23_io_x_px; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179034.4]
  wire  pma_checker_OptimizationBarrier_23_io_x_pr; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179034.4]
  wire  pma_checker_OptimizationBarrier_23_io_x_ppp; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179034.4]
  wire  pma_checker_OptimizationBarrier_23_io_x_pal; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179034.4]
  wire  pma_checker_OptimizationBarrier_23_io_x_paa; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179034.4]
  wire  pma_checker_OptimizationBarrier_23_io_x_eff; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179034.4]
  wire  pma_checker_OptimizationBarrier_23_io_x_c; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179034.4]
  wire [19:0] pma_checker_OptimizationBarrier_23_io_y_ppn; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179034.4]
  wire  pma_checker_OptimizationBarrier_23_io_y_u; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179034.4]
  wire  pma_checker_OptimizationBarrier_23_io_y_ae; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179034.4]
  wire  pma_checker_OptimizationBarrier_23_io_y_sw; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179034.4]
  wire  pma_checker_OptimizationBarrier_23_io_y_sx; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179034.4]
  wire  pma_checker_OptimizationBarrier_23_io_y_sr; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179034.4]
  wire  pma_checker_OptimizationBarrier_23_io_y_pw; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179034.4]
  wire  pma_checker_OptimizationBarrier_23_io_y_px; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179034.4]
  wire  pma_checker_OptimizationBarrier_23_io_y_pr; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179034.4]
  wire  pma_checker_OptimizationBarrier_23_io_y_ppp; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179034.4]
  wire  pma_checker_OptimizationBarrier_23_io_y_pal; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179034.4]
  wire  pma_checker_OptimizationBarrier_23_io_y_paa; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179034.4]
  wire  pma_checker_OptimizationBarrier_23_io_y_eff; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179034.4]
  wire  pma_checker_OptimizationBarrier_23_io_y_c; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179034.4]
  wire [19:0] pma_checker_OptimizationBarrier_24_io_x_ppn; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179076.4]
  wire  pma_checker_OptimizationBarrier_24_io_x_u; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179076.4]
  wire  pma_checker_OptimizationBarrier_24_io_x_ae; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179076.4]
  wire  pma_checker_OptimizationBarrier_24_io_x_sw; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179076.4]
  wire  pma_checker_OptimizationBarrier_24_io_x_sx; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179076.4]
  wire  pma_checker_OptimizationBarrier_24_io_x_sr; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179076.4]
  wire  pma_checker_OptimizationBarrier_24_io_x_pw; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179076.4]
  wire  pma_checker_OptimizationBarrier_24_io_x_px; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179076.4]
  wire  pma_checker_OptimizationBarrier_24_io_x_pr; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179076.4]
  wire  pma_checker_OptimizationBarrier_24_io_x_ppp; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179076.4]
  wire  pma_checker_OptimizationBarrier_24_io_x_pal; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179076.4]
  wire  pma_checker_OptimizationBarrier_24_io_x_paa; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179076.4]
  wire  pma_checker_OptimizationBarrier_24_io_x_eff; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179076.4]
  wire  pma_checker_OptimizationBarrier_24_io_x_c; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179076.4]
  wire [19:0] pma_checker_OptimizationBarrier_24_io_y_ppn; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179076.4]
  wire  pma_checker_OptimizationBarrier_24_io_y_u; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179076.4]
  wire  pma_checker_OptimizationBarrier_24_io_y_ae; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179076.4]
  wire  pma_checker_OptimizationBarrier_24_io_y_sw; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179076.4]
  wire  pma_checker_OptimizationBarrier_24_io_y_sx; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179076.4]
  wire  pma_checker_OptimizationBarrier_24_io_y_sr; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179076.4]
  wire  pma_checker_OptimizationBarrier_24_io_y_pw; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179076.4]
  wire  pma_checker_OptimizationBarrier_24_io_y_px; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179076.4]
  wire  pma_checker_OptimizationBarrier_24_io_y_pr; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179076.4]
  wire  pma_checker_OptimizationBarrier_24_io_y_ppp; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179076.4]
  wire  pma_checker_OptimizationBarrier_24_io_y_pal; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179076.4]
  wire  pma_checker_OptimizationBarrier_24_io_y_paa; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179076.4]
  wire  pma_checker_OptimizationBarrier_24_io_y_eff; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179076.4]
  wire  pma_checker_OptimizationBarrier_24_io_y_c; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179076.4]
  wire [19:0] pma_checker_OptimizationBarrier_25_io_x_ppn; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179118.4]
  wire  pma_checker_OptimizationBarrier_25_io_x_u; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179118.4]
  wire  pma_checker_OptimizationBarrier_25_io_x_ae; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179118.4]
  wire  pma_checker_OptimizationBarrier_25_io_x_sw; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179118.4]
  wire  pma_checker_OptimizationBarrier_25_io_x_sx; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179118.4]
  wire  pma_checker_OptimizationBarrier_25_io_x_sr; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179118.4]
  wire  pma_checker_OptimizationBarrier_25_io_x_pw; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179118.4]
  wire  pma_checker_OptimizationBarrier_25_io_x_px; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179118.4]
  wire  pma_checker_OptimizationBarrier_25_io_x_pr; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179118.4]
  wire  pma_checker_OptimizationBarrier_25_io_x_ppp; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179118.4]
  wire  pma_checker_OptimizationBarrier_25_io_x_pal; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179118.4]
  wire  pma_checker_OptimizationBarrier_25_io_x_paa; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179118.4]
  wire  pma_checker_OptimizationBarrier_25_io_x_eff; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179118.4]
  wire  pma_checker_OptimizationBarrier_25_io_x_c; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179118.4]
  wire [19:0] pma_checker_OptimizationBarrier_25_io_y_ppn; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179118.4]
  wire  pma_checker_OptimizationBarrier_25_io_y_u; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179118.4]
  wire  pma_checker_OptimizationBarrier_25_io_y_ae; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179118.4]
  wire  pma_checker_OptimizationBarrier_25_io_y_sw; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179118.4]
  wire  pma_checker_OptimizationBarrier_25_io_y_sx; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179118.4]
  wire  pma_checker_OptimizationBarrier_25_io_y_sr; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179118.4]
  wire  pma_checker_OptimizationBarrier_25_io_y_pw; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179118.4]
  wire  pma_checker_OptimizationBarrier_25_io_y_px; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179118.4]
  wire  pma_checker_OptimizationBarrier_25_io_y_pr; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179118.4]
  wire  pma_checker_OptimizationBarrier_25_io_y_ppp; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179118.4]
  wire  pma_checker_OptimizationBarrier_25_io_y_pal; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179118.4]
  wire  pma_checker_OptimizationBarrier_25_io_y_paa; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179118.4]
  wire  pma_checker_OptimizationBarrier_25_io_y_eff; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179118.4]
  wire  pma_checker_OptimizationBarrier_25_io_y_c; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179118.4]
  wire [19:0] pma_checker_OptimizationBarrier_26_io_x_ppn; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179160.4]
  wire  pma_checker_OptimizationBarrier_26_io_x_u; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179160.4]
  wire  pma_checker_OptimizationBarrier_26_io_x_ae; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179160.4]
  wire  pma_checker_OptimizationBarrier_26_io_x_sw; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179160.4]
  wire  pma_checker_OptimizationBarrier_26_io_x_sx; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179160.4]
  wire  pma_checker_OptimizationBarrier_26_io_x_sr; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179160.4]
  wire  pma_checker_OptimizationBarrier_26_io_x_pw; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179160.4]
  wire  pma_checker_OptimizationBarrier_26_io_x_px; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179160.4]
  wire  pma_checker_OptimizationBarrier_26_io_x_pr; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179160.4]
  wire  pma_checker_OptimizationBarrier_26_io_x_ppp; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179160.4]
  wire  pma_checker_OptimizationBarrier_26_io_x_pal; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179160.4]
  wire  pma_checker_OptimizationBarrier_26_io_x_paa; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179160.4]
  wire  pma_checker_OptimizationBarrier_26_io_x_eff; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179160.4]
  wire  pma_checker_OptimizationBarrier_26_io_x_c; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179160.4]
  wire [19:0] pma_checker_OptimizationBarrier_26_io_y_ppn; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179160.4]
  wire  pma_checker_OptimizationBarrier_26_io_y_u; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179160.4]
  wire  pma_checker_OptimizationBarrier_26_io_y_ae; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179160.4]
  wire  pma_checker_OptimizationBarrier_26_io_y_sw; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179160.4]
  wire  pma_checker_OptimizationBarrier_26_io_y_sx; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179160.4]
  wire  pma_checker_OptimizationBarrier_26_io_y_sr; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179160.4]
  wire  pma_checker_OptimizationBarrier_26_io_y_pw; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179160.4]
  wire  pma_checker_OptimizationBarrier_26_io_y_px; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179160.4]
  wire  pma_checker_OptimizationBarrier_26_io_y_pr; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179160.4]
  wire  pma_checker_OptimizationBarrier_26_io_y_ppp; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179160.4]
  wire  pma_checker_OptimizationBarrier_26_io_y_pal; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179160.4]
  wire  pma_checker_OptimizationBarrier_26_io_y_paa; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179160.4]
  wire  pma_checker_OptimizationBarrier_26_io_y_eff; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179160.4]
  wire  pma_checker_OptimizationBarrier_26_io_y_c; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179160.4]
  wire [19:0] pma_checker_OptimizationBarrier_27_io_x_ppn; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179203.4]
  wire  pma_checker_OptimizationBarrier_27_io_x_u; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179203.4]
  wire  pma_checker_OptimizationBarrier_27_io_x_ae; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179203.4]
  wire  pma_checker_OptimizationBarrier_27_io_x_sw; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179203.4]
  wire  pma_checker_OptimizationBarrier_27_io_x_sx; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179203.4]
  wire  pma_checker_OptimizationBarrier_27_io_x_sr; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179203.4]
  wire  pma_checker_OptimizationBarrier_27_io_x_pw; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179203.4]
  wire  pma_checker_OptimizationBarrier_27_io_x_px; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179203.4]
  wire  pma_checker_OptimizationBarrier_27_io_x_pr; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179203.4]
  wire  pma_checker_OptimizationBarrier_27_io_x_ppp; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179203.4]
  wire  pma_checker_OptimizationBarrier_27_io_x_pal; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179203.4]
  wire  pma_checker_OptimizationBarrier_27_io_x_paa; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179203.4]
  wire  pma_checker_OptimizationBarrier_27_io_x_eff; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179203.4]
  wire  pma_checker_OptimizationBarrier_27_io_x_c; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179203.4]
  wire [19:0] pma_checker_OptimizationBarrier_27_io_y_ppn; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179203.4]
  wire  pma_checker_OptimizationBarrier_27_io_y_u; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179203.4]
  wire  pma_checker_OptimizationBarrier_27_io_y_ae; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179203.4]
  wire  pma_checker_OptimizationBarrier_27_io_y_sw; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179203.4]
  wire  pma_checker_OptimizationBarrier_27_io_y_sx; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179203.4]
  wire  pma_checker_OptimizationBarrier_27_io_y_sr; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179203.4]
  wire  pma_checker_OptimizationBarrier_27_io_y_pw; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179203.4]
  wire  pma_checker_OptimizationBarrier_27_io_y_px; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179203.4]
  wire  pma_checker_OptimizationBarrier_27_io_y_pr; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179203.4]
  wire  pma_checker_OptimizationBarrier_27_io_y_ppp; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179203.4]
  wire  pma_checker_OptimizationBarrier_27_io_y_pal; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179203.4]
  wire  pma_checker_OptimizationBarrier_27_io_y_paa; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179203.4]
  wire  pma_checker_OptimizationBarrier_27_io_y_eff; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179203.4]
  wire  pma_checker_OptimizationBarrier_27_io_y_c; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179203.4]
  wire [19:0] pma_checker_OptimizationBarrier_28_io_x_ppn; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179246.4]
  wire  pma_checker_OptimizationBarrier_28_io_x_u; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179246.4]
  wire  pma_checker_OptimizationBarrier_28_io_x_ae; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179246.4]
  wire  pma_checker_OptimizationBarrier_28_io_x_sw; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179246.4]
  wire  pma_checker_OptimizationBarrier_28_io_x_sx; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179246.4]
  wire  pma_checker_OptimizationBarrier_28_io_x_sr; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179246.4]
  wire  pma_checker_OptimizationBarrier_28_io_x_pw; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179246.4]
  wire  pma_checker_OptimizationBarrier_28_io_x_px; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179246.4]
  wire  pma_checker_OptimizationBarrier_28_io_x_pr; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179246.4]
  wire  pma_checker_OptimizationBarrier_28_io_x_ppp; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179246.4]
  wire  pma_checker_OptimizationBarrier_28_io_x_pal; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179246.4]
  wire  pma_checker_OptimizationBarrier_28_io_x_paa; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179246.4]
  wire  pma_checker_OptimizationBarrier_28_io_x_eff; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179246.4]
  wire  pma_checker_OptimizationBarrier_28_io_x_c; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179246.4]
  wire [19:0] pma_checker_OptimizationBarrier_28_io_y_ppn; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179246.4]
  wire  pma_checker_OptimizationBarrier_28_io_y_u; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179246.4]
  wire  pma_checker_OptimizationBarrier_28_io_y_ae; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179246.4]
  wire  pma_checker_OptimizationBarrier_28_io_y_sw; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179246.4]
  wire  pma_checker_OptimizationBarrier_28_io_y_sx; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179246.4]
  wire  pma_checker_OptimizationBarrier_28_io_y_sr; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179246.4]
  wire  pma_checker_OptimizationBarrier_28_io_y_pw; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179246.4]
  wire  pma_checker_OptimizationBarrier_28_io_y_px; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179246.4]
  wire  pma_checker_OptimizationBarrier_28_io_y_pr; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179246.4]
  wire  pma_checker_OptimizationBarrier_28_io_y_ppp; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179246.4]
  wire  pma_checker_OptimizationBarrier_28_io_y_pal; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179246.4]
  wire  pma_checker_OptimizationBarrier_28_io_y_paa; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179246.4]
  wire  pma_checker_OptimizationBarrier_28_io_y_eff; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179246.4]
  wire  pma_checker_OptimizationBarrier_28_io_y_c; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179246.4]
  wire [19:0] pma_checker_OptimizationBarrier_29_io_x_ppn; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179289.4]
  wire  pma_checker_OptimizationBarrier_29_io_x_u; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179289.4]
  wire  pma_checker_OptimizationBarrier_29_io_x_ae; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179289.4]
  wire  pma_checker_OptimizationBarrier_29_io_x_sw; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179289.4]
  wire  pma_checker_OptimizationBarrier_29_io_x_sx; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179289.4]
  wire  pma_checker_OptimizationBarrier_29_io_x_sr; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179289.4]
  wire  pma_checker_OptimizationBarrier_29_io_x_pw; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179289.4]
  wire  pma_checker_OptimizationBarrier_29_io_x_px; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179289.4]
  wire  pma_checker_OptimizationBarrier_29_io_x_pr; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179289.4]
  wire  pma_checker_OptimizationBarrier_29_io_x_ppp; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179289.4]
  wire  pma_checker_OptimizationBarrier_29_io_x_pal; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179289.4]
  wire  pma_checker_OptimizationBarrier_29_io_x_paa; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179289.4]
  wire  pma_checker_OptimizationBarrier_29_io_x_eff; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179289.4]
  wire  pma_checker_OptimizationBarrier_29_io_x_c; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179289.4]
  wire [19:0] pma_checker_OptimizationBarrier_29_io_y_ppn; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179289.4]
  wire  pma_checker_OptimizationBarrier_29_io_y_u; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179289.4]
  wire  pma_checker_OptimizationBarrier_29_io_y_ae; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179289.4]
  wire  pma_checker_OptimizationBarrier_29_io_y_sw; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179289.4]
  wire  pma_checker_OptimizationBarrier_29_io_y_sx; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179289.4]
  wire  pma_checker_OptimizationBarrier_29_io_y_sr; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179289.4]
  wire  pma_checker_OptimizationBarrier_29_io_y_pw; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179289.4]
  wire  pma_checker_OptimizationBarrier_29_io_y_px; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179289.4]
  wire  pma_checker_OptimizationBarrier_29_io_y_pr; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179289.4]
  wire  pma_checker_OptimizationBarrier_29_io_y_ppp; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179289.4]
  wire  pma_checker_OptimizationBarrier_29_io_y_pal; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179289.4]
  wire  pma_checker_OptimizationBarrier_29_io_y_paa; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179289.4]
  wire  pma_checker_OptimizationBarrier_29_io_y_eff; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179289.4]
  wire  pma_checker_OptimizationBarrier_29_io_y_c; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179289.4]
  wire [19:0] pma_checker_OptimizationBarrier_30_io_x_ppn; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179332.4]
  wire  pma_checker_OptimizationBarrier_30_io_x_u; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179332.4]
  wire  pma_checker_OptimizationBarrier_30_io_x_ae; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179332.4]
  wire  pma_checker_OptimizationBarrier_30_io_x_sw; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179332.4]
  wire  pma_checker_OptimizationBarrier_30_io_x_sx; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179332.4]
  wire  pma_checker_OptimizationBarrier_30_io_x_sr; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179332.4]
  wire  pma_checker_OptimizationBarrier_30_io_x_pw; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179332.4]
  wire  pma_checker_OptimizationBarrier_30_io_x_px; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179332.4]
  wire  pma_checker_OptimizationBarrier_30_io_x_pr; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179332.4]
  wire  pma_checker_OptimizationBarrier_30_io_x_ppp; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179332.4]
  wire  pma_checker_OptimizationBarrier_30_io_x_pal; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179332.4]
  wire  pma_checker_OptimizationBarrier_30_io_x_paa; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179332.4]
  wire  pma_checker_OptimizationBarrier_30_io_x_eff; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179332.4]
  wire  pma_checker_OptimizationBarrier_30_io_x_c; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179332.4]
  wire [19:0] pma_checker_OptimizationBarrier_30_io_y_ppn; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179332.4]
  wire  pma_checker_OptimizationBarrier_30_io_y_u; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179332.4]
  wire  pma_checker_OptimizationBarrier_30_io_y_ae; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179332.4]
  wire  pma_checker_OptimizationBarrier_30_io_y_sw; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179332.4]
  wire  pma_checker_OptimizationBarrier_30_io_y_sx; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179332.4]
  wire  pma_checker_OptimizationBarrier_30_io_y_sr; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179332.4]
  wire  pma_checker_OptimizationBarrier_30_io_y_pw; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179332.4]
  wire  pma_checker_OptimizationBarrier_30_io_y_px; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179332.4]
  wire  pma_checker_OptimizationBarrier_30_io_y_pr; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179332.4]
  wire  pma_checker_OptimizationBarrier_30_io_y_ppp; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179332.4]
  wire  pma_checker_OptimizationBarrier_30_io_y_pal; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179332.4]
  wire  pma_checker_OptimizationBarrier_30_io_y_paa; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179332.4]
  wire  pma_checker_OptimizationBarrier_30_io_y_eff; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179332.4]
  wire  pma_checker_OptimizationBarrier_30_io_y_c; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179332.4]
  wire [19:0] pma_checker_OptimizationBarrier_31_io_x_ppn; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179375.4]
  wire  pma_checker_OptimizationBarrier_31_io_x_u; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179375.4]
  wire  pma_checker_OptimizationBarrier_31_io_x_ae; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179375.4]
  wire  pma_checker_OptimizationBarrier_31_io_x_sw; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179375.4]
  wire  pma_checker_OptimizationBarrier_31_io_x_sx; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179375.4]
  wire  pma_checker_OptimizationBarrier_31_io_x_sr; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179375.4]
  wire  pma_checker_OptimizationBarrier_31_io_x_pw; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179375.4]
  wire  pma_checker_OptimizationBarrier_31_io_x_px; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179375.4]
  wire  pma_checker_OptimizationBarrier_31_io_x_pr; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179375.4]
  wire  pma_checker_OptimizationBarrier_31_io_x_ppp; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179375.4]
  wire  pma_checker_OptimizationBarrier_31_io_x_pal; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179375.4]
  wire  pma_checker_OptimizationBarrier_31_io_x_paa; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179375.4]
  wire  pma_checker_OptimizationBarrier_31_io_x_eff; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179375.4]
  wire  pma_checker_OptimizationBarrier_31_io_x_c; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179375.4]
  wire [19:0] pma_checker_OptimizationBarrier_31_io_y_ppn; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179375.4]
  wire  pma_checker_OptimizationBarrier_31_io_y_u; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179375.4]
  wire  pma_checker_OptimizationBarrier_31_io_y_ae; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179375.4]
  wire  pma_checker_OptimizationBarrier_31_io_y_sw; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179375.4]
  wire  pma_checker_OptimizationBarrier_31_io_y_sx; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179375.4]
  wire  pma_checker_OptimizationBarrier_31_io_y_sr; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179375.4]
  wire  pma_checker_OptimizationBarrier_31_io_y_pw; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179375.4]
  wire  pma_checker_OptimizationBarrier_31_io_y_px; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179375.4]
  wire  pma_checker_OptimizationBarrier_31_io_y_pr; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179375.4]
  wire  pma_checker_OptimizationBarrier_31_io_y_ppp; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179375.4]
  wire  pma_checker_OptimizationBarrier_31_io_y_pal; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179375.4]
  wire  pma_checker_OptimizationBarrier_31_io_y_paa; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179375.4]
  wire  pma_checker_OptimizationBarrier_31_io_y_eff; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179375.4]
  wire  pma_checker_OptimizationBarrier_31_io_y_c; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179375.4]
  wire [19:0] pma_checker_OptimizationBarrier_32_io_x_ppn; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179418.4]
  wire  pma_checker_OptimizationBarrier_32_io_x_u; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179418.4]
  wire  pma_checker_OptimizationBarrier_32_io_x_ae; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179418.4]
  wire  pma_checker_OptimizationBarrier_32_io_x_sw; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179418.4]
  wire  pma_checker_OptimizationBarrier_32_io_x_sx; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179418.4]
  wire  pma_checker_OptimizationBarrier_32_io_x_sr; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179418.4]
  wire  pma_checker_OptimizationBarrier_32_io_x_pw; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179418.4]
  wire  pma_checker_OptimizationBarrier_32_io_x_px; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179418.4]
  wire  pma_checker_OptimizationBarrier_32_io_x_pr; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179418.4]
  wire  pma_checker_OptimizationBarrier_32_io_x_ppp; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179418.4]
  wire  pma_checker_OptimizationBarrier_32_io_x_pal; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179418.4]
  wire  pma_checker_OptimizationBarrier_32_io_x_paa; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179418.4]
  wire  pma_checker_OptimizationBarrier_32_io_x_eff; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179418.4]
  wire  pma_checker_OptimizationBarrier_32_io_x_c; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179418.4]
  wire [19:0] pma_checker_OptimizationBarrier_32_io_y_ppn; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179418.4]
  wire  pma_checker_OptimizationBarrier_32_io_y_u; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179418.4]
  wire  pma_checker_OptimizationBarrier_32_io_y_ae; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179418.4]
  wire  pma_checker_OptimizationBarrier_32_io_y_sw; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179418.4]
  wire  pma_checker_OptimizationBarrier_32_io_y_sx; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179418.4]
  wire  pma_checker_OptimizationBarrier_32_io_y_sr; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179418.4]
  wire  pma_checker_OptimizationBarrier_32_io_y_pw; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179418.4]
  wire  pma_checker_OptimizationBarrier_32_io_y_px; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179418.4]
  wire  pma_checker_OptimizationBarrier_32_io_y_pr; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179418.4]
  wire  pma_checker_OptimizationBarrier_32_io_y_ppp; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179418.4]
  wire  pma_checker_OptimizationBarrier_32_io_y_pal; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179418.4]
  wire  pma_checker_OptimizationBarrier_32_io_y_paa; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179418.4]
  wire  pma_checker_OptimizationBarrier_32_io_y_eff; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179418.4]
  wire  pma_checker_OptimizationBarrier_32_io_y_c; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179418.4]
  wire [19:0] pma_checker_OptimizationBarrier_33_io_x_ppn; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179461.4]
  wire  pma_checker_OptimizationBarrier_33_io_x_u; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179461.4]
  wire  pma_checker_OptimizationBarrier_33_io_x_ae; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179461.4]
  wire  pma_checker_OptimizationBarrier_33_io_x_sw; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179461.4]
  wire  pma_checker_OptimizationBarrier_33_io_x_sx; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179461.4]
  wire  pma_checker_OptimizationBarrier_33_io_x_sr; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179461.4]
  wire  pma_checker_OptimizationBarrier_33_io_x_pw; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179461.4]
  wire  pma_checker_OptimizationBarrier_33_io_x_px; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179461.4]
  wire  pma_checker_OptimizationBarrier_33_io_x_pr; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179461.4]
  wire  pma_checker_OptimizationBarrier_33_io_x_ppp; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179461.4]
  wire  pma_checker_OptimizationBarrier_33_io_x_pal; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179461.4]
  wire  pma_checker_OptimizationBarrier_33_io_x_paa; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179461.4]
  wire  pma_checker_OptimizationBarrier_33_io_x_eff; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179461.4]
  wire  pma_checker_OptimizationBarrier_33_io_x_c; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179461.4]
  wire [19:0] pma_checker_OptimizationBarrier_33_io_y_ppn; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179461.4]
  wire  pma_checker_OptimizationBarrier_33_io_y_u; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179461.4]
  wire  pma_checker_OptimizationBarrier_33_io_y_ae; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179461.4]
  wire  pma_checker_OptimizationBarrier_33_io_y_sw; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179461.4]
  wire  pma_checker_OptimizationBarrier_33_io_y_sx; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179461.4]
  wire  pma_checker_OptimizationBarrier_33_io_y_sr; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179461.4]
  wire  pma_checker_OptimizationBarrier_33_io_y_pw; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179461.4]
  wire  pma_checker_OptimizationBarrier_33_io_y_px; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179461.4]
  wire  pma_checker_OptimizationBarrier_33_io_y_pr; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179461.4]
  wire  pma_checker_OptimizationBarrier_33_io_y_ppp; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179461.4]
  wire  pma_checker_OptimizationBarrier_33_io_y_pal; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179461.4]
  wire  pma_checker_OptimizationBarrier_33_io_y_paa; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179461.4]
  wire  pma_checker_OptimizationBarrier_33_io_y_eff; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179461.4]
  wire  pma_checker_OptimizationBarrier_33_io_y_c; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179461.4]
  wire [19:0] pma_checker_OptimizationBarrier_34_io_x_ppn; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179504.4]
  wire  pma_checker_OptimizationBarrier_34_io_x_u; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179504.4]
  wire  pma_checker_OptimizationBarrier_34_io_x_ae; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179504.4]
  wire  pma_checker_OptimizationBarrier_34_io_x_sw; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179504.4]
  wire  pma_checker_OptimizationBarrier_34_io_x_sx; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179504.4]
  wire  pma_checker_OptimizationBarrier_34_io_x_sr; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179504.4]
  wire  pma_checker_OptimizationBarrier_34_io_x_pw; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179504.4]
  wire  pma_checker_OptimizationBarrier_34_io_x_px; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179504.4]
  wire  pma_checker_OptimizationBarrier_34_io_x_pr; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179504.4]
  wire  pma_checker_OptimizationBarrier_34_io_x_ppp; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179504.4]
  wire  pma_checker_OptimizationBarrier_34_io_x_pal; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179504.4]
  wire  pma_checker_OptimizationBarrier_34_io_x_paa; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179504.4]
  wire  pma_checker_OptimizationBarrier_34_io_x_eff; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179504.4]
  wire  pma_checker_OptimizationBarrier_34_io_x_c; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179504.4]
  wire [19:0] pma_checker_OptimizationBarrier_34_io_y_ppn; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179504.4]
  wire  pma_checker_OptimizationBarrier_34_io_y_u; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179504.4]
  wire  pma_checker_OptimizationBarrier_34_io_y_ae; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179504.4]
  wire  pma_checker_OptimizationBarrier_34_io_y_sw; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179504.4]
  wire  pma_checker_OptimizationBarrier_34_io_y_sx; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179504.4]
  wire  pma_checker_OptimizationBarrier_34_io_y_sr; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179504.4]
  wire  pma_checker_OptimizationBarrier_34_io_y_pw; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179504.4]
  wire  pma_checker_OptimizationBarrier_34_io_y_px; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179504.4]
  wire  pma_checker_OptimizationBarrier_34_io_y_pr; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179504.4]
  wire  pma_checker_OptimizationBarrier_34_io_y_ppp; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179504.4]
  wire  pma_checker_OptimizationBarrier_34_io_y_pal; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179504.4]
  wire  pma_checker_OptimizationBarrier_34_io_y_paa; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179504.4]
  wire  pma_checker_OptimizationBarrier_34_io_y_eff; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179504.4]
  wire  pma_checker_OptimizationBarrier_34_io_y_c; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179504.4]
  wire [19:0] pma_checker_OptimizationBarrier_35_io_x_ppn; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179546.4]
  wire  pma_checker_OptimizationBarrier_35_io_x_u; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179546.4]
  wire  pma_checker_OptimizationBarrier_35_io_x_ae; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179546.4]
  wire  pma_checker_OptimizationBarrier_35_io_x_sw; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179546.4]
  wire  pma_checker_OptimizationBarrier_35_io_x_sx; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179546.4]
  wire  pma_checker_OptimizationBarrier_35_io_x_sr; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179546.4]
  wire  pma_checker_OptimizationBarrier_35_io_x_pw; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179546.4]
  wire  pma_checker_OptimizationBarrier_35_io_x_px; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179546.4]
  wire  pma_checker_OptimizationBarrier_35_io_x_pr; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179546.4]
  wire  pma_checker_OptimizationBarrier_35_io_x_ppp; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179546.4]
  wire  pma_checker_OptimizationBarrier_35_io_x_pal; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179546.4]
  wire  pma_checker_OptimizationBarrier_35_io_x_paa; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179546.4]
  wire  pma_checker_OptimizationBarrier_35_io_x_eff; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179546.4]
  wire  pma_checker_OptimizationBarrier_35_io_x_c; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179546.4]
  wire [19:0] pma_checker_OptimizationBarrier_35_io_y_ppn; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179546.4]
  wire  pma_checker_OptimizationBarrier_35_io_y_u; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179546.4]
  wire  pma_checker_OptimizationBarrier_35_io_y_ae; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179546.4]
  wire  pma_checker_OptimizationBarrier_35_io_y_sw; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179546.4]
  wire  pma_checker_OptimizationBarrier_35_io_y_sx; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179546.4]
  wire  pma_checker_OptimizationBarrier_35_io_y_sr; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179546.4]
  wire  pma_checker_OptimizationBarrier_35_io_y_pw; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179546.4]
  wire  pma_checker_OptimizationBarrier_35_io_y_px; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179546.4]
  wire  pma_checker_OptimizationBarrier_35_io_y_pr; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179546.4]
  wire  pma_checker_OptimizationBarrier_35_io_y_ppp; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179546.4]
  wire  pma_checker_OptimizationBarrier_35_io_y_pal; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179546.4]
  wire  pma_checker_OptimizationBarrier_35_io_y_paa; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179546.4]
  wire  pma_checker_OptimizationBarrier_35_io_y_eff; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179546.4]
  wire  pma_checker_OptimizationBarrier_35_io_y_c; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179546.4]
  wire [19:0] pma_checker_OptimizationBarrier_36_io_x_ppn; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179588.4]
  wire  pma_checker_OptimizationBarrier_36_io_x_u; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179588.4]
  wire  pma_checker_OptimizationBarrier_36_io_x_ae; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179588.4]
  wire  pma_checker_OptimizationBarrier_36_io_x_sw; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179588.4]
  wire  pma_checker_OptimizationBarrier_36_io_x_sx; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179588.4]
  wire  pma_checker_OptimizationBarrier_36_io_x_sr; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179588.4]
  wire  pma_checker_OptimizationBarrier_36_io_x_pw; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179588.4]
  wire  pma_checker_OptimizationBarrier_36_io_x_px; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179588.4]
  wire  pma_checker_OptimizationBarrier_36_io_x_pr; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179588.4]
  wire  pma_checker_OptimizationBarrier_36_io_x_ppp; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179588.4]
  wire  pma_checker_OptimizationBarrier_36_io_x_pal; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179588.4]
  wire  pma_checker_OptimizationBarrier_36_io_x_paa; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179588.4]
  wire  pma_checker_OptimizationBarrier_36_io_x_eff; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179588.4]
  wire  pma_checker_OptimizationBarrier_36_io_x_c; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179588.4]
  wire [19:0] pma_checker_OptimizationBarrier_36_io_y_ppn; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179588.4]
  wire  pma_checker_OptimizationBarrier_36_io_y_u; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179588.4]
  wire  pma_checker_OptimizationBarrier_36_io_y_ae; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179588.4]
  wire  pma_checker_OptimizationBarrier_36_io_y_sw; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179588.4]
  wire  pma_checker_OptimizationBarrier_36_io_y_sx; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179588.4]
  wire  pma_checker_OptimizationBarrier_36_io_y_sr; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179588.4]
  wire  pma_checker_OptimizationBarrier_36_io_y_pw; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179588.4]
  wire  pma_checker_OptimizationBarrier_36_io_y_px; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179588.4]
  wire  pma_checker_OptimizationBarrier_36_io_y_pr; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179588.4]
  wire  pma_checker_OptimizationBarrier_36_io_y_ppp; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179588.4]
  wire  pma_checker_OptimizationBarrier_36_io_y_pal; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179588.4]
  wire  pma_checker_OptimizationBarrier_36_io_y_paa; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179588.4]
  wire  pma_checker_OptimizationBarrier_36_io_y_eff; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179588.4]
  wire  pma_checker_OptimizationBarrier_36_io_y_c; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179588.4]
  wire [19:0] pma_checker_OptimizationBarrier_37_io_x_ppn; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179630.4]
  wire  pma_checker_OptimizationBarrier_37_io_x_u; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179630.4]
  wire  pma_checker_OptimizationBarrier_37_io_x_ae; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179630.4]
  wire  pma_checker_OptimizationBarrier_37_io_x_sw; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179630.4]
  wire  pma_checker_OptimizationBarrier_37_io_x_sx; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179630.4]
  wire  pma_checker_OptimizationBarrier_37_io_x_sr; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179630.4]
  wire  pma_checker_OptimizationBarrier_37_io_x_pw; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179630.4]
  wire  pma_checker_OptimizationBarrier_37_io_x_px; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179630.4]
  wire  pma_checker_OptimizationBarrier_37_io_x_pr; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179630.4]
  wire  pma_checker_OptimizationBarrier_37_io_x_ppp; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179630.4]
  wire  pma_checker_OptimizationBarrier_37_io_x_pal; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179630.4]
  wire  pma_checker_OptimizationBarrier_37_io_x_paa; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179630.4]
  wire  pma_checker_OptimizationBarrier_37_io_x_eff; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179630.4]
  wire  pma_checker_OptimizationBarrier_37_io_x_c; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179630.4]
  wire [19:0] pma_checker_OptimizationBarrier_37_io_y_ppn; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179630.4]
  wire  pma_checker_OptimizationBarrier_37_io_y_u; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179630.4]
  wire  pma_checker_OptimizationBarrier_37_io_y_ae; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179630.4]
  wire  pma_checker_OptimizationBarrier_37_io_y_sw; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179630.4]
  wire  pma_checker_OptimizationBarrier_37_io_y_sx; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179630.4]
  wire  pma_checker_OptimizationBarrier_37_io_y_sr; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179630.4]
  wire  pma_checker_OptimizationBarrier_37_io_y_pw; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179630.4]
  wire  pma_checker_OptimizationBarrier_37_io_y_px; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179630.4]
  wire  pma_checker_OptimizationBarrier_37_io_y_pr; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179630.4]
  wire  pma_checker_OptimizationBarrier_37_io_y_ppp; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179630.4]
  wire  pma_checker_OptimizationBarrier_37_io_y_pal; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179630.4]
  wire  pma_checker_OptimizationBarrier_37_io_y_paa; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179630.4]
  wire  pma_checker_OptimizationBarrier_37_io_y_eff; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179630.4]
  wire  pma_checker_OptimizationBarrier_37_io_y_c; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179630.4]
  wire [19:0] pma_checker_OptimizationBarrier_38_io_x_ppn; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179672.4]
  wire  pma_checker_OptimizationBarrier_38_io_x_u; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179672.4]
  wire  pma_checker_OptimizationBarrier_38_io_x_ae; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179672.4]
  wire  pma_checker_OptimizationBarrier_38_io_x_sw; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179672.4]
  wire  pma_checker_OptimizationBarrier_38_io_x_sx; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179672.4]
  wire  pma_checker_OptimizationBarrier_38_io_x_sr; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179672.4]
  wire  pma_checker_OptimizationBarrier_38_io_x_pw; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179672.4]
  wire  pma_checker_OptimizationBarrier_38_io_x_px; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179672.4]
  wire  pma_checker_OptimizationBarrier_38_io_x_pr; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179672.4]
  wire  pma_checker_OptimizationBarrier_38_io_x_ppp; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179672.4]
  wire  pma_checker_OptimizationBarrier_38_io_x_pal; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179672.4]
  wire  pma_checker_OptimizationBarrier_38_io_x_paa; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179672.4]
  wire  pma_checker_OptimizationBarrier_38_io_x_eff; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179672.4]
  wire  pma_checker_OptimizationBarrier_38_io_x_c; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179672.4]
  wire [19:0] pma_checker_OptimizationBarrier_38_io_y_ppn; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179672.4]
  wire  pma_checker_OptimizationBarrier_38_io_y_u; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179672.4]
  wire  pma_checker_OptimizationBarrier_38_io_y_ae; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179672.4]
  wire  pma_checker_OptimizationBarrier_38_io_y_sw; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179672.4]
  wire  pma_checker_OptimizationBarrier_38_io_y_sx; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179672.4]
  wire  pma_checker_OptimizationBarrier_38_io_y_sr; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179672.4]
  wire  pma_checker_OptimizationBarrier_38_io_y_pw; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179672.4]
  wire  pma_checker_OptimizationBarrier_38_io_y_px; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179672.4]
  wire  pma_checker_OptimizationBarrier_38_io_y_pr; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179672.4]
  wire  pma_checker_OptimizationBarrier_38_io_y_ppp; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179672.4]
  wire  pma_checker_OptimizationBarrier_38_io_y_pal; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179672.4]
  wire  pma_checker_OptimizationBarrier_38_io_y_paa; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179672.4]
  wire  pma_checker_OptimizationBarrier_38_io_y_eff; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179672.4]
  wire  pma_checker_OptimizationBarrier_38_io_y_c; // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179672.4]
  wire  pma_checker__T_2026; // @[OneHot.scala 32:14:freechips.rocketchip.system.DefaultRV32Config.fir@180088.8]
  wire  MaxPeriodFibonacciLFSR_clock; // @[PRNG.scala 82:22:freechips.rocketchip.system.DefaultRV32Config.fir@192119.4]
  wire  MaxPeriodFibonacciLFSR_reset; // @[PRNG.scala 82:22:freechips.rocketchip.system.DefaultRV32Config.fir@192119.4]
  wire  MaxPeriodFibonacciLFSR_io_increment; // @[PRNG.scala 82:22:freechips.rocketchip.system.DefaultRV32Config.fir@192119.4]
  wire  MaxPeriodFibonacciLFSR_io_out_0; // @[PRNG.scala 82:22:freechips.rocketchip.system.DefaultRV32Config.fir@192119.4]
  wire  MaxPeriodFibonacciLFSR_io_out_1; // @[PRNG.scala 82:22:freechips.rocketchip.system.DefaultRV32Config.fir@192119.4]
  wire  MaxPeriodFibonacciLFSR_io_out_2; // @[PRNG.scala 82:22:freechips.rocketchip.system.DefaultRV32Config.fir@192119.4]
  wire  MaxPeriodFibonacciLFSR_io_out_3; // @[PRNG.scala 82:22:freechips.rocketchip.system.DefaultRV32Config.fir@192119.4]
  wire  MaxPeriodFibonacciLFSR_io_out_4; // @[PRNG.scala 82:22:freechips.rocketchip.system.DefaultRV32Config.fir@192119.4]
  wire  MaxPeriodFibonacciLFSR_io_out_5; // @[PRNG.scala 82:22:freechips.rocketchip.system.DefaultRV32Config.fir@192119.4]
  wire  MaxPeriodFibonacciLFSR_io_out_6; // @[PRNG.scala 82:22:freechips.rocketchip.system.DefaultRV32Config.fir@192119.4]
  wire  MaxPeriodFibonacciLFSR_io_out_7; // @[PRNG.scala 82:22:freechips.rocketchip.system.DefaultRV32Config.fir@192119.4]
  wire  MaxPeriodFibonacciLFSR_io_out_8; // @[PRNG.scala 82:22:freechips.rocketchip.system.DefaultRV32Config.fir@192119.4]
  wire  MaxPeriodFibonacciLFSR_io_out_9; // @[PRNG.scala 82:22:freechips.rocketchip.system.DefaultRV32Config.fir@192119.4]
  wire  MaxPeriodFibonacciLFSR_io_out_10; // @[PRNG.scala 82:22:freechips.rocketchip.system.DefaultRV32Config.fir@192119.4]
  wire  MaxPeriodFibonacciLFSR_io_out_11; // @[PRNG.scala 82:22:freechips.rocketchip.system.DefaultRV32Config.fir@192119.4]
  wire  MaxPeriodFibonacciLFSR_io_out_12; // @[PRNG.scala 82:22:freechips.rocketchip.system.DefaultRV32Config.fir@192119.4]
  wire  MaxPeriodFibonacciLFSR_io_out_13; // @[PRNG.scala 82:22:freechips.rocketchip.system.DefaultRV32Config.fir@192119.4]
  wire  MaxPeriodFibonacciLFSR_io_out_14; // @[PRNG.scala 82:22:freechips.rocketchip.system.DefaultRV32Config.fir@192119.4]
  wire  MaxPeriodFibonacciLFSR_io_out_15; // @[PRNG.scala 82:22:freechips.rocketchip.system.DefaultRV32Config.fir@192119.4]
  wire  metaArb_io_in_0_valid; // @[:freechips.rocketchip.system.DefaultRV32Config.fir@191714.4]
  wire [31:0] metaArb_io_in_0_bits_addr; // @[:freechips.rocketchip.system.DefaultRV32Config.fir@191714.4]
  wire [5:0] metaArb_io_in_0_bits_idx; // @[:freechips.rocketchip.system.DefaultRV32Config.fir@191714.4]
  wire [21:0] metaArb_io_in_0_bits_data; // @[:freechips.rocketchip.system.DefaultRV32Config.fir@191714.4]
  wire  metaArb_io_in_1_valid; // @[:freechips.rocketchip.system.DefaultRV32Config.fir@191714.4]
  wire [31:0] metaArb_io_in_1_bits_addr; // @[:freechips.rocketchip.system.DefaultRV32Config.fir@191714.4]
  wire [5:0] metaArb_io_in_1_bits_idx; // @[:freechips.rocketchip.system.DefaultRV32Config.fir@191714.4]
  wire [21:0] metaArb_io_in_1_bits_data; // @[:freechips.rocketchip.system.DefaultRV32Config.fir@191714.4]
  wire  metaArb_io_in_2_valid; // @[:freechips.rocketchip.system.DefaultRV32Config.fir@191714.4]
  wire [31:0] metaArb_io_in_2_bits_addr; // @[:freechips.rocketchip.system.DefaultRV32Config.fir@191714.4]
  wire [5:0] metaArb_io_in_2_bits_idx; // @[:freechips.rocketchip.system.DefaultRV32Config.fir@191714.4]
  wire [3:0] metaArb_io_in_2_bits_way_en; // @[:freechips.rocketchip.system.DefaultRV32Config.fir@191714.4]
  wire [21:0] metaArb_io_in_2_bits_data; // @[:freechips.rocketchip.system.DefaultRV32Config.fir@191714.4]
  wire  metaArb_io_in_3_valid; // @[:freechips.rocketchip.system.DefaultRV32Config.fir@191714.4]
  wire [31:0] metaArb_io_in_3_bits_addr; // @[:freechips.rocketchip.system.DefaultRV32Config.fir@191714.4]
  wire [5:0] metaArb_io_in_3_bits_idx; // @[:freechips.rocketchip.system.DefaultRV32Config.fir@191714.4]
  wire [3:0] metaArb_io_in_3_bits_way_en; // @[:freechips.rocketchip.system.DefaultRV32Config.fir@191714.4]
  wire [21:0] metaArb_io_in_3_bits_data; // @[:freechips.rocketchip.system.DefaultRV32Config.fir@191714.4]
  wire  metaArb_io_in_4_ready; // @[:freechips.rocketchip.system.DefaultRV32Config.fir@191714.4]
  wire  metaArb_io_in_4_valid; // @[:freechips.rocketchip.system.DefaultRV32Config.fir@191714.4]
  wire [31:0] metaArb_io_in_4_bits_addr; // @[:freechips.rocketchip.system.DefaultRV32Config.fir@191714.4]
  wire [5:0] metaArb_io_in_4_bits_idx; // @[:freechips.rocketchip.system.DefaultRV32Config.fir@191714.4]
  wire [3:0] metaArb_io_in_4_bits_way_en; // @[:freechips.rocketchip.system.DefaultRV32Config.fir@191714.4]
  wire [21:0] metaArb_io_in_4_bits_data; // @[:freechips.rocketchip.system.DefaultRV32Config.fir@191714.4]
  wire [31:0] metaArb_io_in_5_bits_addr; // @[:freechips.rocketchip.system.DefaultRV32Config.fir@191714.4]
  wire [5:0] metaArb_io_in_5_bits_idx; // @[:freechips.rocketchip.system.DefaultRV32Config.fir@191714.4]
  wire  metaArb_io_in_6_ready; // @[:freechips.rocketchip.system.DefaultRV32Config.fir@191714.4]
  wire  metaArb_io_in_6_valid; // @[:freechips.rocketchip.system.DefaultRV32Config.fir@191714.4]
  wire [31:0] metaArb_io_in_6_bits_addr; // @[:freechips.rocketchip.system.DefaultRV32Config.fir@191714.4]
  wire [5:0] metaArb_io_in_6_bits_idx; // @[:freechips.rocketchip.system.DefaultRV32Config.fir@191714.4]
  wire [3:0] metaArb_io_in_6_bits_way_en; // @[:freechips.rocketchip.system.DefaultRV32Config.fir@191714.4]
  wire [21:0] metaArb_io_in_6_bits_data; // @[:freechips.rocketchip.system.DefaultRV32Config.fir@191714.4]
  wire  metaArb_io_in_7_ready; // @[:freechips.rocketchip.system.DefaultRV32Config.fir@191714.4]
  wire  metaArb_io_in_7_valid; // @[:freechips.rocketchip.system.DefaultRV32Config.fir@191714.4]
  wire [31:0] metaArb_io_in_7_bits_addr; // @[:freechips.rocketchip.system.DefaultRV32Config.fir@191714.4]
  wire [5:0] metaArb_io_in_7_bits_idx; // @[:freechips.rocketchip.system.DefaultRV32Config.fir@191714.4]
  wire [3:0] metaArb_io_in_7_bits_way_en; // @[:freechips.rocketchip.system.DefaultRV32Config.fir@191714.4]
  wire [21:0] metaArb_io_in_7_bits_data; // @[:freechips.rocketchip.system.DefaultRV32Config.fir@191714.4]
  wire  metaArb_io_out_valid; // @[:freechips.rocketchip.system.DefaultRV32Config.fir@191714.4]
  wire  metaArb_io_out_bits_write; // @[:freechips.rocketchip.system.DefaultRV32Config.fir@191714.4]
  wire [31:0] metaArb_io_out_bits_addr; // @[:freechips.rocketchip.system.DefaultRV32Config.fir@191714.4]
  wire [5:0] metaArb_io_out_bits_idx; // @[:freechips.rocketchip.system.DefaultRV32Config.fir@191714.4]
  wire [3:0] metaArb_io_out_bits_way_en; // @[:freechips.rocketchip.system.DefaultRV32Config.fir@191714.4]
  wire [21:0] metaArb_io_out_bits_data; // @[:freechips.rocketchip.system.DefaultRV32Config.fir@191714.4]
  wire [21:0] metaArb__GEN_1; // @[Arbiter.scala 126:27:freechips.rocketchip.system.DefaultRV32Config.fir@191722.4]
  wire [3:0] metaArb__GEN_2; // @[Arbiter.scala 126:27:freechips.rocketchip.system.DefaultRV32Config.fir@191722.4]
  wire [5:0] metaArb__GEN_3; // @[Arbiter.scala 126:27:freechips.rocketchip.system.DefaultRV32Config.fir@191722.4]
  wire [31:0] metaArb__GEN_4; // @[Arbiter.scala 126:27:freechips.rocketchip.system.DefaultRV32Config.fir@191722.4]
  wire [21:0] metaArb__GEN_13; // @[Arbiter.scala 126:27:freechips.rocketchip.system.DefaultRV32Config.fir@191738.4]
  wire [3:0] metaArb__GEN_14; // @[Arbiter.scala 126:27:freechips.rocketchip.system.DefaultRV32Config.fir@191738.4]
  wire [5:0] metaArb__GEN_15; // @[Arbiter.scala 126:27:freechips.rocketchip.system.DefaultRV32Config.fir@191738.4]
  wire [31:0] metaArb__GEN_16; // @[Arbiter.scala 126:27:freechips.rocketchip.system.DefaultRV32Config.fir@191738.4]
  wire [21:0] metaArb__GEN_19; // @[Arbiter.scala 126:27:freechips.rocketchip.system.DefaultRV32Config.fir@191746.4]
  wire [3:0] metaArb__GEN_20; // @[Arbiter.scala 126:27:freechips.rocketchip.system.DefaultRV32Config.fir@191746.4]
  wire [5:0] metaArb__GEN_21; // @[Arbiter.scala 126:27:freechips.rocketchip.system.DefaultRV32Config.fir@191746.4]
  wire [31:0] metaArb__GEN_22; // @[Arbiter.scala 126:27:freechips.rocketchip.system.DefaultRV32Config.fir@191746.4]
  wire  metaArb__GEN_23; // @[Arbiter.scala 126:27:freechips.rocketchip.system.DefaultRV32Config.fir@191746.4]
  wire [21:0] metaArb__GEN_25; // @[Arbiter.scala 126:27:freechips.rocketchip.system.DefaultRV32Config.fir@191754.4]
  wire [3:0] metaArb__GEN_26; // @[Arbiter.scala 126:27:freechips.rocketchip.system.DefaultRV32Config.fir@191754.4]
  wire [5:0] metaArb__GEN_27; // @[Arbiter.scala 126:27:freechips.rocketchip.system.DefaultRV32Config.fir@191754.4]
  wire [31:0] metaArb__GEN_28; // @[Arbiter.scala 126:27:freechips.rocketchip.system.DefaultRV32Config.fir@191754.4]
  wire  metaArb__GEN_29; // @[Arbiter.scala 126:27:freechips.rocketchip.system.DefaultRV32Config.fir@191754.4]
  wire [21:0] metaArb__GEN_31; // @[Arbiter.scala 126:27:freechips.rocketchip.system.DefaultRV32Config.fir@191762.4]
  wire [3:0] metaArb__GEN_32; // @[Arbiter.scala 126:27:freechips.rocketchip.system.DefaultRV32Config.fir@191762.4]
  wire [5:0] metaArb__GEN_33; // @[Arbiter.scala 126:27:freechips.rocketchip.system.DefaultRV32Config.fir@191762.4]
  wire [31:0] metaArb__GEN_34; // @[Arbiter.scala 126:27:freechips.rocketchip.system.DefaultRV32Config.fir@191762.4]
  wire  metaArb__GEN_35; // @[Arbiter.scala 126:27:freechips.rocketchip.system.DefaultRV32Config.fir@191762.4]
  wire  metaArb__T; // @[Arbiter.scala 31:68:freechips.rocketchip.system.DefaultRV32Config.fir@191778.4]
  wire  metaArb__T_1; // @[Arbiter.scala 31:68:freechips.rocketchip.system.DefaultRV32Config.fir@191779.4]
  wire  metaArb__T_2; // @[Arbiter.scala 31:68:freechips.rocketchip.system.DefaultRV32Config.fir@191780.4]
  wire  metaArb__T_3; // @[Arbiter.scala 31:68:freechips.rocketchip.system.DefaultRV32Config.fir@191781.4]
  wire  metaArb__T_5; // @[Arbiter.scala 31:68:freechips.rocketchip.system.DefaultRV32Config.fir@191783.4]
  wire  metaArb_grant_7; // @[Arbiter.scala 31:78:freechips.rocketchip.system.DefaultRV32Config.fir@191790.4]
  wire  metaArb__T_14; // @[Arbiter.scala 135:19:freechips.rocketchip.system.DefaultRV32Config.fir@191807.4]
  wire [5:0] tag_array_RW0_addr; // @[DescribedSRAM.scala 23:26:freechips.rocketchip.system.DefaultRV32Config.fir@192159.4]
  wire  tag_array_RW0_en; // @[DescribedSRAM.scala 23:26:freechips.rocketchip.system.DefaultRV32Config.fir@192159.4]
  wire  tag_array_RW0_clk; // @[DescribedSRAM.scala 23:26:freechips.rocketchip.system.DefaultRV32Config.fir@192159.4]
  wire  tag_array_RW0_wmode; // @[DescribedSRAM.scala 23:26:freechips.rocketchip.system.DefaultRV32Config.fir@192159.4]
  wire [21:0] tag_array_RW0_wdata_0; // @[DescribedSRAM.scala 23:26:freechips.rocketchip.system.DefaultRV32Config.fir@192159.4]
  wire [21:0] tag_array_RW0_wdata_1; // @[DescribedSRAM.scala 23:26:freechips.rocketchip.system.DefaultRV32Config.fir@192159.4]
  wire [21:0] tag_array_RW0_wdata_2; // @[DescribedSRAM.scala 23:26:freechips.rocketchip.system.DefaultRV32Config.fir@192159.4]
  wire [21:0] tag_array_RW0_wdata_3; // @[DescribedSRAM.scala 23:26:freechips.rocketchip.system.DefaultRV32Config.fir@192159.4]
  wire [21:0] tag_array_RW0_rdata_0; // @[DescribedSRAM.scala 23:26:freechips.rocketchip.system.DefaultRV32Config.fir@192159.4]
  wire [21:0] tag_array_RW0_rdata_1; // @[DescribedSRAM.scala 23:26:freechips.rocketchip.system.DefaultRV32Config.fir@192159.4]
  wire [21:0] tag_array_RW0_rdata_2; // @[DescribedSRAM.scala 23:26:freechips.rocketchip.system.DefaultRV32Config.fir@192159.4]
  wire [21:0] tag_array_RW0_rdata_3; // @[DescribedSRAM.scala 23:26:freechips.rocketchip.system.DefaultRV32Config.fir@192159.4]
  wire  tag_array_RW0_wmask_0; // @[DescribedSRAM.scala 23:26:freechips.rocketchip.system.DefaultRV32Config.fir@192159.4]
  wire  tag_array_RW0_wmask_1; // @[DescribedSRAM.scala 23:26:freechips.rocketchip.system.DefaultRV32Config.fir@192159.4]
  wire  tag_array_RW0_wmask_2; // @[DescribedSRAM.scala 23:26:freechips.rocketchip.system.DefaultRV32Config.fir@192159.4]
  wire  tag_array_RW0_wmask_3; // @[DescribedSRAM.scala 23:26:freechips.rocketchip.system.DefaultRV32Config.fir@192159.4]
  wire  data_clock; // @[DCache.scala 130:20:freechips.rocketchip.system.DefaultRV32Config.fir@192160.4]
  wire  data_io_req_valid; // @[DCache.scala 130:20:freechips.rocketchip.system.DefaultRV32Config.fir@192160.4]
  wire [11:0] data_io_req_bits_addr; // @[DCache.scala 130:20:freechips.rocketchip.system.DefaultRV32Config.fir@192160.4]
  wire  data_io_req_bits_write; // @[DCache.scala 130:20:freechips.rocketchip.system.DefaultRV32Config.fir@192160.4]
  wire [31:0] data_io_req_bits_wdata; // @[DCache.scala 130:20:freechips.rocketchip.system.DefaultRV32Config.fir@192160.4]
  wire [3:0] data_io_req_bits_eccMask; // @[DCache.scala 130:20:freechips.rocketchip.system.DefaultRV32Config.fir@192160.4]
  wire [3:0] data_io_req_bits_way_en; // @[DCache.scala 130:20:freechips.rocketchip.system.DefaultRV32Config.fir@192160.4]
  wire [31:0] data_io_resp_0; // @[DCache.scala 130:20:freechips.rocketchip.system.DefaultRV32Config.fir@192160.4]
  wire [31:0] data_io_resp_1; // @[DCache.scala 130:20:freechips.rocketchip.system.DefaultRV32Config.fir@192160.4]
  wire [31:0] data_io_resp_2; // @[DCache.scala 130:20:freechips.rocketchip.system.DefaultRV32Config.fir@192160.4]
  wire [31:0] data_io_resp_3; // @[DCache.scala 130:20:freechips.rocketchip.system.DefaultRV32Config.fir@192160.4]
  wire  dataArb_io_in_0_valid; // @[:freechips.rocketchip.system.DefaultRV32Config.fir@191966.4]
  wire [11:0] dataArb_io_in_0_bits_addr; // @[:freechips.rocketchip.system.DefaultRV32Config.fir@191966.4]
  wire  dataArb_io_in_0_bits_write; // @[:freechips.rocketchip.system.DefaultRV32Config.fir@191966.4]
  wire [31:0] dataArb_io_in_0_bits_wdata; // @[:freechips.rocketchip.system.DefaultRV32Config.fir@191966.4]
  wire [3:0] dataArb_io_in_0_bits_eccMask; // @[:freechips.rocketchip.system.DefaultRV32Config.fir@191966.4]
  wire [3:0] dataArb_io_in_0_bits_way_en; // @[:freechips.rocketchip.system.DefaultRV32Config.fir@191966.4]
  wire  dataArb_io_in_1_ready; // @[:freechips.rocketchip.system.DefaultRV32Config.fir@191966.4]
  wire  dataArb_io_in_1_valid; // @[:freechips.rocketchip.system.DefaultRV32Config.fir@191966.4]
  wire [11:0] dataArb_io_in_1_bits_addr; // @[:freechips.rocketchip.system.DefaultRV32Config.fir@191966.4]
  wire  dataArb_io_in_1_bits_write; // @[:freechips.rocketchip.system.DefaultRV32Config.fir@191966.4]
  wire [31:0] dataArb_io_in_1_bits_wdata; // @[:freechips.rocketchip.system.DefaultRV32Config.fir@191966.4]
  wire [3:0] dataArb_io_in_1_bits_way_en; // @[:freechips.rocketchip.system.DefaultRV32Config.fir@191966.4]
  wire  dataArb_io_in_2_ready; // @[:freechips.rocketchip.system.DefaultRV32Config.fir@191966.4]
  wire  dataArb_io_in_2_valid; // @[:freechips.rocketchip.system.DefaultRV32Config.fir@191966.4]
  wire [11:0] dataArb_io_in_2_bits_addr; // @[:freechips.rocketchip.system.DefaultRV32Config.fir@191966.4]
  wire [31:0] dataArb_io_in_2_bits_wdata; // @[:freechips.rocketchip.system.DefaultRV32Config.fir@191966.4]
  wire  dataArb_io_in_3_ready; // @[:freechips.rocketchip.system.DefaultRV32Config.fir@191966.4]
  wire  dataArb_io_in_3_valid; // @[:freechips.rocketchip.system.DefaultRV32Config.fir@191966.4]
  wire [11:0] dataArb_io_in_3_bits_addr; // @[:freechips.rocketchip.system.DefaultRV32Config.fir@191966.4]
  wire [31:0] dataArb_io_in_3_bits_wdata; // @[:freechips.rocketchip.system.DefaultRV32Config.fir@191966.4]
  wire  dataArb_io_out_valid; // @[:freechips.rocketchip.system.DefaultRV32Config.fir@191966.4]
  wire [11:0] dataArb_io_out_bits_addr; // @[:freechips.rocketchip.system.DefaultRV32Config.fir@191966.4]
  wire  dataArb_io_out_bits_write; // @[:freechips.rocketchip.system.DefaultRV32Config.fir@191966.4]
  wire [31:0] dataArb_io_out_bits_wdata; // @[:freechips.rocketchip.system.DefaultRV32Config.fir@191966.4]
  wire [3:0] dataArb_io_out_bits_eccMask; // @[:freechips.rocketchip.system.DefaultRV32Config.fir@191966.4]
  wire [3:0] dataArb_io_out_bits_way_en; // @[:freechips.rocketchip.system.DefaultRV32Config.fir@191966.4]
  wire [31:0] dataArb__GEN_4; // @[Arbiter.scala 126:27:freechips.rocketchip.system.DefaultRV32Config.fir@191975.4]
  wire [11:0] dataArb__GEN_6; // @[Arbiter.scala 126:27:freechips.rocketchip.system.DefaultRV32Config.fir@191975.4]
  wire [3:0] dataArb__GEN_8; // @[Arbiter.scala 126:27:freechips.rocketchip.system.DefaultRV32Config.fir@191984.4]
  wire [31:0] dataArb__GEN_11; // @[Arbiter.scala 126:27:freechips.rocketchip.system.DefaultRV32Config.fir@191984.4]
  wire  dataArb__GEN_12; // @[Arbiter.scala 126:27:freechips.rocketchip.system.DefaultRV32Config.fir@191984.4]
  wire [11:0] dataArb__GEN_13; // @[Arbiter.scala 126:27:freechips.rocketchip.system.DefaultRV32Config.fir@191984.4]
  wire  dataArb__T; // @[Arbiter.scala 31:68:freechips.rocketchip.system.DefaultRV32Config.fir@192002.4]
  wire  dataArb__T_1; // @[Arbiter.scala 31:68:freechips.rocketchip.system.DefaultRV32Config.fir@192003.4]
  wire  dataArb_grant_3; // @[Arbiter.scala 31:78:freechips.rocketchip.system.DefaultRV32Config.fir@192006.4]
  wire  dataArb__T_6; // @[Arbiter.scala 135:19:freechips.rocketchip.system.DefaultRV32Config.fir@192015.4]
  wire [3:0] amoalu_io_mask; // @[DCache.scala 881:26:freechips.rocketchip.system.DefaultRV32Config.fir@195706.4]
  wire [4:0] amoalu_io_cmd; // @[DCache.scala 881:26:freechips.rocketchip.system.DefaultRV32Config.fir@195706.4]
  wire [31:0] amoalu_io_lhs; // @[DCache.scala 881:26:freechips.rocketchip.system.DefaultRV32Config.fir@195706.4]
  wire [31:0] amoalu_io_rhs; // @[DCache.scala 881:26:freechips.rocketchip.system.DefaultRV32Config.fir@195706.4]
  wire [31:0] amoalu_io_out; // @[DCache.scala 881:26:freechips.rocketchip.system.DefaultRV32Config.fir@195706.4]
  wire [7:0] _T_7; // @[PRNG.scala 86:17:freechips.rocketchip.system.DefaultRV32Config.fir@192146.4]
  wire [15:0] _T_15; // @[PRNG.scala 86:17:freechips.rocketchip.system.DefaultRV32Config.fir@192154.4]
  wire  _T_16; // @[Decoupled.scala 40:37:freechips.rocketchip.system.DefaultRV32Config.fir@192188.4]
  reg  s1_valid; // @[DCache.scala 159:21:freechips.rocketchip.system.DefaultRV32Config.fir@192189.4]
  reg [2:0] blockProbeAfterGrantCount; // @[DCache.scala 611:38:freechips.rocketchip.system.DefaultRV32Config.fir@195083.4]
  wire  _T_2338; // @[DCache.scala 709:65:freechips.rocketchip.system.DefaultRV32Config.fir@195310.4]
  reg [6:0] lrscCount; // @[DCache.scala 423:22:freechips.rocketchip.system.DefaultRV32Config.fir@193432.4]
  wire  lrscValid; // @[DCache.scala 424:29:freechips.rocketchip.system.DefaultRV32Config.fir@193433.4]
  wire  block_probe_for_core_progress; // @[DCache.scala 709:69:freechips.rocketchip.system.DefaultRV32Config.fir@195311.4]
  reg  s1_probe; // @[DCache.scala 160:21:freechips.rocketchip.system.DefaultRV32Config.fir@192192.4]
  reg  s2_probe; // @[DCache.scala 285:21:freechips.rocketchip.system.DefaultRV32Config.fir@192766.4]
  wire  _T_365; // @[DCache.scala 286:34:freechips.rocketchip.system.DefaultRV32Config.fir@192768.4]
  reg [2:0] release_state; // @[DCache.scala 199:26:freechips.rocketchip.system.DefaultRV32Config.fir@192324.4]
  wire  _T_366; // @[DCache.scala 286:63:freechips.rocketchip.system.DefaultRV32Config.fir@192769.4]
  wire  releaseInFlight; // @[DCache.scala 286:46:freechips.rocketchip.system.DefaultRV32Config.fir@192770.4]
  reg  release_ack_wait; // @[DCache.scala 197:29:freechips.rocketchip.system.DefaultRV32Config.fir@192322.4]
  reg [31:0] release_ack_addr; // @[DCache.scala 198:29:freechips.rocketchip.system.DefaultRV32Config.fir@192323.4]
  wire [31:0] _T_2339; // @[DCache.scala 710:88:freechips.rocketchip.system.DefaultRV32Config.fir@195312.4]
  wire  _T_2341; // @[DCache.scala 710:124:freechips.rocketchip.system.DefaultRV32Config.fir@195314.4]
  wire  block_probe_for_pending_release_ack; // @[DCache.scala 710:62:freechips.rocketchip.system.DefaultRV32Config.fir@195315.4]
  wire  _T_2342; // @[DCache.scala 711:50:freechips.rocketchip.system.DefaultRV32Config.fir@195316.4]
  reg  grantInProgress; // @[DCache.scala 610:28:freechips.rocketchip.system.DefaultRV32Config.fir@195082.4]
  wire  block_probe_for_ordering; // @[DCache.scala 711:89:freechips.rocketchip.system.DefaultRV32Config.fir@195317.4]
  wire  _T_2346; // @[DCache.scala 713:79:freechips.rocketchip.system.DefaultRV32Config.fir@195322.4]
  wire  _T_2347; // @[DCache.scala 713:107:freechips.rocketchip.system.DefaultRV32Config.fir@195323.4]
  reg  s2_valid; // @[DCache.scala 283:21:freechips.rocketchip.system.DefaultRV32Config.fir@192756.4]
  wire  _T_2348; // @[DCache.scala 713:119:freechips.rocketchip.system.DefaultRV32Config.fir@195324.4]
  wire  _T_2349; // @[DCache.scala 713:47:freechips.rocketchip.system.DefaultRV32Config.fir@195325.4]
  wire  tl_out__b_ready; // @[DCache.scala 713:44:freechips.rocketchip.system.DefaultRV32Config.fir@195326.4]
  wire  _T_17; // @[Decoupled.scala 40:37:freechips.rocketchip.system.DefaultRV32Config.fir@192191.4]
  reg [1:0] probe_bits_param; // @[Reg.scala 15:16:freechips.rocketchip.system.DefaultRV32Config.fir@192195.4]
  reg [3:0] probe_bits_size; // @[Reg.scala 15:16:freechips.rocketchip.system.DefaultRV32Config.fir@192195.4]
  reg  probe_bits_source; // @[Reg.scala 15:16:freechips.rocketchip.system.DefaultRV32Config.fir@192195.4]
  reg [31:0] probe_bits_address; // @[Reg.scala 15:16:freechips.rocketchip.system.DefaultRV32Config.fir@192195.4]
  wire  _T_19; // @[DCache.scala 163:37:freechips.rocketchip.system.DefaultRV32Config.fir@192209.4]
  wire  s1_valid_masked; // @[DCache.scala 163:34:freechips.rocketchip.system.DefaultRV32Config.fir@192210.4]
  reg [1:0] s2_probe_state_state; // @[Reg.scala 15:16:freechips.rocketchip.system.DefaultRV32Config.fir@192989.4]
  wire [3:0] _T_640; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@193206.4]
  wire  _T_697; // @[Misc.scala 55:20:freechips.rocketchip.system.DefaultRV32Config.fir@193263.4]
  wire  _T_693; // @[Misc.scala 55:20:freechips.rocketchip.system.DefaultRV32Config.fir@193259.4]
  wire  _T_689; // @[Misc.scala 55:20:freechips.rocketchip.system.DefaultRV32Config.fir@193255.4]
  wire  _T_685; // @[Misc.scala 55:20:freechips.rocketchip.system.DefaultRV32Config.fir@193251.4]
  wire  _T_681; // @[Misc.scala 55:20:freechips.rocketchip.system.DefaultRV32Config.fir@193247.4]
  wire  _T_677; // @[Misc.scala 55:20:freechips.rocketchip.system.DefaultRV32Config.fir@193243.4]
  wire  _T_673; // @[Misc.scala 55:20:freechips.rocketchip.system.DefaultRV32Config.fir@193239.4]
  wire  _T_669; // @[Misc.scala 55:20:freechips.rocketchip.system.DefaultRV32Config.fir@193235.4]
  wire  _T_665; // @[Misc.scala 55:20:freechips.rocketchip.system.DefaultRV32Config.fir@193231.4]
  wire  _T_661; // @[Misc.scala 55:20:freechips.rocketchip.system.DefaultRV32Config.fir@193227.4]
  wire  _T_657; // @[Misc.scala 55:20:freechips.rocketchip.system.DefaultRV32Config.fir@193223.4]
  wire  _T_653; // @[Misc.scala 55:20:freechips.rocketchip.system.DefaultRV32Config.fir@193219.4]
  wire  _T_670; // @[Misc.scala 37:9:freechips.rocketchip.system.DefaultRV32Config.fir@193236.4]
  wire  _T_674; // @[Misc.scala 37:9:freechips.rocketchip.system.DefaultRV32Config.fir@193240.4]
  wire  _T_678; // @[Misc.scala 37:9:freechips.rocketchip.system.DefaultRV32Config.fir@193244.4]
  wire  _T_682; // @[Misc.scala 37:9:freechips.rocketchip.system.DefaultRV32Config.fir@193248.4]
  wire  _T_686; // @[Misc.scala 37:9:freechips.rocketchip.system.DefaultRV32Config.fir@193252.4]
  wire  _T_690; // @[Misc.scala 37:9:freechips.rocketchip.system.DefaultRV32Config.fir@193256.4]
  wire  _T_694; // @[Misc.scala 37:9:freechips.rocketchip.system.DefaultRV32Config.fir@193260.4]
  wire  s2_prb_ack_data; // @[Misc.scala 37:9:freechips.rocketchip.system.DefaultRV32Config.fir@193264.4]
  wire  _T_2399; // @[Metadata.scala 50:45:freechips.rocketchip.system.DefaultRV32Config.fir@195454.10]
  reg [9:0] _T_2362; // @[Edges.scala 230:27:freechips.rocketchip.system.DefaultRV32Config.fir@195344.4]
  wire  _T_2365; // @[Edges.scala 233:25:freechips.rocketchip.system.DefaultRV32Config.fir@195348.4]
  wire  _T_2410; // @[package.scala 15:47:freechips.rocketchip.system.DefaultRV32Config.fir@195507.4]
  wire  _T_2411; // @[package.scala 15:47:freechips.rocketchip.system.DefaultRV32Config.fir@195508.4]
  wire  _T_2412; // @[package.scala 64:59:freechips.rocketchip.system.DefaultRV32Config.fir@195509.4]
  wire  _T_2409; // @[DCache.scala 779:25:freechips.rocketchip.system.DefaultRV32Config.fir@195500.4]
  wire  _T_2408; // @[DCache.scala 774:25:freechips.rocketchip.system.DefaultRV32Config.fir@195492.4]
  wire [2:0] _GEN_310; // @[DCache.scala 779:48:freechips.rocketchip.system.DefaultRV32Config.fir@195501.4]
  wire [2:0] tl_out__c_bits_opcode; // @[DCache.scala 783:81:freechips.rocketchip.system.DefaultRV32Config.fir@195510.4]
  wire [3:0] tl_out__c_bits_size; // @[DCache.scala 783:81:freechips.rocketchip.system.DefaultRV32Config.fir@195510.4]
  wire [26:0] _T_2356; // @[package.scala 207:77:freechips.rocketchip.system.DefaultRV32Config.fir@195338.4]
  wire [11:0] _T_2358; // @[package.scala 207:46:freechips.rocketchip.system.DefaultRV32Config.fir@195340.4]
  wire [9:0] _T_2361; // @[Edges.scala 222:14:freechips.rocketchip.system.DefaultRV32Config.fir@195343.4]
  wire  _T_2366; // @[Edges.scala 233:47:freechips.rocketchip.system.DefaultRV32Config.fir@195349.4]
  wire  c_last; // @[Edges.scala 233:37:freechips.rocketchip.system.DefaultRV32Config.fir@195350.4]
  wire  _T_2407; // @[DCache.scala 770:25:freechips.rocketchip.system.DefaultRV32Config.fir@195485.4]
  reg  s2_release_data_valid; // @[DCache.scala 724:34:freechips.rocketchip.system.DefaultRV32Config.fir@195365.4]
  wire  c_first; // @[Edges.scala 232:25:freechips.rocketchip.system.DefaultRV32Config.fir@195347.4]
  wire  _T_2381; // @[DCache.scala 732:56:freechips.rocketchip.system.DefaultRV32Config.fir@195405.4]
  wire  _T_2382; // @[DCache.scala 732:46:freechips.rocketchip.system.DefaultRV32Config.fir@195406.4]
  wire  _T_2383; // @[DCache.scala 732:43:freechips.rocketchip.system.DefaultRV32Config.fir@195407.4]
  wire  _GEN_259; // @[DCache.scala 748:36:freechips.rocketchip.system.DefaultRV32Config.fir@195450.8]
  wire  _GEN_269; // @[DCache.scala 746:28:freechips.rocketchip.system.DefaultRV32Config.fir@195446.6]
  wire  _GEN_280; // @[DCache.scala 744:21:freechips.rocketchip.system.DefaultRV32Config.fir@195442.4]
  wire  _GEN_297; // @[DCache.scala 770:47:freechips.rocketchip.system.DefaultRV32Config.fir@195486.4]
  wire  tl_out__c_valid; // @[DCache.scala 774:48:freechips.rocketchip.system.DefaultRV32Config.fir@195493.4]
  wire  _T_2354; // @[Decoupled.scala 40:37:freechips.rocketchip.system.DefaultRV32Config.fir@195336.4]
  wire  releaseDone; // @[Edges.scala 234:22:freechips.rocketchip.system.DefaultRV32Config.fir@195351.4]
  wire  _T_2401; // @[DCache.scala 756:22:freechips.rocketchip.system.DefaultRV32Config.fir@195463.12]
  wire  _GEN_257; // @[DCache.scala 750:45:freechips.rocketchip.system.DefaultRV32Config.fir@195455.10]
  wire  _GEN_267; // @[DCache.scala 748:36:freechips.rocketchip.system.DefaultRV32Config.fir@195450.8]
  wire  probeNack; // @[DCache.scala 746:28:freechips.rocketchip.system.DefaultRV32Config.fir@195446.6]
  reg [4:0] s1_req_cmd; // @[Reg.scala 15:16:freechips.rocketchip.system.DefaultRV32Config.fir@192231.4]
  wire  _T_30; // @[Consts.scala 82:31:freechips.rocketchip.system.DefaultRV32Config.fir@192264.4]
  wire  _T_31; // @[Consts.scala 82:48:freechips.rocketchip.system.DefaultRV32Config.fir@192265.4]
  wire  _T_32; // @[Consts.scala 82:41:freechips.rocketchip.system.DefaultRV32Config.fir@192266.4]
  wire  _T_33; // @[Consts.scala 82:65:freechips.rocketchip.system.DefaultRV32Config.fir@192267.4]
  wire  _T_34; // @[Consts.scala 82:58:freechips.rocketchip.system.DefaultRV32Config.fir@192268.4]
  wire  _T_35; // @[package.scala 15:47:freechips.rocketchip.system.DefaultRV32Config.fir@192269.4]
  wire  _T_36; // @[package.scala 15:47:freechips.rocketchip.system.DefaultRV32Config.fir@192270.4]
  wire  _T_39; // @[package.scala 64:59:freechips.rocketchip.system.DefaultRV32Config.fir@192273.4]
  wire  _T_37; // @[package.scala 15:47:freechips.rocketchip.system.DefaultRV32Config.fir@192271.4]
  wire  _T_40; // @[package.scala 64:59:freechips.rocketchip.system.DefaultRV32Config.fir@192274.4]
  wire  _T_38; // @[package.scala 15:47:freechips.rocketchip.system.DefaultRV32Config.fir@192272.4]
  wire  _T_41; // @[package.scala 64:59:freechips.rocketchip.system.DefaultRV32Config.fir@192275.4]
  wire  _T_42; // @[package.scala 15:47:freechips.rocketchip.system.DefaultRV32Config.fir@192276.4]
  wire  _T_43; // @[package.scala 15:47:freechips.rocketchip.system.DefaultRV32Config.fir@192277.4]
  wire  _T_47; // @[package.scala 64:59:freechips.rocketchip.system.DefaultRV32Config.fir@192281.4]
  wire  _T_44; // @[package.scala 15:47:freechips.rocketchip.system.DefaultRV32Config.fir@192278.4]
  wire  _T_48; // @[package.scala 64:59:freechips.rocketchip.system.DefaultRV32Config.fir@192282.4]
  wire  _T_45; // @[package.scala 15:47:freechips.rocketchip.system.DefaultRV32Config.fir@192279.4]
  wire  _T_49; // @[package.scala 64:59:freechips.rocketchip.system.DefaultRV32Config.fir@192283.4]
  wire  _T_46; // @[package.scala 15:47:freechips.rocketchip.system.DefaultRV32Config.fir@192280.4]
  wire  _T_50; // @[package.scala 64:59:freechips.rocketchip.system.DefaultRV32Config.fir@192284.4]
  wire  _T_51; // @[Consts.scala 80:44:freechips.rocketchip.system.DefaultRV32Config.fir@192285.4]
  wire  s1_read; // @[Consts.scala 82:75:freechips.rocketchip.system.DefaultRV32Config.fir@192286.4]
  reg [4:0] s2_req_cmd; // @[DCache.scala 291:19:freechips.rocketchip.system.DefaultRV32Config.fir@192778.4]
  wire  _T_402; // @[Consts.scala 83:32:freechips.rocketchip.system.DefaultRV32Config.fir@192828.4]
  wire  _T_403; // @[Consts.scala 83:49:freechips.rocketchip.system.DefaultRV32Config.fir@192829.4]
  wire  _T_404; // @[Consts.scala 83:42:freechips.rocketchip.system.DefaultRV32Config.fir@192830.4]
  wire  _T_405; // @[Consts.scala 83:66:freechips.rocketchip.system.DefaultRV32Config.fir@192831.4]
  wire  _T_406; // @[Consts.scala 83:59:freechips.rocketchip.system.DefaultRV32Config.fir@192832.4]
  wire  _T_407; // @[package.scala 15:47:freechips.rocketchip.system.DefaultRV32Config.fir@192833.4]
  wire  _T_408; // @[package.scala 15:47:freechips.rocketchip.system.DefaultRV32Config.fir@192834.4]
  wire  _T_411; // @[package.scala 64:59:freechips.rocketchip.system.DefaultRV32Config.fir@192837.4]
  wire  _T_409; // @[package.scala 15:47:freechips.rocketchip.system.DefaultRV32Config.fir@192835.4]
  wire  _T_412; // @[package.scala 64:59:freechips.rocketchip.system.DefaultRV32Config.fir@192838.4]
  wire  _T_410; // @[package.scala 15:47:freechips.rocketchip.system.DefaultRV32Config.fir@192836.4]
  wire  _T_413; // @[package.scala 64:59:freechips.rocketchip.system.DefaultRV32Config.fir@192839.4]
  wire  _T_414; // @[package.scala 15:47:freechips.rocketchip.system.DefaultRV32Config.fir@192840.4]
  wire  _T_415; // @[package.scala 15:47:freechips.rocketchip.system.DefaultRV32Config.fir@192841.4]
  wire  _T_419; // @[package.scala 64:59:freechips.rocketchip.system.DefaultRV32Config.fir@192845.4]
  wire  _T_416; // @[package.scala 15:47:freechips.rocketchip.system.DefaultRV32Config.fir@192842.4]
  wire  _T_420; // @[package.scala 64:59:freechips.rocketchip.system.DefaultRV32Config.fir@192846.4]
  wire  _T_417; // @[package.scala 15:47:freechips.rocketchip.system.DefaultRV32Config.fir@192843.4]
  wire  _T_421; // @[package.scala 64:59:freechips.rocketchip.system.DefaultRV32Config.fir@192847.4]
  wire  _T_418; // @[package.scala 15:47:freechips.rocketchip.system.DefaultRV32Config.fir@192844.4]
  wire  _T_422; // @[package.scala 64:59:freechips.rocketchip.system.DefaultRV32Config.fir@192848.4]
  wire  _T_423; // @[Consts.scala 80:44:freechips.rocketchip.system.DefaultRV32Config.fir@192849.4]
  wire  s2_write; // @[Consts.scala 83:76:freechips.rocketchip.system.DefaultRV32Config.fir@192850.4]
  wire  _T_977; // @[DCache.scala 456:39:freechips.rocketchip.system.DefaultRV32Config.fir@193647.4]
  reg  pstore1_held; // @[DCache.scala 455:25:freechips.rocketchip.system.DefaultRV32Config.fir@193646.4]
  wire  pstore1_valid_likely; // @[DCache.scala 456:51:freechips.rocketchip.system.DefaultRV32Config.fir@193648.4]
  reg [31:0] pstore1_addr; // @[Reg.scala 15:16:freechips.rocketchip.system.DefaultRV32Config.fir@193484.4]
  reg [31:0] s1_req_addr; // @[Reg.scala 15:16:freechips.rocketchip.system.DefaultRV32Config.fir@192231.4]
  wire  _T_1094; // @[DCache.scala 508:31:freechips.rocketchip.system.DefaultRV32Config.fir@193812.4]
  wire  _T_52; // @[Consts.scala 83:32:freechips.rocketchip.system.DefaultRV32Config.fir@192287.4]
  wire  _T_53; // @[Consts.scala 83:49:freechips.rocketchip.system.DefaultRV32Config.fir@192288.4]
  wire  _T_54; // @[Consts.scala 83:42:freechips.rocketchip.system.DefaultRV32Config.fir@192289.4]
  wire  _T_56; // @[Consts.scala 83:59:freechips.rocketchip.system.DefaultRV32Config.fir@192291.4]
  wire  s1_write; // @[Consts.scala 83:76:freechips.rocketchip.system.DefaultRV32Config.fir@192309.4]
  reg [3:0] pstore1_mask; // @[Reg.scala 15:16:freechips.rocketchip.system.DefaultRV32Config.fir@193499.4]
  wire  _T_1102; // @[DCache.scala 1076:66:freechips.rocketchip.system.DefaultRV32Config.fir@193820.4]
  wire  _T_1101; // @[DCache.scala 1076:66:freechips.rocketchip.system.DefaultRV32Config.fir@193819.4]
  wire  _T_1100; // @[DCache.scala 1076:66:freechips.rocketchip.system.DefaultRV32Config.fir@193818.4]
  wire  _T_1099; // @[DCache.scala 1076:66:freechips.rocketchip.system.DefaultRV32Config.fir@193817.4]
  wire [3:0] _T_1105; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@193823.4]
  wire [3:0] _T_1112; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@193830.4]
  reg [1:0] s1_req_size; // @[Reg.scala 15:16:freechips.rocketchip.system.DefaultRV32Config.fir@192231.4]
  wire  _T_332; // @[AMOALU.scala 17:57:freechips.rocketchip.system.DefaultRV32Config.fir@192724.4]
  wire  _T_334; // @[AMOALU.scala 17:46:freechips.rocketchip.system.DefaultRV32Config.fir@192726.4]
  wire  _T_336; // @[AMOALU.scala 18:22:freechips.rocketchip.system.DefaultRV32Config.fir@192728.4]
  wire [1:0] _T_337; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@192729.4]
  wire [1:0] _T_339; // @[AMOALU.scala 17:22:freechips.rocketchip.system.DefaultRV32Config.fir@192731.4]
  wire  _T_340; // @[AMOALU.scala 17:57:freechips.rocketchip.system.DefaultRV32Config.fir@192732.4]
  wire [1:0] _T_341; // @[AMOALU.scala 17:51:freechips.rocketchip.system.DefaultRV32Config.fir@192733.4]
  wire [1:0] _T_342; // @[AMOALU.scala 17:46:freechips.rocketchip.system.DefaultRV32Config.fir@192734.4]
  wire [1:0] _T_344; // @[AMOALU.scala 18:22:freechips.rocketchip.system.DefaultRV32Config.fir@192736.4]
  wire [3:0] s1_mask_xwr; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@192737.4]
  wire  _T_1120; // @[DCache.scala 1076:66:freechips.rocketchip.system.DefaultRV32Config.fir@193838.4]
  wire  _T_1119; // @[DCache.scala 1076:66:freechips.rocketchip.system.DefaultRV32Config.fir@193837.4]
  wire  _T_1118; // @[DCache.scala 1076:66:freechips.rocketchip.system.DefaultRV32Config.fir@193836.4]
  wire  _T_1117; // @[DCache.scala 1076:66:freechips.rocketchip.system.DefaultRV32Config.fir@193835.4]
  wire [3:0] _T_1123; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@193841.4]
  wire [3:0] _T_1130; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@193848.4]
  wire [3:0] _T_1131; // @[DCache.scala 509:38:freechips.rocketchip.system.DefaultRV32Config.fir@193849.4]
  wire  _T_1132; // @[DCache.scala 509:66:freechips.rocketchip.system.DefaultRV32Config.fir@193850.4]
  wire [3:0] _T_1133; // @[DCache.scala 509:77:freechips.rocketchip.system.DefaultRV32Config.fir@193851.4]
  wire  _T_1134; // @[DCache.scala 509:92:freechips.rocketchip.system.DefaultRV32Config.fir@193852.4]
  wire  _T_1135; // @[DCache.scala 509:8:freechips.rocketchip.system.DefaultRV32Config.fir@193853.4]
  wire  _T_1136; // @[DCache.scala 508:68:freechips.rocketchip.system.DefaultRV32Config.fir@193854.4]
  wire  _T_1137; // @[DCache.scala 511:27:freechips.rocketchip.system.DefaultRV32Config.fir@193855.4]
  reg  pstore2_valid; // @[DCache.scala 452:26:freechips.rocketchip.system.DefaultRV32Config.fir@193571.4]
  reg [31:0] pstore2_addr; // @[Reg.scala 15:16:freechips.rocketchip.system.DefaultRV32Config.fir@193710.4]
  wire  _T_1140; // @[DCache.scala 508:31:freechips.rocketchip.system.DefaultRV32Config.fir@193858.4]
  reg [3:0] mask; // @[DCache.scala 482:19:freechips.rocketchip.system.DefaultRV32Config.fir@193754.4]
  wire  _T_1148; // @[DCache.scala 1076:66:freechips.rocketchip.system.DefaultRV32Config.fir@193866.4]
  wire  _T_1147; // @[DCache.scala 1076:66:freechips.rocketchip.system.DefaultRV32Config.fir@193865.4]
  wire  _T_1146; // @[DCache.scala 1076:66:freechips.rocketchip.system.DefaultRV32Config.fir@193864.4]
  wire  _T_1145; // @[DCache.scala 1076:66:freechips.rocketchip.system.DefaultRV32Config.fir@193863.4]
  wire [3:0] _T_1151; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@193869.4]
  wire [3:0] _T_1158; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@193876.4]
  wire [3:0] _T_1177; // @[DCache.scala 509:38:freechips.rocketchip.system.DefaultRV32Config.fir@193895.4]
  wire  _T_1178; // @[DCache.scala 509:66:freechips.rocketchip.system.DefaultRV32Config.fir@193896.4]
  wire [3:0] _T_1179; // @[DCache.scala 509:77:freechips.rocketchip.system.DefaultRV32Config.fir@193897.4]
  wire  _T_1180; // @[DCache.scala 509:92:freechips.rocketchip.system.DefaultRV32Config.fir@193898.4]
  wire  _T_1181; // @[DCache.scala 509:8:freechips.rocketchip.system.DefaultRV32Config.fir@193899.4]
  wire  _T_1182; // @[DCache.scala 508:68:freechips.rocketchip.system.DefaultRV32Config.fir@193900.4]
  wire  _T_1183; // @[DCache.scala 512:21:freechips.rocketchip.system.DefaultRV32Config.fir@193901.4]
  wire  s1_hazard; // @[DCache.scala 511:69:freechips.rocketchip.system.DefaultRV32Config.fir@193902.4]
  wire  s1_raw_hazard; // @[DCache.scala 513:31:freechips.rocketchip.system.DefaultRV32Config.fir@193903.4]
  wire  _T_1184; // @[DCache.scala 518:18:freechips.rocketchip.system.DefaultRV32Config.fir@193905.4]
  wire [5:0] _T_362; // @[DCache.scala 284:54:freechips.rocketchip.system.DefaultRV32Config.fir@192762.4]
  wire  _T_363; // @[DCache.scala 284:61:freechips.rocketchip.system.DefaultRV32Config.fir@192763.4]
  wire  _T_364; // @[DCache.scala 284:38:freechips.rocketchip.system.DefaultRV32Config.fir@192764.4]
  wire  s2_valid_no_xcpt; // @[DCache.scala 284:35:freechips.rocketchip.system.DefaultRV32Config.fir@192765.4]
  reg  s2_not_nacked_in_s1; // @[DCache.scala 287:36:freechips.rocketchip.system.DefaultRV32Config.fir@192772.4]
  wire  s2_valid_masked; // @[DCache.scala 289:42:freechips.rocketchip.system.DefaultRV32Config.fir@192775.4]
  wire  _T_603; // @[DCache.scala 349:74:freechips.rocketchip.system.DefaultRV32Config.fir@193144.4]
  wire  _T_604; // @[DCache.scala 349:71:freechips.rocketchip.system.DefaultRV32Config.fir@193145.4]
  wire  _T_523; // @[Consts.scala 84:54:freechips.rocketchip.system.DefaultRV32Config.fir@193055.4]
  wire  _T_524; // @[Consts.scala 84:47:freechips.rocketchip.system.DefaultRV32Config.fir@193056.4]
  wire  _T_525; // @[Consts.scala 84:71:freechips.rocketchip.system.DefaultRV32Config.fir@193057.4]
  wire  _T_526; // @[Consts.scala 84:64:freechips.rocketchip.system.DefaultRV32Config.fir@193058.4]
  reg [1:0] s2_hit_state_state; // @[Reg.scala 15:16:freechips.rocketchip.system.DefaultRV32Config.fir@192998.4]
  wire [3:0] _T_528; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@193060.4]
  wire  _T_586; // @[Misc.scala 48:20:freechips.rocketchip.system.DefaultRV32Config.fir@193118.4]
  wire  _T_583; // @[Misc.scala 48:20:freechips.rocketchip.system.DefaultRV32Config.fir@193115.4]
  wire  _T_580; // @[Misc.scala 48:20:freechips.rocketchip.system.DefaultRV32Config.fir@193112.4]
  wire  _T_577; // @[Misc.scala 48:20:freechips.rocketchip.system.DefaultRV32Config.fir@193109.4]
  wire  _T_574; // @[Misc.scala 48:20:freechips.rocketchip.system.DefaultRV32Config.fir@193106.4]
  wire  _T_571; // @[Misc.scala 48:20:freechips.rocketchip.system.DefaultRV32Config.fir@193103.4]
  wire  _T_568; // @[Misc.scala 48:20:freechips.rocketchip.system.DefaultRV32Config.fir@193100.4]
  wire  _T_565; // @[Misc.scala 48:20:freechips.rocketchip.system.DefaultRV32Config.fir@193097.4]
  wire  _T_562; // @[Misc.scala 48:20:freechips.rocketchip.system.DefaultRV32Config.fir@193094.4]
  wire  _T_559; // @[Misc.scala 48:20:freechips.rocketchip.system.DefaultRV32Config.fir@193091.4]
  wire  _T_556; // @[Misc.scala 48:20:freechips.rocketchip.system.DefaultRV32Config.fir@193088.4]
  wire  _T_553; // @[Misc.scala 48:20:freechips.rocketchip.system.DefaultRV32Config.fir@193085.4]
  wire  _T_572; // @[Misc.scala 34:9:freechips.rocketchip.system.DefaultRV32Config.fir@193104.4]
  wire  _T_575; // @[Misc.scala 34:9:freechips.rocketchip.system.DefaultRV32Config.fir@193107.4]
  wire  _T_578; // @[Misc.scala 34:9:freechips.rocketchip.system.DefaultRV32Config.fir@193110.4]
  wire  _T_581; // @[Misc.scala 34:9:freechips.rocketchip.system.DefaultRV32Config.fir@193113.4]
  wire  _T_584; // @[Misc.scala 34:9:freechips.rocketchip.system.DefaultRV32Config.fir@193116.4]
  wire  s2_hit; // @[Misc.scala 34:9:freechips.rocketchip.system.DefaultRV32Config.fir@193119.4]
  wire  s2_valid_hit_maybe_flush_pre_data_ecc_and_waw; // @[DCache.scala 349:89:freechips.rocketchip.system.DefaultRV32Config.fir@193146.4]
  wire  _T_380; // @[Consts.scala 82:31:freechips.rocketchip.system.DefaultRV32Config.fir@192805.4]
  wire  _T_382; // @[Consts.scala 82:41:freechips.rocketchip.system.DefaultRV32Config.fir@192807.4]
  wire  _T_384; // @[Consts.scala 82:58:freechips.rocketchip.system.DefaultRV32Config.fir@192809.4]
  wire  s2_read; // @[Consts.scala 82:75:freechips.rocketchip.system.DefaultRV32Config.fir@192827.4]
  wire  s2_readwrite; // @[DCache.scala 306:30:freechips.rocketchip.system.DefaultRV32Config.fir@192851.4]
  wire  s2_valid_hit_pre_data_ecc_and_waw; // @[DCache.scala 370:89:freechips.rocketchip.system.DefaultRV32Config.fir@193147.4]
  wire [1:0] _T_555; // @[Misc.scala 34:36:freechips.rocketchip.system.DefaultRV32Config.fir@193087.4]
  wire [1:0] _T_558; // @[Misc.scala 34:36:freechips.rocketchip.system.DefaultRV32Config.fir@193090.4]
  wire [1:0] _T_561; // @[Misc.scala 34:36:freechips.rocketchip.system.DefaultRV32Config.fir@193093.4]
  wire [1:0] _T_564; // @[Misc.scala 34:36:freechips.rocketchip.system.DefaultRV32Config.fir@193096.4]
  wire [1:0] _T_567; // @[Misc.scala 34:36:freechips.rocketchip.system.DefaultRV32Config.fir@193099.4]
  wire [1:0] _T_570; // @[Misc.scala 34:36:freechips.rocketchip.system.DefaultRV32Config.fir@193102.4]
  wire [1:0] _T_573; // @[Misc.scala 34:36:freechips.rocketchip.system.DefaultRV32Config.fir@193105.4]
  wire [1:0] _T_576; // @[Misc.scala 34:36:freechips.rocketchip.system.DefaultRV32Config.fir@193108.4]
  wire [1:0] _T_579; // @[Misc.scala 34:36:freechips.rocketchip.system.DefaultRV32Config.fir@193111.4]
  wire [1:0] _T_582; // @[Misc.scala 34:36:freechips.rocketchip.system.DefaultRV32Config.fir@193114.4]
  wire [1:0] _T_585; // @[Misc.scala 34:36:freechips.rocketchip.system.DefaultRV32Config.fir@193117.4]
  wire [1:0] s2_grow_param; // @[Misc.scala 34:36:freechips.rocketchip.system.DefaultRV32Config.fir@193120.4]
  wire  _T_764; // @[Metadata.scala 46:46:freechips.rocketchip.system.DefaultRV32Config.fir@193340.4]
  wire  s2_update_meta; // @[Metadata.scala 47:40:freechips.rocketchip.system.DefaultRV32Config.fir@193341.4]
  wire  _T_783; // @[DCache.scala 397:62:freechips.rocketchip.system.DefaultRV32Config.fir@193363.4]
  wire  _T_784; // @[DCache.scala 397:24:freechips.rocketchip.system.DefaultRV32Config.fir@193364.4]
  wire  s1_readwrite; // @[DCache.scala 185:30:freechips.rocketchip.system.DefaultRV32Config.fir@192310.4]
  wire  _T_74; // @[DCache.scala 187:34:freechips.rocketchip.system.DefaultRV32Config.fir@192312.4]
  wire  s1_flush_line; // @[DCache.scala 187:50:freechips.rocketchip.system.DefaultRV32Config.fir@192314.4]
  wire  _T_227; // @[DCache.scala 229:38:freechips.rocketchip.system.DefaultRV32Config.fir@192517.4]
  wire  _T_228; // @[DCache.scala 229:69:freechips.rocketchip.system.DefaultRV32Config.fir@192518.4]
  wire  s1_cmd_uses_tlb; // @[DCache.scala 229:55:freechips.rocketchip.system.DefaultRV32Config.fir@192519.4]
  wire  _T_242; // @[DCache.scala 235:39:freechips.rocketchip.system.DefaultRV32Config.fir@192540.4]
  wire  _T_243; // @[DCache.scala 235:58:freechips.rocketchip.system.DefaultRV32Config.fir@192541.4]
  wire  _GEN_118; // @[DCache.scala 397:82:freechips.rocketchip.system.DefaultRV32Config.fir@193365.4]
  wire  _GEN_138; // @[DCache.scala 518:36:freechips.rocketchip.system.DefaultRV32Config.fir@193906.4]
  wire  _GEN_278; // @[DCache.scala 759:24:freechips.rocketchip.system.DefaultRV32Config.fir@195468.6]
  wire  s1_nack; // @[DCache.scala 744:21:freechips.rocketchip.system.DefaultRV32Config.fir@195442.4]
  wire  _T_20; // @[DCache.scala 164:41:freechips.rocketchip.system.DefaultRV32Config.fir@192211.4]
  wire  s1_valid_not_nacked; // @[DCache.scala 164:38:freechips.rocketchip.system.DefaultRV32Config.fir@192212.4]
  wire  _T_22; // @[DCache.scala 167:43:freechips.rocketchip.system.DefaultRV32Config.fir@192218.4]
  wire  s0_clk_en; // @[DCache.scala 167:40:freechips.rocketchip.system.DefaultRV32Config.fir@192219.4]
  wire [31:0] s0_req_addr; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@192225.4]
  wire  _T_26; // @[DCache.scala 171:9:freechips.rocketchip.system.DefaultRV32Config.fir@192227.4]
  wire  s0_req_phys; // @[DCache.scala 171:34:freechips.rocketchip.system.DefaultRV32Config.fir@192228.4]
  reg [6:0] s1_req_tag; // @[Reg.scala 15:16:freechips.rocketchip.system.DefaultRV32Config.fir@192231.4]
  reg  s1_req_signed; // @[Reg.scala 15:16:freechips.rocketchip.system.DefaultRV32Config.fir@192231.4]
  reg [1:0] s1_req_dprv; // @[Reg.scala 15:16:freechips.rocketchip.system.DefaultRV32Config.fir@192231.4]
  reg [31:0] s1_tlb_req_vaddr; // @[Reg.scala 15:16:freechips.rocketchip.system.DefaultRV32Config.fir@192257.4]
  reg  s1_tlb_req_passthrough; // @[Reg.scala 15:16:freechips.rocketchip.system.DefaultRV32Config.fir@192257.4]
  reg [1:0] s1_tlb_req_size; // @[Reg.scala 15:16:freechips.rocketchip.system.DefaultRV32Config.fir@192257.4]
  reg [4:0] s1_tlb_req_cmd; // @[Reg.scala 15:16:freechips.rocketchip.system.DefaultRV32Config.fir@192257.4]
  wire  s1_sfence; // @[DCache.scala 186:30:freechips.rocketchip.system.DefaultRV32Config.fir@192311.4]
  reg  cached_grant_wait; // @[DCache.scala 196:30:freechips.rocketchip.system.DefaultRV32Config.fir@192321.4]
  wire  inWriteback; // @[package.scala 64:59:freechips.rocketchip.system.DefaultRV32Config.fir@192329.4]
  wire  _T_78; // @[DCache.scala 203:38:freechips.rocketchip.system.DefaultRV32Config.fir@192332.4]
  wire  _T_79; // @[DCache.scala 203:54:freechips.rocketchip.system.DefaultRV32Config.fir@192333.4]
  wire  _T_80; // @[DCache.scala 203:51:freechips.rocketchip.system.DefaultRV32Config.fir@192334.4]
  wire  _T_82; // @[DCache.scala 203:73:freechips.rocketchip.system.DefaultRV32Config.fir@192336.4]
  reg  uncachedInFlight_0; // @[DCache.scala 206:33:freechips.rocketchip.system.DefaultRV32Config.fir@192341.4]
  reg [31:0] uncachedReqs_0_addr; // @[DCache.scala 207:25:freechips.rocketchip.system.DefaultRV32Config.fir@192342.4]
  reg [6:0] uncachedReqs_0_tag; // @[DCache.scala 207:25:freechips.rocketchip.system.DefaultRV32Config.fir@192342.4]
  reg [1:0] uncachedReqs_0_size; // @[DCache.scala 207:25:freechips.rocketchip.system.DefaultRV32Config.fir@192342.4]
  reg  uncachedReqs_0_signed; // @[DCache.scala 207:25:freechips.rocketchip.system.DefaultRV32Config.fir@192342.4]
  wire  _T_84; // @[Consts.scala 82:31:freechips.rocketchip.system.DefaultRV32Config.fir@192346.4]
  wire  _T_85; // @[Consts.scala 82:48:freechips.rocketchip.system.DefaultRV32Config.fir@192347.4]
  wire  _T_86; // @[Consts.scala 82:41:freechips.rocketchip.system.DefaultRV32Config.fir@192348.4]
  wire  _T_87; // @[Consts.scala 82:65:freechips.rocketchip.system.DefaultRV32Config.fir@192349.4]
  wire  _T_88; // @[Consts.scala 82:58:freechips.rocketchip.system.DefaultRV32Config.fir@192350.4]
  wire  _T_89; // @[package.scala 15:47:freechips.rocketchip.system.DefaultRV32Config.fir@192351.4]
  wire  _T_90; // @[package.scala 15:47:freechips.rocketchip.system.DefaultRV32Config.fir@192352.4]
  wire  _T_91; // @[package.scala 15:47:freechips.rocketchip.system.DefaultRV32Config.fir@192353.4]
  wire  _T_92; // @[package.scala 15:47:freechips.rocketchip.system.DefaultRV32Config.fir@192354.4]
  wire  _T_93; // @[package.scala 64:59:freechips.rocketchip.system.DefaultRV32Config.fir@192355.4]
  wire  _T_94; // @[package.scala 64:59:freechips.rocketchip.system.DefaultRV32Config.fir@192356.4]
  wire  _T_95; // @[package.scala 64:59:freechips.rocketchip.system.DefaultRV32Config.fir@192357.4]
  wire  _T_96; // @[package.scala 15:47:freechips.rocketchip.system.DefaultRV32Config.fir@192358.4]
  wire  _T_97; // @[package.scala 15:47:freechips.rocketchip.system.DefaultRV32Config.fir@192359.4]
  wire  _T_98; // @[package.scala 15:47:freechips.rocketchip.system.DefaultRV32Config.fir@192360.4]
  wire  _T_99; // @[package.scala 15:47:freechips.rocketchip.system.DefaultRV32Config.fir@192361.4]
  wire  _T_100; // @[package.scala 15:47:freechips.rocketchip.system.DefaultRV32Config.fir@192362.4]
  wire  _T_101; // @[package.scala 64:59:freechips.rocketchip.system.DefaultRV32Config.fir@192363.4]
  wire  _T_102; // @[package.scala 64:59:freechips.rocketchip.system.DefaultRV32Config.fir@192364.4]
  wire  _T_103; // @[package.scala 64:59:freechips.rocketchip.system.DefaultRV32Config.fir@192365.4]
  wire  _T_104; // @[package.scala 64:59:freechips.rocketchip.system.DefaultRV32Config.fir@192366.4]
  wire  _T_105; // @[Consts.scala 80:44:freechips.rocketchip.system.DefaultRV32Config.fir@192367.4]
  wire  s0_read; // @[Consts.scala 82:75:freechips.rocketchip.system.DefaultRV32Config.fir@192368.4]
  wire  _T_106; // @[package.scala 15:47:freechips.rocketchip.system.DefaultRV32Config.fir@192369.4]
  wire  _T_107; // @[package.scala 15:47:freechips.rocketchip.system.DefaultRV32Config.fir@192370.4]
  wire  _T_108; // @[package.scala 64:59:freechips.rocketchip.system.DefaultRV32Config.fir@192371.4]
  wire  res; // @[DCache.scala 1080:15:freechips.rocketchip.system.DefaultRV32Config.fir@192372.4]
  wire  _T_135; // @[Consts.scala 83:49:freechips.rocketchip.system.DefaultRV32Config.fir@192399.4]
  wire  _T_136; // @[Consts.scala 83:42:freechips.rocketchip.system.DefaultRV32Config.fir@192400.4]
  wire  _T_138; // @[Consts.scala 83:59:freechips.rocketchip.system.DefaultRV32Config.fir@192402.4]
  wire  _T_156; // @[Consts.scala 83:76:freechips.rocketchip.system.DefaultRV32Config.fir@192420.4]
  wire  _T_160; // @[DCache.scala 1086:23:freechips.rocketchip.system.DefaultRV32Config.fir@192424.4]
  wire  _T_161; // @[DCache.scala 1085:21:freechips.rocketchip.system.DefaultRV32Config.fir@192425.4]
  wire  _T_162; // @[DCache.scala 1081:12:freechips.rocketchip.system.DefaultRV32Config.fir@192426.4]
  wire  _T_163; // @[DCache.scala 1081:28:freechips.rocketchip.system.DefaultRV32Config.fir@192427.4]
  wire  _T_165; // @[DCache.scala 1081:11:freechips.rocketchip.system.DefaultRV32Config.fir@192429.4]
  wire  _T_166; // @[DCache.scala 1081:11:freechips.rocketchip.system.DefaultRV32Config.fir@192430.4]
  wire  _T_167; // @[DCache.scala 212:46:freechips.rocketchip.system.DefaultRV32Config.fir@192435.4]
  wire  _T_170; // @[DCache.scala 218:9:freechips.rocketchip.system.DefaultRV32Config.fir@192444.4]
  wire  _T_171; // @[DCache.scala 218:33:freechips.rocketchip.system.DefaultRV32Config.fir@192445.4]
  wire  _GEN_28; // @[DCache.scala 218:45:freechips.rocketchip.system.DefaultRV32Config.fir@192446.4]
  wire  _T_223; // @[DCache.scala 219:75:freechips.rocketchip.system.DefaultRV32Config.fir@192500.4]
  wire  _T_224; // @[DCache.scala 219:54:freechips.rocketchip.system.DefaultRV32Config.fir@192501.4]
  reg  s1_did_read; // @[Reg.scala 15:16:freechips.rocketchip.system.DefaultRV32Config.fir@192502.4]
  wire  _GEN_30; // @[DCache.scala 226:34:freechips.rocketchip.system.DefaultRV32Config.fir@192514.4]
  wire  _T_235; // @[DCache.scala 234:9:freechips.rocketchip.system.DefaultRV32Config.fir@192530.4]
  wire  _T_236; // @[DCache.scala 234:30:freechips.rocketchip.system.DefaultRV32Config.fir@192531.4]
  wire  _T_237; // @[DCache.scala 234:27:freechips.rocketchip.system.DefaultRV32Config.fir@192532.4]
  wire  _T_238; // @[DCache.scala 234:56:freechips.rocketchip.system.DefaultRV32Config.fir@192533.4]
  wire  _T_239; // @[DCache.scala 234:53:freechips.rocketchip.system.DefaultRV32Config.fir@192534.4]
  wire  _GEN_31; // @[DCache.scala 234:79:freechips.rocketchip.system.DefaultRV32Config.fir@192535.4]
  wire [31:0] s1_paddr; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@192570.4]
  wire [1:0] s1_victim_way; // @[package.scala 138:13:freechips.rocketchip.system.DefaultRV32Config.fir@192571.4]
  wire  _T_258; // @[DCache.scala 262:27:freechips.rocketchip.system.DefaultRV32Config.fir@192575.4]
  wire [21:0] _T_266; // @[:freechips.rocketchip.system.DefaultRV32Config.fir@192614.4 :freechips.rocketchip.system.DefaultRV32Config.fir@192616.4]
  wire [19:0] s1_meta_uncorrected_0_tag; // @[DCache.scala 267:80:freechips.rocketchip.system.DefaultRV32Config.fir@192617.4]
  wire [1:0] s1_meta_uncorrected_0_coh_state; // @[DCache.scala 267:80:freechips.rocketchip.system.DefaultRV32Config.fir@192619.4]
  wire [21:0] _T_269; // @[:freechips.rocketchip.system.DefaultRV32Config.fir@192623.4 :freechips.rocketchip.system.DefaultRV32Config.fir@192625.4]
  wire [19:0] s1_meta_uncorrected_1_tag; // @[DCache.scala 267:80:freechips.rocketchip.system.DefaultRV32Config.fir@192626.4]
  wire [1:0] s1_meta_uncorrected_1_coh_state; // @[DCache.scala 267:80:freechips.rocketchip.system.DefaultRV32Config.fir@192628.4]
  wire [21:0] _T_272; // @[:freechips.rocketchip.system.DefaultRV32Config.fir@192632.4 :freechips.rocketchip.system.DefaultRV32Config.fir@192634.4]
  wire [19:0] s1_meta_uncorrected_2_tag; // @[DCache.scala 267:80:freechips.rocketchip.system.DefaultRV32Config.fir@192635.4]
  wire [1:0] s1_meta_uncorrected_2_coh_state; // @[DCache.scala 267:80:freechips.rocketchip.system.DefaultRV32Config.fir@192637.4]
  wire [21:0] _T_275; // @[:freechips.rocketchip.system.DefaultRV32Config.fir@192641.4 :freechips.rocketchip.system.DefaultRV32Config.fir@192643.4]
  wire [19:0] s1_meta_uncorrected_3_tag; // @[DCache.scala 267:80:freechips.rocketchip.system.DefaultRV32Config.fir@192644.4]
  wire [1:0] s1_meta_uncorrected_3_coh_state; // @[DCache.scala 267:80:freechips.rocketchip.system.DefaultRV32Config.fir@192646.4]
  wire [19:0] s1_tag; // @[DCache.scala 268:29:freechips.rocketchip.system.DefaultRV32Config.fir@192648.4]
  wire  _T_278; // @[Metadata.scala 50:45:freechips.rocketchip.system.DefaultRV32Config.fir@192649.4]
  wire  _T_279; // @[DCache.scala 269:83:freechips.rocketchip.system.DefaultRV32Config.fir@192650.4]
  wire  _T_280; // @[DCache.scala 269:74:freechips.rocketchip.system.DefaultRV32Config.fir@192651.4]
  wire  _T_281; // @[Metadata.scala 50:45:freechips.rocketchip.system.DefaultRV32Config.fir@192652.4]
  wire  _T_282; // @[DCache.scala 269:83:freechips.rocketchip.system.DefaultRV32Config.fir@192653.4]
  wire  _T_283; // @[DCache.scala 269:74:freechips.rocketchip.system.DefaultRV32Config.fir@192654.4]
  wire  _T_284; // @[Metadata.scala 50:45:freechips.rocketchip.system.DefaultRV32Config.fir@192655.4]
  wire  _T_285; // @[DCache.scala 269:83:freechips.rocketchip.system.DefaultRV32Config.fir@192656.4]
  wire  _T_286; // @[DCache.scala 269:74:freechips.rocketchip.system.DefaultRV32Config.fir@192657.4]
  wire  _T_287; // @[Metadata.scala 50:45:freechips.rocketchip.system.DefaultRV32Config.fir@192658.4]
  wire  _T_288; // @[DCache.scala 269:83:freechips.rocketchip.system.DefaultRV32Config.fir@192659.4]
  wire  _T_289; // @[DCache.scala 269:74:freechips.rocketchip.system.DefaultRV32Config.fir@192660.4]
  wire [3:0] s1_meta_hit_way; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@192663.4]
  wire [1:0] _T_296; // @[DCache.scala 271:41:freechips.rocketchip.system.DefaultRV32Config.fir@192670.4]
  wire [1:0] _T_300; // @[DCache.scala 271:41:freechips.rocketchip.system.DefaultRV32Config.fir@192674.4]
  wire [1:0] _T_304; // @[DCache.scala 271:41:freechips.rocketchip.system.DefaultRV32Config.fir@192678.4]
  wire [1:0] _T_308; // @[DCache.scala 271:41:freechips.rocketchip.system.DefaultRV32Config.fir@192682.4]
  wire [1:0] _T_309; // @[DCache.scala 272:19:freechips.rocketchip.system.DefaultRV32Config.fir@192683.4]
  wire [1:0] _T_310; // @[DCache.scala 272:19:freechips.rocketchip.system.DefaultRV32Config.fir@192684.4]
  wire [1:0] s1_meta_hit_state_state; // @[DCache.scala 272:19:freechips.rocketchip.system.DefaultRV32Config.fir@192685.4]
  wire  _T_316; // @[package.scala 32:86:freechips.rocketchip.system.DefaultRV32Config.fir@192695.4]
  wire  _T_318; // @[package.scala 32:86:freechips.rocketchip.system.DefaultRV32Config.fir@192697.4]
  wire  _T_320; // @[package.scala 32:86:freechips.rocketchip.system.DefaultRV32Config.fir@192699.4]
  wire  s2_hit_valid; // @[Metadata.scala 50:45:freechips.rocketchip.system.DefaultRV32Config.fir@193008.4]
  reg [3:0] s2_hit_way; // @[Reg.scala 15:16:freechips.rocketchip.system.DefaultRV32Config.fir@192993.4]
  reg [1:0] _T_632; // @[Reg.scala 15:16:freechips.rocketchip.system.DefaultRV32Config.fir@193186.4]
  wire [3:0] _T_633; // @[OneHot.scala 58:35:freechips.rocketchip.system.DefaultRV32Config.fir@193190.4]
  wire [3:0] s2_victim_way; // @[DCache.scala 383:26:freechips.rocketchip.system.DefaultRV32Config.fir@193191.4]
  reg [3:0] s2_probe_way; // @[Reg.scala 15:16:freechips.rocketchip.system.DefaultRV32Config.fir@192985.4]
  wire [3:0] releaseWay; // @[DCache.scala 783:81:freechips.rocketchip.system.DefaultRV32Config.fir@195510.4]
  wire [3:0] _T_321; // @[DCache.scala 275:61:freechips.rocketchip.system.DefaultRV32Config.fir@192701.4]
  wire [15:0] _T_326; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@192709.4]
  wire [15:0] _T_327; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@192710.4]
  wire [31:0] _T_328; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@192711.4]
  wire  _T_347; // @[DCache.scala 281:28:freechips.rocketchip.system.DefaultRV32Config.fir@192741.4]
  wire  _T_348; // @[DCache.scala 281:10:freechips.rocketchip.system.DefaultRV32Config.fir@192742.4]
  wire [3:0] _T_349; // @[DCache.scala 281:71:freechips.rocketchip.system.DefaultRV32Config.fir@192743.4]
  wire [3:0] _T_350; // @[DCache.scala 281:69:freechips.rocketchip.system.DefaultRV32Config.fir@192744.4]
  wire  _T_351; // @[DCache.scala 281:93:freechips.rocketchip.system.DefaultRV32Config.fir@192745.4]
  wire  _T_352; // @[DCache.scala 281:53:freechips.rocketchip.system.DefaultRV32Config.fir@192746.4]
  wire  _T_354; // @[DCache.scala 281:9:freechips.rocketchip.system.DefaultRV32Config.fir@192748.4]
  wire  _T_355; // @[DCache.scala 281:9:freechips.rocketchip.system.DefaultRV32Config.fir@192749.4]
  wire  _T_356; // @[DCache.scala 283:46:freechips.rocketchip.system.DefaultRV32Config.fir@192754.4]
  wire  _T_357; // @[DCache.scala 283:43:freechips.rocketchip.system.DefaultRV32Config.fir@192755.4]
  reg [31:0] s2_req_addr; // @[DCache.scala 291:19:freechips.rocketchip.system.DefaultRV32Config.fir@192778.4]
  reg [6:0] s2_req_tag; // @[DCache.scala 291:19:freechips.rocketchip.system.DefaultRV32Config.fir@192778.4]
  reg [1:0] s2_req_size; // @[DCache.scala 291:19:freechips.rocketchip.system.DefaultRV32Config.fir@192778.4]
  reg  s2_req_signed; // @[DCache.scala 291:19:freechips.rocketchip.system.DefaultRV32Config.fir@192778.4]
  reg [1:0] s2_req_dprv; // @[DCache.scala 291:19:freechips.rocketchip.system.DefaultRV32Config.fir@192778.4]
  wire  _T_369; // @[DCache.scala 292:37:freechips.rocketchip.system.DefaultRV32Config.fir@192779.4]
  wire  s2_cmd_flush_line; // @[DCache.scala 293:54:freechips.rocketchip.system.DefaultRV32Config.fir@192785.4]
  reg  s2_tlb_xcpt_pf_ld; // @[DCache.scala 294:24:freechips.rocketchip.system.DefaultRV32Config.fir@192786.4]
  reg  s2_tlb_xcpt_pf_st; // @[DCache.scala 294:24:freechips.rocketchip.system.DefaultRV32Config.fir@192786.4]
  reg  s2_tlb_xcpt_ae_ld; // @[DCache.scala 294:24:freechips.rocketchip.system.DefaultRV32Config.fir@192786.4]
  reg  s2_tlb_xcpt_ae_st; // @[DCache.scala 294:24:freechips.rocketchip.system.DefaultRV32Config.fir@192786.4]
  reg  s2_tlb_xcpt_ma_ld; // @[DCache.scala 294:24:freechips.rocketchip.system.DefaultRV32Config.fir@192786.4]
  reg  s2_tlb_xcpt_ma_st; // @[DCache.scala 294:24:freechips.rocketchip.system.DefaultRV32Config.fir@192786.4]
  reg  s2_pma_cacheable; // @[DCache.scala 295:19:freechips.rocketchip.system.DefaultRV32Config.fir@192787.4]
  reg [31:0] s2_uncached_resp_addr; // @[DCache.scala 296:34:freechips.rocketchip.system.DefaultRV32Config.fir@192788.4]
  reg [31:0] _T_377; // @[Reg.scala 15:16:freechips.rocketchip.system.DefaultRV32Config.fir@192798.4]
  wire [31:0] s2_vaddr; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@192804.4]
  wire  s1_meta_clk_en; // @[DCache.scala 309:62:freechips.rocketchip.system.DefaultRV32Config.fir@192855.4]
  reg [21:0] _T_449; // @[Reg.scala 15:16:freechips.rocketchip.system.DefaultRV32Config.fir@192934.4]
  wire [19:0] s2_meta_corrected_3_tag; // @[DCache.scala 313:99:freechips.rocketchip.system.DefaultRV32Config.fir@192943.4]
  wire [1:0] s2_meta_corrected_3_coh_state; // @[DCache.scala 313:99:freechips.rocketchip.system.DefaultRV32Config.fir@192945.4]
  wire  _T_455; // @[DCache.scala 318:23:freechips.rocketchip.system.DefaultRV32Config.fir@192951.4]
  wire  en; // @[DCache.scala 318:38:freechips.rocketchip.system.DefaultRV32Config.fir@192952.4]
  wire  _T_456; // @[DCache.scala 319:64:freechips.rocketchip.system.DefaultRV32Config.fir@192953.4]
  wire  _T_457; // @[DCache.scala 319:63:freechips.rocketchip.system.DefaultRV32Config.fir@192954.4]
  wire  word_en; // @[DCache.scala 319:22:freechips.rocketchip.system.DefaultRV32Config.fir@192955.4]
  wire [31:0] s1_all_data_ways_0; // @[DCache.scala 277:29:freechips.rocketchip.system.DefaultRV32Config.fir@192714.4 DCache.scala 277:29:freechips.rocketchip.system.DefaultRV32Config.fir@192716.4]
  wire [31:0] s1_all_data_ways_1; // @[DCache.scala 277:29:freechips.rocketchip.system.DefaultRV32Config.fir@192714.4 DCache.scala 277:29:freechips.rocketchip.system.DefaultRV32Config.fir@192717.4]
  wire [31:0] s1_all_data_ways_2; // @[DCache.scala 277:29:freechips.rocketchip.system.DefaultRV32Config.fir@192714.4 DCache.scala 277:29:freechips.rocketchip.system.DefaultRV32Config.fir@192718.4]
  wire [31:0] s1_all_data_ways_3; // @[DCache.scala 277:29:freechips.rocketchip.system.DefaultRV32Config.fir@192714.4 DCache.scala 277:29:freechips.rocketchip.system.DefaultRV32Config.fir@192719.4]
  wire  _T_458; // @[DCache.scala 329:28:freechips.rocketchip.system.DefaultRV32Config.fir@192961.4]
  wire  s1_word_en; // @[DCache.scala 329:27:freechips.rocketchip.system.DefaultRV32Config.fir@192962.4]
  wire  grantIsUncachedData; // @[package.scala 15:47:freechips.rocketchip.system.DefaultRV32Config.fir@195063.4]
  reg  blockUncachedGrant; // @[DCache.scala 693:33:freechips.rocketchip.system.DefaultRV32Config.fir@195294.4]
  wire  _T_2333; // @[DCache.scala 695:54:freechips.rocketchip.system.DefaultRV32Config.fir@195296.4]
  wire  _T_2334; // @[DCache.scala 695:31:freechips.rocketchip.system.DefaultRV32Config.fir@195297.4]
  wire  grantIsRefill; // @[DCache.scala 609:29:freechips.rocketchip.system.DefaultRV32Config.fir@195081.4]
  wire  _T_2247; // @[DCache.scala 665:26:freechips.rocketchip.system.DefaultRV32Config.fir@195187.4]
  wire  _T_2248; // @[DCache.scala 665:23:freechips.rocketchip.system.DefaultRV32Config.fir@195188.4]
  wire  _T_2201; // @[package.scala 15:47:freechips.rocketchip.system.DefaultRV32Config.fir@195077.4]
  wire  grantIsCached; // @[package.scala 64:59:freechips.rocketchip.system.DefaultRV32Config.fir@195079.4]
  reg [9:0] _T_2177; // @[Edges.scala 230:27:freechips.rocketchip.system.DefaultRV32Config.fir@195043.4]
  wire  d_first; // @[Edges.scala 232:25:freechips.rocketchip.system.DefaultRV32Config.fir@195046.4]
  wire  _T_2209; // @[DCache.scala 614:41:freechips.rocketchip.system.DefaultRV32Config.fir@195094.4]
  wire  _T_2210; // @[DCache.scala 614:50:freechips.rocketchip.system.DefaultRV32Config.fir@195095.4]
  wire  canAcceptCachedGrant; // @[DCache.scala 613:30:freechips.rocketchip.system.DefaultRV32Config.fir@195093.4]
  wire  _T_2211; // @[DCache.scala 614:69:freechips.rocketchip.system.DefaultRV32Config.fir@195096.4]
  wire  _T_2212; // @[DCache.scala 614:24:freechips.rocketchip.system.DefaultRV32Config.fir@195097.4]
  wire  _GEN_228; // @[DCache.scala 665:51:freechips.rocketchip.system.DefaultRV32Config.fir@195189.4]
  wire  tl_out__d_ready; // @[DCache.scala 695:68:freechips.rocketchip.system.DefaultRV32Config.fir@195298.4]
  wire  _T_2217; // @[Decoupled.scala 40:37:freechips.rocketchip.system.DefaultRV32Config.fir@195105.4]
  wire  _T_2186; // @[package.scala 15:47:freechips.rocketchip.system.DefaultRV32Config.fir@195059.4]
  wire  _T_2188; // @[package.scala 64:59:freechips.rocketchip.system.DefaultRV32Config.fir@195061.4]
  wire  _T_2187; // @[package.scala 15:47:freechips.rocketchip.system.DefaultRV32Config.fir@195060.4]
  wire  grantIsUncached; // @[package.scala 64:59:freechips.rocketchip.system.DefaultRV32Config.fir@195062.4]
  wire [4:0] _GEN_184; // @[DCache.scala 634:34:freechips.rocketchip.system.DefaultRV32Config.fir@195137.10]
  wire [4:0] _GEN_193; // @[DCache.scala 627:35:freechips.rocketchip.system.DefaultRV32Config.fir@195124.8]
  wire [4:0] _GEN_206; // @[DCache.scala 618:26:freechips.rocketchip.system.DefaultRV32Config.fir@195107.6]
  wire [4:0] s1_data_way; // @[DCache.scala 617:26:freechips.rocketchip.system.DefaultRV32Config.fir@195106.4]
  wire [4:0] _T_460; // @[DCache.scala 331:28:freechips.rocketchip.system.DefaultRV32Config.fir@192964.4]
  wire [31:0] _T_466; // @[Mux.scala 27:72:freechips.rocketchip.system.DefaultRV32Config.fir@192970.4]
  wire [31:0] _T_467; // @[Mux.scala 27:72:freechips.rocketchip.system.DefaultRV32Config.fir@192971.4]
  wire [31:0] _T_468; // @[Mux.scala 27:72:freechips.rocketchip.system.DefaultRV32Config.fir@192972.4]
  wire [31:0] _T_469; // @[Mux.scala 27:72:freechips.rocketchip.system.DefaultRV32Config.fir@192973.4]
  wire [31:0] _T_470; // @[Mux.scala 27:72:freechips.rocketchip.system.DefaultRV32Config.fir@192974.4]
  wire [31:0] _T_471; // @[Mux.scala 27:72:freechips.rocketchip.system.DefaultRV32Config.fir@192975.4]
  wire [31:0] _T_472; // @[Mux.scala 27:72:freechips.rocketchip.system.DefaultRV32Config.fir@192976.4]
  wire [31:0] _T_473; // @[Mux.scala 27:72:freechips.rocketchip.system.DefaultRV32Config.fir@192977.4]
  wire [31:0] _T_474; // @[Mux.scala 27:72:freechips.rocketchip.system.DefaultRV32Config.fir@192978.4]
  reg [31:0] s2_data; // @[Reg.scala 15:16:freechips.rocketchip.system.DefaultRV32Config.fir@192981.4]
  wire [15:0] _T_599; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@193138.4]
  wire [15:0] _T_600; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@193139.4]
  wire [31:0] s2_data_corrected; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@193140.4]
  wire  s2_valid_flush_line; // @[DCache.scala 371:75:freechips.rocketchip.system.DefaultRV32Config.fir@193150.4]
  wire  _T_610; // @[DCache.scala 375:39:freechips.rocketchip.system.DefaultRV32Config.fir@193157.4]
  wire  _T_612; // @[DCache.scala 375:55:freechips.rocketchip.system.DefaultRV32Config.fir@193159.4]
  wire  _T_613; // @[DCache.scala 375:76:freechips.rocketchip.system.DefaultRV32Config.fir@193160.4]
  wire  s2_valid_miss; // @[DCache.scala 375:73:freechips.rocketchip.system.DefaultRV32Config.fir@193161.4]
  wire  s2_uncached; // @[DCache.scala 376:21:freechips.rocketchip.system.DefaultRV32Config.fir@193162.4]
  wire  _T_619; // @[DCache.scala 377:47:freechips.rocketchip.system.DefaultRV32Config.fir@193168.4]
  wire  _T_620; // @[DCache.scala 377:44:freechips.rocketchip.system.DefaultRV32Config.fir@193169.4]
  wire  _T_621; // @[DCache.scala 377:88:freechips.rocketchip.system.DefaultRV32Config.fir@193170.4]
  wire  _T_622; // @[DCache.scala 377:63:freechips.rocketchip.system.DefaultRV32Config.fir@193171.4]
  wire  s2_valid_cached_miss; // @[DCache.scala 377:60:freechips.rocketchip.system.DefaultRV32Config.fir@193172.4]
  wire  s2_want_victimize; // @[DCache.scala 379:79:freechips.rocketchip.system.DefaultRV32Config.fir@193173.4]
  wire  _T_628; // @[DCache.scala 382:49:freechips.rocketchip.system.DefaultRV32Config.fir@193181.4]
  wire  _T_629; // @[DCache.scala 382:92:freechips.rocketchip.system.DefaultRV32Config.fir@193182.4]
  wire  _T_630; // @[DCache.scala 382:67:freechips.rocketchip.system.DefaultRV32Config.fir@193183.4]
  wire  s2_valid_uncached_pending; // @[DCache.scala 382:64:freechips.rocketchip.system.DefaultRV32Config.fir@193184.4]
  reg [19:0] _T_637; // @[Reg.scala 15:16:freechips.rocketchip.system.DefaultRV32Config.fir@193195.4]
  wire [19:0] s2_victim_tag; // @[DCache.scala 384:26:freechips.rocketchip.system.DefaultRV32Config.fir@193199.4]
  reg [1:0] _T_639_state; // @[Reg.scala 15:16:freechips.rocketchip.system.DefaultRV32Config.fir@193201.4]
  wire [1:0] s2_victim_state_state; // @[DCache.scala 385:28:freechips.rocketchip.system.DefaultRV32Config.fir@193205.4]
  wire [2:0] _T_655; // @[Misc.scala 37:36:freechips.rocketchip.system.DefaultRV32Config.fir@193221.4]
  wire [2:0] _T_659; // @[Misc.scala 37:36:freechips.rocketchip.system.DefaultRV32Config.fir@193225.4]
  wire [2:0] _T_663; // @[Misc.scala 37:36:freechips.rocketchip.system.DefaultRV32Config.fir@193229.4]
  wire [2:0] _T_667; // @[Misc.scala 37:36:freechips.rocketchip.system.DefaultRV32Config.fir@193233.4]
  wire [2:0] _T_671; // @[Misc.scala 37:36:freechips.rocketchip.system.DefaultRV32Config.fir@193237.4]
  wire [2:0] _T_675; // @[Misc.scala 37:36:freechips.rocketchip.system.DefaultRV32Config.fir@193241.4]
  wire [1:0] _T_676; // @[Misc.scala 37:63:freechips.rocketchip.system.DefaultRV32Config.fir@193242.4]
  wire [2:0] _T_679; // @[Misc.scala 37:36:freechips.rocketchip.system.DefaultRV32Config.fir@193245.4]
  wire [1:0] _T_680; // @[Misc.scala 37:63:freechips.rocketchip.system.DefaultRV32Config.fir@193246.4]
  wire [2:0] _T_683; // @[Misc.scala 37:36:freechips.rocketchip.system.DefaultRV32Config.fir@193249.4]
  wire [1:0] _T_684; // @[Misc.scala 37:63:freechips.rocketchip.system.DefaultRV32Config.fir@193250.4]
  wire [2:0] _T_687; // @[Misc.scala 37:36:freechips.rocketchip.system.DefaultRV32Config.fir@193253.4]
  wire [1:0] _T_688; // @[Misc.scala 37:63:freechips.rocketchip.system.DefaultRV32Config.fir@193254.4]
  wire [2:0] _T_691; // @[Misc.scala 37:36:freechips.rocketchip.system.DefaultRV32Config.fir@193257.4]
  wire [1:0] _T_692; // @[Misc.scala 37:63:freechips.rocketchip.system.DefaultRV32Config.fir@193258.4]
  wire [2:0] _T_695; // @[Misc.scala 37:36:freechips.rocketchip.system.DefaultRV32Config.fir@193261.4]
  wire [1:0] _T_696; // @[Misc.scala 37:63:freechips.rocketchip.system.DefaultRV32Config.fir@193262.4]
  wire [2:0] s2_report_param; // @[Misc.scala 37:36:freechips.rocketchip.system.DefaultRV32Config.fir@193265.4]
  wire [1:0] probeNewCoh_state; // @[Misc.scala 37:63:freechips.rocketchip.system.DefaultRV32Config.fir@193266.4]
  wire [3:0] _T_705; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@193276.4]
  wire  _T_718; // @[Misc.scala 55:20:freechips.rocketchip.system.DefaultRV32Config.fir@193289.4]
  wire [2:0] _T_720; // @[Misc.scala 37:36:freechips.rocketchip.system.DefaultRV32Config.fir@193291.4]
  wire  _T_722; // @[Misc.scala 55:20:freechips.rocketchip.system.DefaultRV32Config.fir@193293.4]
  wire [2:0] _T_724; // @[Misc.scala 37:36:freechips.rocketchip.system.DefaultRV32Config.fir@193295.4]
  wire  _T_726; // @[Misc.scala 55:20:freechips.rocketchip.system.DefaultRV32Config.fir@193297.4]
  wire [2:0] _T_728; // @[Misc.scala 37:36:freechips.rocketchip.system.DefaultRV32Config.fir@193299.4]
  wire  _T_730; // @[Misc.scala 55:20:freechips.rocketchip.system.DefaultRV32Config.fir@193301.4]
  wire [2:0] _T_732; // @[Misc.scala 37:36:freechips.rocketchip.system.DefaultRV32Config.fir@193303.4]
  wire  _T_734; // @[Misc.scala 55:20:freechips.rocketchip.system.DefaultRV32Config.fir@193305.4]
  wire  _T_735; // @[Misc.scala 37:9:freechips.rocketchip.system.DefaultRV32Config.fir@193306.4]
  wire [2:0] _T_736; // @[Misc.scala 37:36:freechips.rocketchip.system.DefaultRV32Config.fir@193307.4]
  wire  _T_738; // @[Misc.scala 55:20:freechips.rocketchip.system.DefaultRV32Config.fir@193309.4]
  wire  _T_739; // @[Misc.scala 37:9:freechips.rocketchip.system.DefaultRV32Config.fir@193310.4]
  wire [2:0] _T_740; // @[Misc.scala 37:36:freechips.rocketchip.system.DefaultRV32Config.fir@193311.4]
  wire [1:0] _T_741; // @[Misc.scala 37:63:freechips.rocketchip.system.DefaultRV32Config.fir@193312.4]
  wire  _T_742; // @[Misc.scala 55:20:freechips.rocketchip.system.DefaultRV32Config.fir@193313.4]
  wire  _T_743; // @[Misc.scala 37:9:freechips.rocketchip.system.DefaultRV32Config.fir@193314.4]
  wire [2:0] _T_744; // @[Misc.scala 37:36:freechips.rocketchip.system.DefaultRV32Config.fir@193315.4]
  wire [1:0] _T_745; // @[Misc.scala 37:63:freechips.rocketchip.system.DefaultRV32Config.fir@193316.4]
  wire  _T_746; // @[Misc.scala 55:20:freechips.rocketchip.system.DefaultRV32Config.fir@193317.4]
  wire  _T_747; // @[Misc.scala 37:9:freechips.rocketchip.system.DefaultRV32Config.fir@193318.4]
  wire [2:0] _T_748; // @[Misc.scala 37:36:freechips.rocketchip.system.DefaultRV32Config.fir@193319.4]
  wire [1:0] _T_749; // @[Misc.scala 37:63:freechips.rocketchip.system.DefaultRV32Config.fir@193320.4]
  wire  _T_750; // @[Misc.scala 55:20:freechips.rocketchip.system.DefaultRV32Config.fir@193321.4]
  wire  _T_751; // @[Misc.scala 37:9:freechips.rocketchip.system.DefaultRV32Config.fir@193322.4]
  wire [2:0] _T_752; // @[Misc.scala 37:36:freechips.rocketchip.system.DefaultRV32Config.fir@193323.4]
  wire [1:0] _T_753; // @[Misc.scala 37:63:freechips.rocketchip.system.DefaultRV32Config.fir@193324.4]
  wire  _T_754; // @[Misc.scala 55:20:freechips.rocketchip.system.DefaultRV32Config.fir@193325.4]
  wire  _T_755; // @[Misc.scala 37:9:freechips.rocketchip.system.DefaultRV32Config.fir@193326.4]
  wire [2:0] _T_756; // @[Misc.scala 37:36:freechips.rocketchip.system.DefaultRV32Config.fir@193327.4]
  wire [1:0] _T_757; // @[Misc.scala 37:63:freechips.rocketchip.system.DefaultRV32Config.fir@193328.4]
  wire  _T_758; // @[Misc.scala 55:20:freechips.rocketchip.system.DefaultRV32Config.fir@193329.4]
  wire  _T_759; // @[Misc.scala 37:9:freechips.rocketchip.system.DefaultRV32Config.fir@193330.4]
  wire [2:0] _T_760; // @[Misc.scala 37:36:freechips.rocketchip.system.DefaultRV32Config.fir@193331.4]
  wire [1:0] _T_761; // @[Misc.scala 37:63:freechips.rocketchip.system.DefaultRV32Config.fir@193332.4]
  wire  _T_762; // @[Misc.scala 55:20:freechips.rocketchip.system.DefaultRV32Config.fir@193333.4]
  wire  s2_victim_dirty; // @[Misc.scala 37:9:freechips.rocketchip.system.DefaultRV32Config.fir@193334.4]
  wire [2:0] s2_shrink_param; // @[Misc.scala 37:36:freechips.rocketchip.system.DefaultRV32Config.fir@193335.4]
  wire [1:0] voluntaryNewCoh_state; // @[Misc.scala 37:63:freechips.rocketchip.system.DefaultRV32Config.fir@193336.4]
  wire  s2_dont_nack_uncached; // @[DCache.scala 391:57:freechips.rocketchip.system.DefaultRV32Config.fir@193342.4]
  wire  _T_775; // @[DCache.scala 395:17:freechips.rocketchip.system.DefaultRV32Config.fir@193353.4]
  wire  s2_dont_nack_misc; // @[DCache.scala 392:61:freechips.rocketchip.system.DefaultRV32Config.fir@193355.4]
  wire  _T_777; // @[DCache.scala 396:41:freechips.rocketchip.system.DefaultRV32Config.fir@193356.4]
  wire  _T_778; // @[DCache.scala 396:38:freechips.rocketchip.system.DefaultRV32Config.fir@193357.4]
  wire  _T_779; // @[DCache.scala 396:67:freechips.rocketchip.system.DefaultRV32Config.fir@193358.4]
  wire  _T_780; // @[DCache.scala 396:64:freechips.rocketchip.system.DefaultRV32Config.fir@193359.4]
  wire  _T_781; // @[DCache.scala 396:89:freechips.rocketchip.system.DefaultRV32Config.fir@193360.4]
  wire  _T_792; // @[DCache.scala 401:93:freechips.rocketchip.system.DefaultRV32Config.fir@193376.4]
  wire [11:0] _T_808; // @[DCache.scala 405:98:freechips.rocketchip.system.DefaultRV32Config.fir@193396.4]
  wire [1:0] new_meta_coh_state; // @[DCache.scala 408:40:freechips.rocketchip.system.DefaultRV32Config.fir@193402.4]
  wire  _T_823; // @[DCache.scala 425:34:freechips.rocketchip.system.DefaultRV32Config.fir@193434.4]
  wire  _T_824; // @[DCache.scala 425:41:freechips.rocketchip.system.DefaultRV32Config.fir@193435.4]
  wire  lrscBackingOff; // @[DCache.scala 425:38:freechips.rocketchip.system.DefaultRV32Config.fir@193436.4]
  reg [25:0] lrscAddr; // @[DCache.scala 426:21:freechips.rocketchip.system.DefaultRV32Config.fir@193437.4]
  wire  lrscAddrMatch; // @[DCache.scala 427:32:freechips.rocketchip.system.DefaultRV32Config.fir@193439.4]
  wire  _T_826; // @[DCache.scala 428:41:freechips.rocketchip.system.DefaultRV32Config.fir@193440.4]
  wire  _T_827; // @[DCache.scala 428:29:freechips.rocketchip.system.DefaultRV32Config.fir@193441.4]
  wire  s2_sc_fail; // @[DCache.scala 428:26:freechips.rocketchip.system.DefaultRV32Config.fir@193442.4]
  wire  _T_828; // @[DCache.scala 429:23:freechips.rocketchip.system.DefaultRV32Config.fir@193443.4]
  wire  _T_830; // @[DCache.scala 429:32:freechips.rocketchip.system.DefaultRV32Config.fir@193445.4]
  wire  _T_831; // @[DCache.scala 429:54:freechips.rocketchip.system.DefaultRV32Config.fir@193446.4]
  wire [6:0] _T_838; // @[DCache.scala 433:49:freechips.rocketchip.system.DefaultRV32Config.fir@193458.6]
  wire  _T_839; // @[DCache.scala 434:29:freechips.rocketchip.system.DefaultRV32Config.fir@193461.4]
  wire  _T_847; // @[DCache.scala 443:63:freechips.rocketchip.system.DefaultRV32Config.fir@193478.4]
  reg [4:0] pstore1_cmd; // @[Reg.scala 15:16:freechips.rocketchip.system.DefaultRV32Config.fir@193479.4]
  reg [31:0] pstore1_data; // @[Reg.scala 15:16:freechips.rocketchip.system.DefaultRV32Config.fir@193489.4]
  reg [3:0] pstore1_way; // @[Reg.scala 15:16:freechips.rocketchip.system.DefaultRV32Config.fir@193494.4]
  wire  _T_901; // @[DCache.scala 1086:23:freechips.rocketchip.system.DefaultRV32Config.fir@193555.4]
  wire  _T_902; // @[DCache.scala 1085:21:freechips.rocketchip.system.DefaultRV32Config.fir@193556.4]
  reg  pstore1_rmw; // @[Reg.scala 15:16:freechips.rocketchip.system.DefaultRV32Config.fir@193558.4]
  wire  _T_906; // @[DCache.scala 441:46:freechips.rocketchip.system.DefaultRV32Config.fir@193565.4]
  wire  _T_907; // @[DCache.scala 441:61:freechips.rocketchip.system.DefaultRV32Config.fir@193566.4]
  wire  _T_908; // @[DCache.scala 441:58:freechips.rocketchip.system.DefaultRV32Config.fir@193567.4]
  wire  pstore_drain_opportunistic; // @[DCache.scala 453:36:freechips.rocketchip.system.DefaultRV32Config.fir@193639.4]
  reg  _T_976; // @[DCache.scala 454:56:freechips.rocketchip.system.DefaultRV32Config.fir@193643.4]
  wire  pstore_drain_on_miss; // @[DCache.scala 454:46:freechips.rocketchip.system.DefaultRV32Config.fir@193645.4]
  wire  pstore1_valid; // @[DCache.scala 458:38:freechips.rocketchip.system.DefaultRV32Config.fir@193654.4]
  wire  _T_984; // @[DCache.scala 460:54:freechips.rocketchip.system.DefaultRV32Config.fir@193657.4]
  wire  _T_985; // @[DCache.scala 460:85:freechips.rocketchip.system.DefaultRV32Config.fir@193658.4]
  wire  _T_986; // @[DCache.scala 460:98:freechips.rocketchip.system.DefaultRV32Config.fir@193659.4]
  wire  pstore_drain_structural; // @[DCache.scala 460:71:freechips.rocketchip.system.DefaultRV32Config.fir@193660.4]
  wire  _T_990; // @[DCache.scala 457:96:freechips.rocketchip.system.DefaultRV32Config.fir@193664.4]
  wire  _T_991; // @[DCache.scala 461:63:freechips.rocketchip.system.DefaultRV32Config.fir@193665.4]
  wire  _T_992; // @[DCache.scala 461:22:freechips.rocketchip.system.DefaultRV32Config.fir@193666.4]
  wire  _T_994; // @[DCache.scala 461:9:freechips.rocketchip.system.DefaultRV32Config.fir@193668.4]
  wire  _T_995; // @[DCache.scala 461:9:freechips.rocketchip.system.DefaultRV32Config.fir@193669.4]
  wire  _T_1004; // @[DCache.scala 469:44:freechips.rocketchip.system.DefaultRV32Config.fir@193683.4]
  wire  _T_1005; // @[DCache.scala 469:41:freechips.rocketchip.system.DefaultRV32Config.fir@193684.4]
  wire  _T_1006; // @[DCache.scala 469:58:freechips.rocketchip.system.DefaultRV32Config.fir@193685.4]
  wire  _T_1007; // @[DCache.scala 469:107:freechips.rocketchip.system.DefaultRV32Config.fir@193686.4]
  wire  _T_1008; // @[DCache.scala 469:76:freechips.rocketchip.system.DefaultRV32Config.fir@193687.4]
  wire  pstore_drain; // @[DCache.scala 468:48:freechips.rocketchip.system.DefaultRV32Config.fir@193688.4]
  wire  _T_1018; // @[DCache.scala 472:71:freechips.rocketchip.system.DefaultRV32Config.fir@193698.4]
  wire  _T_1019; // @[DCache.scala 472:91:freechips.rocketchip.system.DefaultRV32Config.fir@193699.4]
  wire  _T_1022; // @[DCache.scala 473:79:freechips.rocketchip.system.DefaultRV32Config.fir@193703.4]
  wire  advance_pstore1; // @[DCache.scala 473:61:freechips.rocketchip.system.DefaultRV32Config.fir@193704.4]
  wire  _T_1024; // @[DCache.scala 474:34:freechips.rocketchip.system.DefaultRV32Config.fir@193706.4]
  reg [3:0] pstore2_way; // @[Reg.scala 15:16:freechips.rocketchip.system.DefaultRV32Config.fir@193715.4]
  wire [31:0] pstore1_storegen_data; // @[:freechips.rocketchip.system.DefaultRV32Config.fir@193503.4 :freechips.rocketchip.system.DefaultRV32Config.fir@193505.4 DCache.scala 888:27:freechips.rocketchip.system.DefaultRV32Config.fir@195717.4]
  reg [7:0] _T_1032; // @[Reg.scala 15:16:freechips.rocketchip.system.DefaultRV32Config.fir@193723.4]
  reg [7:0] _T_1037; // @[Reg.scala 15:16:freechips.rocketchip.system.DefaultRV32Config.fir@193731.4]
  reg [7:0] _T_1042; // @[Reg.scala 15:16:freechips.rocketchip.system.DefaultRV32Config.fir@193739.4]
  reg [7:0] _T_1047; // @[Reg.scala 15:16:freechips.rocketchip.system.DefaultRV32Config.fir@193747.4]
  wire [31:0] pstore2_storegen_data; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@193753.4]
  wire [3:0] _T_1052; // @[DCache.scala 485:37:freechips.rocketchip.system.DefaultRV32Config.fir@193759.6]
  wire [3:0] _T_1054; // @[DCache.scala 485:15:freechips.rocketchip.system.DefaultRV32Config.fir@193761.6]
  wire [31:0] _T_1068; // @[DCache.scala 500:36:freechips.rocketchip.system.DefaultRV32Config.fir@193781.4]
  wire [31:0] _T_1070; // @[DCache.scala 502:63:freechips.rocketchip.system.DefaultRV32Config.fir@193785.4]
  wire [15:0] _T_1075; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@193790.4]
  wire [15:0] _T_1076; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@193791.4]
  wire [3:0] _T_1080; // @[DCache.scala 504:47:freechips.rocketchip.system.DefaultRV32Config.fir@193797.4]
  wire  _T_1085; // @[DCache.scala 1076:66:freechips.rocketchip.system.DefaultRV32Config.fir@193802.4]
  wire  _T_1086; // @[DCache.scala 1076:66:freechips.rocketchip.system.DefaultRV32Config.fir@193803.4]
  wire  _T_1087; // @[DCache.scala 1076:66:freechips.rocketchip.system.DefaultRV32Config.fir@193804.4]
  wire  _T_1088; // @[DCache.scala 1076:66:freechips.rocketchip.system.DefaultRV32Config.fir@193805.4]
  wire [1:0] _T_1089; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@193806.4]
  wire [1:0] _T_1090; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@193807.4]
  wire  _T_1190; // @[DCache.scala 524:34:freechips.rocketchip.system.DefaultRV32Config.fir@193916.4]
  wire [1:0] _T_1191; // @[DCache.scala 524:59:freechips.rocketchip.system.DefaultRV32Config.fir@193917.4]
  wire  a_source; // @[Mux.scala 47:69:freechips.rocketchip.system.DefaultRV32Config.fir@193920.4]
  wire [31:0] acquire_address; // @[DCache.scala 525:49:freechips.rocketchip.system.DefaultRV32Config.fir@193922.4]
  wire [18:0] a_mask; // @[DCache.scala 529:29:freechips.rocketchip.system.DefaultRV32Config.fir@193924.4]
  wire [1:0] _T_1250; // @[OneHot.scala 65:12:freechips.rocketchip.system.DefaultRV32Config.fir@193986.4]
  wire [1:0] _T_1252; // @[Misc.scala 201:81:freechips.rocketchip.system.DefaultRV32Config.fir@193988.4]
  wire  _T_1253; // @[Misc.scala 205:21:freechips.rocketchip.system.DefaultRV32Config.fir@193989.4]
  wire  _T_1256; // @[Misc.scala 210:20:freechips.rocketchip.system.DefaultRV32Config.fir@193992.4]
  wire  _T_1258; // @[Misc.scala 214:38:freechips.rocketchip.system.DefaultRV32Config.fir@193994.4]
  wire  _T_1259; // @[Misc.scala 214:29:freechips.rocketchip.system.DefaultRV32Config.fir@193995.4]
  wire  _T_1261; // @[Misc.scala 214:38:freechips.rocketchip.system.DefaultRV32Config.fir@193997.4]
  wire  _T_1262; // @[Misc.scala 214:29:freechips.rocketchip.system.DefaultRV32Config.fir@193998.4]
  wire  _T_1265; // @[Misc.scala 210:20:freechips.rocketchip.system.DefaultRV32Config.fir@194001.4]
  wire  _T_1266; // @[Misc.scala 213:27:freechips.rocketchip.system.DefaultRV32Config.fir@194002.4]
  wire  _T_1267; // @[Misc.scala 214:38:freechips.rocketchip.system.DefaultRV32Config.fir@194003.4]
  wire  _T_1268; // @[Misc.scala 214:29:freechips.rocketchip.system.DefaultRV32Config.fir@194004.4]
  wire  _T_1269; // @[Misc.scala 213:27:freechips.rocketchip.system.DefaultRV32Config.fir@194005.4]
  wire  _T_1270; // @[Misc.scala 214:38:freechips.rocketchip.system.DefaultRV32Config.fir@194006.4]
  wire  _T_1271; // @[Misc.scala 214:29:freechips.rocketchip.system.DefaultRV32Config.fir@194007.4]
  wire  _T_1272; // @[Misc.scala 213:27:freechips.rocketchip.system.DefaultRV32Config.fir@194008.4]
  wire  _T_1273; // @[Misc.scala 214:38:freechips.rocketchip.system.DefaultRV32Config.fir@194009.4]
  wire  _T_1274; // @[Misc.scala 214:29:freechips.rocketchip.system.DefaultRV32Config.fir@194010.4]
  wire  _T_1275; // @[Misc.scala 213:27:freechips.rocketchip.system.DefaultRV32Config.fir@194011.4]
  wire  _T_1276; // @[Misc.scala 214:38:freechips.rocketchip.system.DefaultRV32Config.fir@194012.4]
  wire  _T_1277; // @[Misc.scala 214:29:freechips.rocketchip.system.DefaultRV32Config.fir@194013.4]
  wire [3:0] get_mask; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@194016.4]
  wire  _T_2072; // @[Mux.scala 80:60:freechips.rocketchip.system.DefaultRV32Config.fir@194913.4]
  wire [2:0] _T_2073_opcode; // @[Mux.scala 80:57:freechips.rocketchip.system.DefaultRV32Config.fir@194914.4]
  wire [3:0] _T_1470_size; // @[Edges.scala 515:17:freechips.rocketchip.system.DefaultRV32Config.fir@194230.4 Edges.scala 518:15:freechips.rocketchip.system.DefaultRV32Config.fir@194234.4]
  wire [3:0] _T_2073_size; // @[Mux.scala 80:57:freechips.rocketchip.system.DefaultRV32Config.fir@194914.4]
  wire  _T_2073_source; // @[Mux.scala 80:57:freechips.rocketchip.system.DefaultRV32Config.fir@194914.4]
  wire [31:0] _T_2073_address; // @[Mux.scala 80:57:freechips.rocketchip.system.DefaultRV32Config.fir@194914.4]
  wire [3:0] _T_2073_mask; // @[Mux.scala 80:57:freechips.rocketchip.system.DefaultRV32Config.fir@194914.4]
  wire [31:0] _T_2073_data; // @[Mux.scala 80:57:freechips.rocketchip.system.DefaultRV32Config.fir@194914.4]
  wire  _T_2074; // @[Mux.scala 80:60:freechips.rocketchip.system.DefaultRV32Config.fir@194915.4]
  wire [2:0] _T_2075_opcode; // @[Mux.scala 80:57:freechips.rocketchip.system.DefaultRV32Config.fir@194916.4]
  wire [2:0] _T_2075_param; // @[Mux.scala 80:57:freechips.rocketchip.system.DefaultRV32Config.fir@194916.4]
  wire [3:0] _T_2075_size; // @[Mux.scala 80:57:freechips.rocketchip.system.DefaultRV32Config.fir@194916.4]
  wire  _T_2075_source; // @[Mux.scala 80:57:freechips.rocketchip.system.DefaultRV32Config.fir@194916.4]
  wire [31:0] _T_2075_address; // @[Mux.scala 80:57:freechips.rocketchip.system.DefaultRV32Config.fir@194916.4]
  wire [3:0] _T_2075_mask; // @[Mux.scala 80:57:freechips.rocketchip.system.DefaultRV32Config.fir@194916.4]
  wire [31:0] _T_2075_data; // @[Mux.scala 80:57:freechips.rocketchip.system.DefaultRV32Config.fir@194916.4]
  wire  _T_2076; // @[Mux.scala 80:60:freechips.rocketchip.system.DefaultRV32Config.fir@194917.4]
  wire [2:0] _T_2077_opcode; // @[Mux.scala 80:57:freechips.rocketchip.system.DefaultRV32Config.fir@194918.4]
  wire [2:0] _T_2077_param; // @[Mux.scala 80:57:freechips.rocketchip.system.DefaultRV32Config.fir@194918.4]
  wire [3:0] _T_2077_size; // @[Mux.scala 80:57:freechips.rocketchip.system.DefaultRV32Config.fir@194918.4]
  wire  _T_2077_source; // @[Mux.scala 80:57:freechips.rocketchip.system.DefaultRV32Config.fir@194918.4]
  wire [31:0] _T_2077_address; // @[Mux.scala 80:57:freechips.rocketchip.system.DefaultRV32Config.fir@194918.4]
  wire [3:0] _T_2077_mask; // @[Mux.scala 80:57:freechips.rocketchip.system.DefaultRV32Config.fir@194918.4]
  wire [31:0] _T_2077_data; // @[Mux.scala 80:57:freechips.rocketchip.system.DefaultRV32Config.fir@194918.4]
  wire  _T_2078; // @[Mux.scala 80:60:freechips.rocketchip.system.DefaultRV32Config.fir@194919.4]
  wire [2:0] _T_2079_opcode; // @[Mux.scala 80:57:freechips.rocketchip.system.DefaultRV32Config.fir@194920.4]
  wire [2:0] _T_2079_param; // @[Mux.scala 80:57:freechips.rocketchip.system.DefaultRV32Config.fir@194920.4]
  wire [3:0] _T_2079_size; // @[Mux.scala 80:57:freechips.rocketchip.system.DefaultRV32Config.fir@194920.4]
  wire  _T_2079_source; // @[Mux.scala 80:57:freechips.rocketchip.system.DefaultRV32Config.fir@194920.4]
  wire [31:0] _T_2079_address; // @[Mux.scala 80:57:freechips.rocketchip.system.DefaultRV32Config.fir@194920.4]
  wire [3:0] _T_2079_mask; // @[Mux.scala 80:57:freechips.rocketchip.system.DefaultRV32Config.fir@194920.4]
  wire [31:0] _T_2079_data; // @[Mux.scala 80:57:freechips.rocketchip.system.DefaultRV32Config.fir@194920.4]
  wire  _T_2080; // @[Mux.scala 80:60:freechips.rocketchip.system.DefaultRV32Config.fir@194921.4]
  wire [2:0] _T_2081_opcode; // @[Mux.scala 80:57:freechips.rocketchip.system.DefaultRV32Config.fir@194922.4]
  wire [2:0] _T_2081_param; // @[Mux.scala 80:57:freechips.rocketchip.system.DefaultRV32Config.fir@194922.4]
  wire [3:0] _T_2081_size; // @[Mux.scala 80:57:freechips.rocketchip.system.DefaultRV32Config.fir@194922.4]
  wire  _T_2081_source; // @[Mux.scala 80:57:freechips.rocketchip.system.DefaultRV32Config.fir@194922.4]
  wire [31:0] _T_2081_address; // @[Mux.scala 80:57:freechips.rocketchip.system.DefaultRV32Config.fir@194922.4]
  wire [3:0] _T_2081_mask; // @[Mux.scala 80:57:freechips.rocketchip.system.DefaultRV32Config.fir@194922.4]
  wire [31:0] _T_2081_data; // @[Mux.scala 80:57:freechips.rocketchip.system.DefaultRV32Config.fir@194922.4]
  wire  _T_2082; // @[Mux.scala 80:60:freechips.rocketchip.system.DefaultRV32Config.fir@194923.4]
  wire [2:0] _T_2083_opcode; // @[Mux.scala 80:57:freechips.rocketchip.system.DefaultRV32Config.fir@194924.4]
  wire [2:0] _T_2083_param; // @[Mux.scala 80:57:freechips.rocketchip.system.DefaultRV32Config.fir@194924.4]
  wire [3:0] _T_2083_size; // @[Mux.scala 80:57:freechips.rocketchip.system.DefaultRV32Config.fir@194924.4]
  wire  _T_2083_source; // @[Mux.scala 80:57:freechips.rocketchip.system.DefaultRV32Config.fir@194924.4]
  wire [31:0] _T_2083_address; // @[Mux.scala 80:57:freechips.rocketchip.system.DefaultRV32Config.fir@194924.4]
  wire [3:0] _T_2083_mask; // @[Mux.scala 80:57:freechips.rocketchip.system.DefaultRV32Config.fir@194924.4]
  wire [31:0] _T_2083_data; // @[Mux.scala 80:57:freechips.rocketchip.system.DefaultRV32Config.fir@194924.4]
  wire  _T_2084; // @[Mux.scala 80:60:freechips.rocketchip.system.DefaultRV32Config.fir@194925.4]
  wire [2:0] _T_2085_opcode; // @[Mux.scala 80:57:freechips.rocketchip.system.DefaultRV32Config.fir@194926.4]
  wire [2:0] _T_2085_param; // @[Mux.scala 80:57:freechips.rocketchip.system.DefaultRV32Config.fir@194926.4]
  wire [3:0] _T_2085_size; // @[Mux.scala 80:57:freechips.rocketchip.system.DefaultRV32Config.fir@194926.4]
  wire  _T_2085_source; // @[Mux.scala 80:57:freechips.rocketchip.system.DefaultRV32Config.fir@194926.4]
  wire [31:0] _T_2085_address; // @[Mux.scala 80:57:freechips.rocketchip.system.DefaultRV32Config.fir@194926.4]
  wire [3:0] _T_2085_mask; // @[Mux.scala 80:57:freechips.rocketchip.system.DefaultRV32Config.fir@194926.4]
  wire [31:0] _T_2085_data; // @[Mux.scala 80:57:freechips.rocketchip.system.DefaultRV32Config.fir@194926.4]
  wire  _T_2086; // @[Mux.scala 80:60:freechips.rocketchip.system.DefaultRV32Config.fir@194927.4]
  wire [2:0] _T_2087_opcode; // @[Mux.scala 80:57:freechips.rocketchip.system.DefaultRV32Config.fir@194928.4]
  wire [2:0] _T_2087_param; // @[Mux.scala 80:57:freechips.rocketchip.system.DefaultRV32Config.fir@194928.4]
  wire [3:0] _T_2087_size; // @[Mux.scala 80:57:freechips.rocketchip.system.DefaultRV32Config.fir@194928.4]
  wire  _T_2087_source; // @[Mux.scala 80:57:freechips.rocketchip.system.DefaultRV32Config.fir@194928.4]
  wire [31:0] _T_2087_address; // @[Mux.scala 80:57:freechips.rocketchip.system.DefaultRV32Config.fir@194928.4]
  wire [3:0] _T_2087_mask; // @[Mux.scala 80:57:freechips.rocketchip.system.DefaultRV32Config.fir@194928.4]
  wire [31:0] _T_2087_data; // @[Mux.scala 80:57:freechips.rocketchip.system.DefaultRV32Config.fir@194928.4]
  wire  _T_2088; // @[Mux.scala 80:60:freechips.rocketchip.system.DefaultRV32Config.fir@194929.4]
  wire [2:0] atomics_opcode; // @[Mux.scala 80:57:freechips.rocketchip.system.DefaultRV32Config.fir@194930.4]
  wire [2:0] atomics_param; // @[Mux.scala 80:57:freechips.rocketchip.system.DefaultRV32Config.fir@194930.4]
  wire [3:0] atomics_size; // @[Mux.scala 80:57:freechips.rocketchip.system.DefaultRV32Config.fir@194930.4]
  wire  atomics_source; // @[Mux.scala 80:57:freechips.rocketchip.system.DefaultRV32Config.fir@194930.4]
  wire [31:0] atomics_address; // @[Mux.scala 80:57:freechips.rocketchip.system.DefaultRV32Config.fir@194930.4]
  wire [3:0] atomics_mask; // @[Mux.scala 80:57:freechips.rocketchip.system.DefaultRV32Config.fir@194930.4]
  wire [31:0] atomics_data; // @[Mux.scala 80:57:freechips.rocketchip.system.DefaultRV32Config.fir@194930.4]
  wire  _T_2090; // @[DCache.scala 551:30:freechips.rocketchip.system.DefaultRV32Config.fir@194932.4]
  wire  _T_2091; // @[DCache.scala 551:27:freechips.rocketchip.system.DefaultRV32Config.fir@194933.4]
  wire  _T_2093; // @[DCache.scala 551:117:freechips.rocketchip.system.DefaultRV32Config.fir@194935.4]
  wire  _T_2095; // @[DCache.scala 551:48:freechips.rocketchip.system.DefaultRV32Config.fir@194937.4]
  wire  tl_out_a_valid; // @[DCache.scala 550:67:freechips.rocketchip.system.DefaultRV32Config.fir@194938.4]
  wire  _T_2154; // @[DCache.scala 553:9:freechips.rocketchip.system.DefaultRV32Config.fir@195006.4]
  wire  _T_2156; // @[DCache.scala 555:9:freechips.rocketchip.system.DefaultRV32Config.fir@195008.4]
  wire [2:0] _T_2157_opcode; // @[DCache.scala 555:8:freechips.rocketchip.system.DefaultRV32Config.fir@195009.4]
  wire [2:0] _T_2157_param; // @[DCache.scala 555:8:freechips.rocketchip.system.DefaultRV32Config.fir@195009.4]
  wire [3:0] _T_2157_size; // @[DCache.scala 555:8:freechips.rocketchip.system.DefaultRV32Config.fir@195009.4]
  wire  _T_2157_source; // @[DCache.scala 555:8:freechips.rocketchip.system.DefaultRV32Config.fir@195009.4]
  wire [31:0] _T_2157_address; // @[DCache.scala 555:8:freechips.rocketchip.system.DefaultRV32Config.fir@195009.4]
  wire [3:0] _T_2157_mask; // @[DCache.scala 555:8:freechips.rocketchip.system.DefaultRV32Config.fir@195009.4]
  wire [31:0] _T_2157_data; // @[DCache.scala 555:8:freechips.rocketchip.system.DefaultRV32Config.fir@195009.4]
  wire [2:0] _T_2158_opcode; // @[DCache.scala 554:8:freechips.rocketchip.system.DefaultRV32Config.fir@195010.4]
  wire [2:0] _T_2158_param; // @[DCache.scala 554:8:freechips.rocketchip.system.DefaultRV32Config.fir@195010.4]
  wire [3:0] _T_2158_size; // @[DCache.scala 554:8:freechips.rocketchip.system.DefaultRV32Config.fir@195010.4]
  wire  _T_2158_source; // @[DCache.scala 554:8:freechips.rocketchip.system.DefaultRV32Config.fir@195010.4]
  wire [31:0] _T_2158_address; // @[DCache.scala 554:8:freechips.rocketchip.system.DefaultRV32Config.fir@195010.4]
  wire [3:0] putpartial_mask; // @[Edges.scala 485:17:freechips.rocketchip.system.DefaultRV32Config.fir@194181.4 Edges.scala 491:15:freechips.rocketchip.system.DefaultRV32Config.fir@194188.4]
  wire [3:0] _T_2158_mask; // @[DCache.scala 554:8:freechips.rocketchip.system.DefaultRV32Config.fir@195010.4]
  wire [31:0] _T_2158_data; // @[DCache.scala 554:8:freechips.rocketchip.system.DefaultRV32Config.fir@195010.4]
  wire [2:0] _T_2159_opcode; // @[DCache.scala 553:8:freechips.rocketchip.system.DefaultRV32Config.fir@195011.4]
  wire [2:0] _T_2159_param; // @[DCache.scala 553:8:freechips.rocketchip.system.DefaultRV32Config.fir@195011.4]
  wire [3:0] _T_2159_size; // @[DCache.scala 553:8:freechips.rocketchip.system.DefaultRV32Config.fir@195011.4]
  wire  _T_2159_source; // @[DCache.scala 553:8:freechips.rocketchip.system.DefaultRV32Config.fir@195011.4]
  wire [31:0] _T_2159_address; // @[DCache.scala 553:8:freechips.rocketchip.system.DefaultRV32Config.fir@195011.4]
  wire [3:0] _T_2159_mask; // @[DCache.scala 553:8:freechips.rocketchip.system.DefaultRV32Config.fir@195011.4]
  wire [31:0] _T_2159_data; // @[DCache.scala 553:8:freechips.rocketchip.system.DefaultRV32Config.fir@195011.4]
  wire [2:0] _T_2120_param; // @[Edges.scala 347:17:freechips.rocketchip.system.DefaultRV32Config.fir@194963.4 Edges.scala 349:15:freechips.rocketchip.system.DefaultRV32Config.fir@194966.4]
  wire [1:0] _T_2162; // @[OneHot.scala 65:12:freechips.rocketchip.system.DefaultRV32Config.fir@195015.4]
  wire  a_sel; // @[DCache.scala 574:66:freechips.rocketchip.system.DefaultRV32Config.fir@195017.4]
  wire  _T_2164; // @[Decoupled.scala 40:37:freechips.rocketchip.system.DefaultRV32Config.fir@195018.4]
  wire  _GEN_139; // @[DCache.scala 578:18:freechips.rocketchip.system.DefaultRV32Config.fir@195022.8]
  wire [26:0] _T_2171; // @[package.scala 207:77:freechips.rocketchip.system.DefaultRV32Config.fir@195037.4]
  wire [11:0] _T_2173; // @[package.scala 207:46:freechips.rocketchip.system.DefaultRV32Config.fir@195039.4]
  wire [9:0] _T_2176; // @[Edges.scala 222:14:freechips.rocketchip.system.DefaultRV32Config.fir@195042.4]
  wire [9:0] _T_2179; // @[Edges.scala 231:28:freechips.rocketchip.system.DefaultRV32Config.fir@195045.4]
  wire  _T_2180; // @[Edges.scala 233:25:freechips.rocketchip.system.DefaultRV32Config.fir@195047.4]
  wire  _T_2181; // @[Edges.scala 233:47:freechips.rocketchip.system.DefaultRV32Config.fir@195048.4]
  wire  d_last; // @[Edges.scala 233:37:freechips.rocketchip.system.DefaultRV32Config.fir@195049.4]
  wire  d_done; // @[Edges.scala 234:22:freechips.rocketchip.system.DefaultRV32Config.fir@195050.4]
  wire [9:0] _T_2182; // @[Edges.scala 235:27:freechips.rocketchip.system.DefaultRV32Config.fir@195051.4]
  wire [9:0] _T_2183; // @[Edges.scala 235:25:freechips.rocketchip.system.DefaultRV32Config.fir@195052.4]
  wire [11:0] d_address_inc; // @[Edges.scala 270:29:freechips.rocketchip.system.DefaultRV32Config.fir@195057.4]
  wire  _T_2192; // @[DCache.scala 606:129:freechips.rocketchip.system.DefaultRV32Config.fir@195067.4]
  wire  grantIsVoluntary; // @[DCache.scala 608:32:freechips.rocketchip.system.DefaultRV32Config.fir@195080.4]
  wire [2:0] _T_2205; // @[DCache.scala 612:97:freechips.rocketchip.system.DefaultRV32Config.fir@195087.6]
  wire [1:0] _T_2214; // @[OneHot.scala 65:12:freechips.rocketchip.system.DefaultRV32Config.fir@195100.4]
  wire  uncachedRespIdxOH; // @[DCache.scala 615:90:freechips.rocketchip.system.DefaultRV32Config.fir@195102.4]
  wire  _T_2219; // @[DCache.scala 620:13:freechips.rocketchip.system.DefaultRV32Config.fir@195110.8]
  wire  _T_2220; // @[DCache.scala 620:13:freechips.rocketchip.system.DefaultRV32Config.fir@195111.8]
  wire  _T_2222; // @[DCache.scala 629:17:freechips.rocketchip.system.DefaultRV32Config.fir@195126.10]
  wire  _T_2224; // @[DCache.scala 630:17:freechips.rocketchip.system.DefaultRV32Config.fir@195129.12]
  wire  _T_2225; // @[DCache.scala 630:17:freechips.rocketchip.system.DefaultRV32Config.fir@195130.12]
  wire [31:0] dontCareBits; // @[DCache.scala 644:55:freechips.rocketchip.system.DefaultRV32Config.fir@195145.12]
  wire [31:0] _GEN_376; // @[DCache.scala 645:26:freechips.rocketchip.system.DefaultRV32Config.fir@195147.12]
  wire [31:0] _T_2229; // @[DCache.scala 645:26:freechips.rocketchip.system.DefaultRV32Config.fir@195147.12]
  wire  _T_2231; // @[DCache.scala 651:13:freechips.rocketchip.system.DefaultRV32Config.fir@195155.12]
  wire  _T_2232; // @[DCache.scala 651:13:freechips.rocketchip.system.DefaultRV32Config.fir@195156.12]
  wire  _GEN_191; // @[DCache.scala 650:36:freechips.rocketchip.system.DefaultRV32Config.fir@195153.10]
  wire  _GEN_200; // @[DCache.scala 627:35:freechips.rocketchip.system.DefaultRV32Config.fir@195124.8]
  wire  _GEN_204; // @[DCache.scala 618:26:freechips.rocketchip.system.DefaultRV32Config.fir@195107.6]
  wire  _GEN_213; // @[DCache.scala 618:26:freechips.rocketchip.system.DefaultRV32Config.fir@195107.6]
  wire  _GEN_226; // @[DCache.scala 617:26:freechips.rocketchip.system.DefaultRV32Config.fir@195106.4]
  wire  _T_2233; // @[DCache.scala 657:36:freechips.rocketchip.system.DefaultRV32Config.fir@195164.4]
  wire  _T_2234; // @[DCache.scala 657:47:freechips.rocketchip.system.DefaultRV32Config.fir@195165.4]
  wire  _T_2235; // @[DCache.scala 657:64:freechips.rocketchip.system.DefaultRV32Config.fir@195166.4]
  wire  tl_out__e_valid; // @[DCache.scala 665:51:freechips.rocketchip.system.DefaultRV32Config.fir@195189.4]
  wire  _T_2237; // @[Decoupled.scala 40:37:freechips.rocketchip.system.DefaultRV32Config.fir@195172.4]
  wire  _T_2239; // @[DCache.scala 659:47:freechips.rocketchip.system.DefaultRV32Config.fir@195174.4]
  wire  _T_2240; // @[DCache.scala 659:58:freechips.rocketchip.system.DefaultRV32Config.fir@195175.4]
  wire  _T_2241; // @[DCache.scala 659:26:freechips.rocketchip.system.DefaultRV32Config.fir@195176.4]
  wire  _T_2243; // @[DCache.scala 659:9:freechips.rocketchip.system.DefaultRV32Config.fir@195178.4]
  wire  _T_2244; // @[DCache.scala 659:9:freechips.rocketchip.system.DefaultRV32Config.fir@195179.4]
  wire  _T_2245; // @[DCache.scala 664:44:freechips.rocketchip.system.DefaultRV32Config.fir@195184.4]
  wire  _T_2246; // @[DCache.scala 664:61:freechips.rocketchip.system.DefaultRV32Config.fir@195185.4]
  wire [31:0] _T_2250; // @[DCache.scala 671:57:freechips.rocketchip.system.DefaultRV32Config.fir@195195.4]
  wire [31:0] _GEN_377; // @[DCache.scala 671:67:freechips.rocketchip.system.DefaultRV32Config.fir@195196.4]
  wire [31:0] _T_2251; // @[DCache.scala 671:67:freechips.rocketchip.system.DefaultRV32Config.fir@195196.4]
  wire  _T_2254; // @[DCache.scala 684:43:freechips.rocketchip.system.DefaultRV32Config.fir@195204.4]
  wire  _T_2255; // @[DCache.scala 684:56:freechips.rocketchip.system.DefaultRV32Config.fir@195205.4]
  wire [3:0] _T_2313; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@195268.4]
  wire  _T_2322; // @[Mux.scala 80:60:freechips.rocketchip.system.DefaultRV32Config.fir@195277.4]
  wire [1:0] _T_2323; // @[Mux.scala 80:57:freechips.rocketchip.system.DefaultRV32Config.fir@195278.4]
  wire  _T_2324; // @[Mux.scala 80:60:freechips.rocketchip.system.DefaultRV32Config.fir@195279.4]
  wire [1:0] _T_2325; // @[Mux.scala 80:57:freechips.rocketchip.system.DefaultRV32Config.fir@195280.4]
  wire  _T_2326; // @[Mux.scala 80:60:freechips.rocketchip.system.DefaultRV32Config.fir@195281.4]
  wire [1:0] _T_2327; // @[Mux.scala 80:57:freechips.rocketchip.system.DefaultRV32Config.fir@195282.4]
  wire  _T_2328; // @[Mux.scala 80:60:freechips.rocketchip.system.DefaultRV32Config.fir@195283.4]
  wire [1:0] _T_2329; // @[Mux.scala 80:57:freechips.rocketchip.system.DefaultRV32Config.fir@195284.4]
  wire  _GEN_229; // @[DCache.scala 698:29:freechips.rocketchip.system.DefaultRV32Config.fir@195300.6]
  wire  _GEN_230; // @[DCache.scala 698:29:freechips.rocketchip.system.DefaultRV32Config.fir@195300.6]
  wire  _GEN_231; // @[DCache.scala 698:29:freechips.rocketchip.system.DefaultRV32Config.fir@195300.6]
  wire  _T_2343; // @[DCache.scala 712:48:freechips.rocketchip.system.DefaultRV32Config.fir@195318.4]
  wire  _T_2344; // @[DCache.scala 712:79:freechips.rocketchip.system.DefaultRV32Config.fir@195319.4]
  wire  _T_2345; // @[DCache.scala 712:44:freechips.rocketchip.system.DefaultRV32Config.fir@195320.4]
  wire [32:0] _T_2353; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@195332.4]
  wire [9:0] _T_2364; // @[Edges.scala 231:28:freechips.rocketchip.system.DefaultRV32Config.fir@195346.4]
  wire [9:0] _T_2367; // @[Edges.scala 235:27:freechips.rocketchip.system.DefaultRV32Config.fir@195352.4]
  wire [9:0] c_count; // @[Edges.scala 235:25:freechips.rocketchip.system.DefaultRV32Config.fir@195353.4]
  reg  s1_release_data_valid; // @[DCache.scala 723:34:freechips.rocketchip.system.DefaultRV32Config.fir@195361.4]
  wire  _T_2373; // @[DCache.scala 725:47:freechips.rocketchip.system.DefaultRV32Config.fir@195368.4]
  wire  releaseRejected; // @[DCache.scala 725:44:freechips.rocketchip.system.DefaultRV32Config.fir@195369.4]
  wire  _T_2370; // @[DCache.scala 724:67:freechips.rocketchip.system.DefaultRV32Config.fir@195363.4]
  wire [10:0] _T_2375; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@195371.4]
  wire [1:0] _T_2376; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@195372.4]
  wire [1:0] _GEN_378; // @[DCache.scala 726:101:freechips.rocketchip.system.DefaultRV32Config.fir@195373.4]
  wire [1:0] _T_2378; // @[DCache.scala 726:101:freechips.rocketchip.system.DefaultRV32Config.fir@195374.4]
  wire [1:0] _T_2379; // @[DCache.scala 726:52:freechips.rocketchip.system.DefaultRV32Config.fir@195375.4]
  wire [10:0] _GEN_379; // @[DCache.scala 726:47:freechips.rocketchip.system.DefaultRV32Config.fir@195376.4]
  wire [10:0] releaseDataBeat; // @[DCache.scala 726:47:freechips.rocketchip.system.DefaultRV32Config.fir@195377.4]
  wire  _T_2385; // @[DCache.scala 739:52:freechips.rocketchip.system.DefaultRV32Config.fir@195416.6]
  wire  _T_2387; // @[DCache.scala 739:13:freechips.rocketchip.system.DefaultRV32Config.fir@195418.6]
  wire  _T_2388; // @[DCache.scala 739:13:freechips.rocketchip.system.DefaultRV32Config.fir@195419.6]
  wire  discard_line; // @[DCache.scala 740:46:freechips.rocketchip.system.DefaultRV32Config.fir@195425.6]
  wire  _T_2393; // @[DCache.scala 741:47:freechips.rocketchip.system.DefaultRV32Config.fir@195429.6]
  wire  _T_2394; // @[DCache.scala 741:44:freechips.rocketchip.system.DefaultRV32Config.fir@195430.6]
  wire [2:0] _T_2395; // @[DCache.scala 741:27:freechips.rocketchip.system.DefaultRV32Config.fir@195431.6]
  wire [25:0] _T_2397; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@195434.6]
  wire [31:0] res_2_address; // @[DCache.scala 742:96:freechips.rocketchip.system.DefaultRV32Config.fir@195435.6]
  wire [2:0] _GEN_239; // @[DCache.scala 738:25:freechips.rocketchip.system.DefaultRV32Config.fir@195414.4]
  wire [2:0] _T_2400; // @[DCache.scala 753:29:freechips.rocketchip.system.DefaultRV32Config.fir@195458.12]
  wire [2:0] _T_2402; // @[DCache.scala 757:29:freechips.rocketchip.system.DefaultRV32Config.fir@195465.12]
  wire [2:0] _GEN_250; // @[DCache.scala 750:45:freechips.rocketchip.system.DefaultRV32Config.fir@195455.10]
  wire [2:0] _GEN_256; // @[DCache.scala 750:45:freechips.rocketchip.system.DefaultRV32Config.fir@195455.10]
  wire [2:0] _GEN_258; // @[DCache.scala 748:36:freechips.rocketchip.system.DefaultRV32Config.fir@195450.8]
  wire [2:0] _GEN_261; // @[DCache.scala 748:36:freechips.rocketchip.system.DefaultRV32Config.fir@195450.8]
  wire [2:0] _GEN_268; // @[DCache.scala 746:28:freechips.rocketchip.system.DefaultRV32Config.fir@195446.6]
  wire [2:0] _GEN_271; // @[DCache.scala 746:28:freechips.rocketchip.system.DefaultRV32Config.fir@195446.6]
  wire [2:0] _GEN_279; // @[DCache.scala 744:21:freechips.rocketchip.system.DefaultRV32Config.fir@195442.4]
  wire [2:0] _GEN_282; // @[DCache.scala 744:21:freechips.rocketchip.system.DefaultRV32Config.fir@195442.4]
  wire  _T_2403; // @[DCache.scala 761:25:freechips.rocketchip.system.DefaultRV32Config.fir@195472.4]
  wire [32:0] _T_2406; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@195478.6]
  wire [2:0] _GEN_289; // @[DCache.scala 765:37:freechips.rocketchip.system.DefaultRV32Config.fir@195480.6]
  wire  _GEN_290; // @[DCache.scala 765:37:freechips.rocketchip.system.DefaultRV32Config.fir@195480.6]
  wire [32:0] _GEN_293; // @[DCache.scala 761:44:freechips.rocketchip.system.DefaultRV32Config.fir@195473.4]
  wire [2:0] _GEN_294; // @[DCache.scala 761:44:freechips.rocketchip.system.DefaultRV32Config.fir@195473.4]
  wire [2:0] _GEN_296; // @[DCache.scala 772:26:freechips.rocketchip.system.DefaultRV32Config.fir@195488.6]
  wire [2:0] _GEN_298; // @[DCache.scala 770:47:freechips.rocketchip.system.DefaultRV32Config.fir@195486.4]
  wire [2:0] _GEN_302; // @[DCache.scala 774:48:freechips.rocketchip.system.DefaultRV32Config.fir@195493.4]
  wire [2:0] _GEN_311; // @[DCache.scala 779:48:freechips.rocketchip.system.DefaultRV32Config.fir@195501.4]
  wire  _T_2434; // @[DCache.scala 792:29:freechips.rocketchip.system.DefaultRV32Config.fir@195546.6]
  wire  _GEN_319; // @[DCache.scala 792:41:freechips.rocketchip.system.DefaultRV32Config.fir@195547.6]
  wire [1:0] newCoh_state; // @[DCache.scala 783:81:freechips.rocketchip.system.DefaultRV32Config.fir@195510.4]
  wire  _T_2436; // @[DCache.scala 803:60:freechips.rocketchip.system.DefaultRV32Config.fir@195557.4]
  wire [11:0] _T_2439; // @[DCache.scala 806:55:freechips.rocketchip.system.DefaultRV32Config.fir@195563.4]
  wire [5:0] _T_2441; // @[DCache.scala 806:117:freechips.rocketchip.system.DefaultRV32Config.fir@195565.4]
  wire [11:0] _GEN_381; // @[DCache.scala 806:72:freechips.rocketchip.system.DefaultRV32Config.fir@195566.4]
  wire  _T_2446; // @[package.scala 15:47:freechips.rocketchip.system.DefaultRV32Config.fir@195573.4]
  wire  _T_2455; // @[Decoupled.scala 40:37:freechips.rocketchip.system.DefaultRV32Config.fir@195591.4]
  wire  _T_2462; // @[DCache.scala 829:57:freechips.rocketchip.system.DefaultRV32Config.fir@195606.4]
  wire  _T_2463; // @[DCache.scala 829:94:freechips.rocketchip.system.DefaultRV32Config.fir@195607.4]
  wire  _T_2465; // @[DCache.scala 829:115:freechips.rocketchip.system.DefaultRV32Config.fir@195609.4]
  reg  _T_2470; // @[DCache.scala 832:32:freechips.rocketchip.system.DefaultRV32Config.fir@195616.4]
  reg  doUncachedResp; // @[DCache.scala 847:27:freechips.rocketchip.system.DefaultRV32Config.fir@195643.4]
  wire  _T_2483; // @[DCache.scala 851:11:freechips.rocketchip.system.DefaultRV32Config.fir@195656.6]
  wire  _T_2484; // @[DCache.scala 851:11:freechips.rocketchip.system.DefaultRV32Config.fir@195657.6]
  wire [15:0] _T_2491; // @[AMOALU.scala 39:24:freechips.rocketchip.system.DefaultRV32Config.fir@195674.4]
  wire  _T_2494; // @[AMOALU.scala 42:26:freechips.rocketchip.system.DefaultRV32Config.fir@195677.4]
  wire  _T_2497; // @[AMOALU.scala 42:76:freechips.rocketchip.system.DefaultRV32Config.fir@195680.4]
  wire [15:0] _T_2499; // @[Bitwise.scala 72:12:freechips.rocketchip.system.DefaultRV32Config.fir@195682.4]
  wire [15:0] _T_2501; // @[AMOALU.scala 42:20:freechips.rocketchip.system.DefaultRV32Config.fir@195684.4]
  wire [31:0] _T_2502; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@195685.4]
  wire [7:0] _T_2506; // @[AMOALU.scala 39:24:freechips.rocketchip.system.DefaultRV32Config.fir@195689.4]
  wire [7:0] _T_2508; // @[AMOALU.scala 41:23:freechips.rocketchip.system.DefaultRV32Config.fir@195691.4]
  wire  _T_2509; // @[AMOALU.scala 42:26:freechips.rocketchip.system.DefaultRV32Config.fir@195692.4]
  wire  _T_2510; // @[AMOALU.scala 42:38:freechips.rocketchip.system.DefaultRV32Config.fir@195693.4]
  wire  _T_2512; // @[AMOALU.scala 42:76:freechips.rocketchip.system.DefaultRV32Config.fir@195695.4]
  wire [23:0] _T_2514; // @[Bitwise.scala 72:12:freechips.rocketchip.system.DefaultRV32Config.fir@195697.4]
  wire [23:0] _T_2516; // @[AMOALU.scala 42:20:freechips.rocketchip.system.DefaultRV32Config.fir@195699.4]
  wire [31:0] _T_2517; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@195700.4]
  wire [31:0] _GEN_382; // @[DCache.scala 873:41:freechips.rocketchip.system.DefaultRV32Config.fir@195701.4]
  reg  resetting; // @[DCache.scala 906:26:freechips.rocketchip.system.DefaultRV32Config.fir@195718.4]
  reg  _T_2523; // @[DCache.scala 908:18:freechips.rocketchip.system.DefaultRV32Config.fir@195720.4]
  wire  _GEN_337; // @[DCache.scala 908:27:freechips.rocketchip.system.DefaultRV32Config.fir@195722.4]
  reg [7:0] flushCounter; // @[DCache.scala 909:25:freechips.rocketchip.system.DefaultRV32Config.fir@195725.4]
  wire [8:0] flushCounterNext; // @[DCache.scala 910:39:freechips.rocketchip.system.DefaultRV32Config.fir@195726.4]
  wire  flushDone; // @[DCache.scala 911:57:freechips.rocketchip.system.DefaultRV32Config.fir@195728.4]
  wire [11:0] _T_2542; // @[DCache.scala 919:98:freechips.rocketchip.system.DefaultRV32Config.fir@195751.4]
  wire [8:0] _GEN_339; // @[DCache.scala 952:20:freechips.rocketchip.system.DefaultRV32Config.fir@195771.4]
  reg [9:0] _T_2604; // @[Edges.scala 230:27:freechips.rocketchip.system.DefaultRV32Config.fir@195837.4]
  wire [9:0] _T_2606; // @[Edges.scala 231:28:freechips.rocketchip.system.DefaultRV32Config.fir@195839.4]
  wire  _T_2607; // @[Edges.scala 232:25:freechips.rocketchip.system.DefaultRV32Config.fir@195840.4]
  wire  _T_2608; // @[Edges.scala 233:25:freechips.rocketchip.system.DefaultRV32Config.fir@195841.4]
  wire  _T_2610; // @[Edges.scala 233:37:freechips.rocketchip.system.DefaultRV32Config.fir@195843.4]
  wire  _T_2725; // @[DCache.scala 1028:35:freechips.rocketchip.system.DefaultRV32Config.fir@195977.4]
  wire  _GEN_385; // @[DCache.scala 620:13:freechips.rocketchip.system.DefaultRV32Config.fir@195113.10]
  wire  _GEN_388; // @[DCache.scala 630:17:freechips.rocketchip.system.DefaultRV32Config.fir@195132.14]
  wire  _GEN_389; // @[DCache.scala 630:17:freechips.rocketchip.system.DefaultRV32Config.fir@195132.14]
  wire  _GEN_390; // @[DCache.scala 630:17:freechips.rocketchip.system.DefaultRV32Config.fir@195132.14]
  wire  _GEN_398; // @[DCache.scala 651:13:freechips.rocketchip.system.DefaultRV32Config.fir@195158.14]
  wire  _GEN_399; // @[DCache.scala 651:13:freechips.rocketchip.system.DefaultRV32Config.fir@195158.14]
  OptimizationBarrier tlb_OptimizationBarrier ( // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@176907.4]
    .io_x_ppn(tlb_OptimizationBarrier_io_x_ppn),
    .io_x_u(tlb_OptimizationBarrier_io_x_u),
    .io_x_ae(tlb_OptimizationBarrier_io_x_ae),
    .io_x_sw(tlb_OptimizationBarrier_io_x_sw),
    .io_x_sx(tlb_OptimizationBarrier_io_x_sx),
    .io_x_sr(tlb_OptimizationBarrier_io_x_sr),
    .io_x_pw(tlb_OptimizationBarrier_io_x_pw),
    .io_x_px(tlb_OptimizationBarrier_io_x_px),
    .io_x_pr(tlb_OptimizationBarrier_io_x_pr),
    .io_x_ppp(tlb_OptimizationBarrier_io_x_ppp),
    .io_x_pal(tlb_OptimizationBarrier_io_x_pal),
    .io_x_paa(tlb_OptimizationBarrier_io_x_paa),
    .io_x_eff(tlb_OptimizationBarrier_io_x_eff),
    .io_x_c(tlb_OptimizationBarrier_io_x_c),
    .io_y_ppn(tlb_OptimizationBarrier_io_y_ppn),
    .io_y_u(tlb_OptimizationBarrier_io_y_u),
    .io_y_ae(tlb_OptimizationBarrier_io_y_ae),
    .io_y_sw(tlb_OptimizationBarrier_io_y_sw),
    .io_y_sx(tlb_OptimizationBarrier_io_y_sx),
    .io_y_sr(tlb_OptimizationBarrier_io_y_sr),
    .io_y_pw(tlb_OptimizationBarrier_io_y_pw),
    .io_y_px(tlb_OptimizationBarrier_io_y_px),
    .io_y_pr(tlb_OptimizationBarrier_io_y_pr),
    .io_y_ppp(tlb_OptimizationBarrier_io_y_ppp),
    .io_y_pal(tlb_OptimizationBarrier_io_y_pal),
    .io_y_paa(tlb_OptimizationBarrier_io_y_paa),
    .io_y_eff(tlb_OptimizationBarrier_io_y_eff),
    .io_y_c(tlb_OptimizationBarrier_io_y_c)
  );
  PMPChecker tlb_pmp ( // @[TLB.scala 190:19:freechips.rocketchip.system.DefaultRV32Config.fir@176928.4]
    .io_prv(tlb_pmp_io_prv),
    .io_pmp_0_cfg_l(tlb_pmp_io_pmp_0_cfg_l),
    .io_pmp_0_cfg_a(tlb_pmp_io_pmp_0_cfg_a),
    .io_pmp_0_cfg_x(tlb_pmp_io_pmp_0_cfg_x),
    .io_pmp_0_cfg_w(tlb_pmp_io_pmp_0_cfg_w),
    .io_pmp_0_cfg_r(tlb_pmp_io_pmp_0_cfg_r),
    .io_pmp_0_addr(tlb_pmp_io_pmp_0_addr),
    .io_pmp_0_mask(tlb_pmp_io_pmp_0_mask),
    .io_pmp_1_cfg_l(tlb_pmp_io_pmp_1_cfg_l),
    .io_pmp_1_cfg_a(tlb_pmp_io_pmp_1_cfg_a),
    .io_pmp_1_cfg_x(tlb_pmp_io_pmp_1_cfg_x),
    .io_pmp_1_cfg_w(tlb_pmp_io_pmp_1_cfg_w),
    .io_pmp_1_cfg_r(tlb_pmp_io_pmp_1_cfg_r),
    .io_pmp_1_addr(tlb_pmp_io_pmp_1_addr),
    .io_pmp_1_mask(tlb_pmp_io_pmp_1_mask),
    .io_pmp_2_cfg_l(tlb_pmp_io_pmp_2_cfg_l),
    .io_pmp_2_cfg_a(tlb_pmp_io_pmp_2_cfg_a),
    .io_pmp_2_cfg_x(tlb_pmp_io_pmp_2_cfg_x),
    .io_pmp_2_cfg_w(tlb_pmp_io_pmp_2_cfg_w),
    .io_pmp_2_cfg_r(tlb_pmp_io_pmp_2_cfg_r),
    .io_pmp_2_addr(tlb_pmp_io_pmp_2_addr),
    .io_pmp_2_mask(tlb_pmp_io_pmp_2_mask),
    .io_pmp_3_cfg_l(tlb_pmp_io_pmp_3_cfg_l),
    .io_pmp_3_cfg_a(tlb_pmp_io_pmp_3_cfg_a),
    .io_pmp_3_cfg_x(tlb_pmp_io_pmp_3_cfg_x),
    .io_pmp_3_cfg_w(tlb_pmp_io_pmp_3_cfg_w),
    .io_pmp_3_cfg_r(tlb_pmp_io_pmp_3_cfg_r),
    .io_pmp_3_addr(tlb_pmp_io_pmp_3_addr),
    .io_pmp_3_mask(tlb_pmp_io_pmp_3_mask),
    .io_pmp_4_cfg_l(tlb_pmp_io_pmp_4_cfg_l),
    .io_pmp_4_cfg_a(tlb_pmp_io_pmp_4_cfg_a),
    .io_pmp_4_cfg_x(tlb_pmp_io_pmp_4_cfg_x),
    .io_pmp_4_cfg_w(tlb_pmp_io_pmp_4_cfg_w),
    .io_pmp_4_cfg_r(tlb_pmp_io_pmp_4_cfg_r),
    .io_pmp_4_addr(tlb_pmp_io_pmp_4_addr),
    .io_pmp_4_mask(tlb_pmp_io_pmp_4_mask),
    .io_pmp_5_cfg_l(tlb_pmp_io_pmp_5_cfg_l),
    .io_pmp_5_cfg_a(tlb_pmp_io_pmp_5_cfg_a),
    .io_pmp_5_cfg_x(tlb_pmp_io_pmp_5_cfg_x),
    .io_pmp_5_cfg_w(tlb_pmp_io_pmp_5_cfg_w),
    .io_pmp_5_cfg_r(tlb_pmp_io_pmp_5_cfg_r),
    .io_pmp_5_addr(tlb_pmp_io_pmp_5_addr),
    .io_pmp_5_mask(tlb_pmp_io_pmp_5_mask),
    .io_pmp_6_cfg_l(tlb_pmp_io_pmp_6_cfg_l),
    .io_pmp_6_cfg_a(tlb_pmp_io_pmp_6_cfg_a),
    .io_pmp_6_cfg_x(tlb_pmp_io_pmp_6_cfg_x),
    .io_pmp_6_cfg_w(tlb_pmp_io_pmp_6_cfg_w),
    .io_pmp_6_cfg_r(tlb_pmp_io_pmp_6_cfg_r),
    .io_pmp_6_addr(tlb_pmp_io_pmp_6_addr),
    .io_pmp_6_mask(tlb_pmp_io_pmp_6_mask),
    .io_pmp_7_cfg_l(tlb_pmp_io_pmp_7_cfg_l),
    .io_pmp_7_cfg_a(tlb_pmp_io_pmp_7_cfg_a),
    .io_pmp_7_cfg_x(tlb_pmp_io_pmp_7_cfg_x),
    .io_pmp_7_cfg_w(tlb_pmp_io_pmp_7_cfg_w),
    .io_pmp_7_cfg_r(tlb_pmp_io_pmp_7_cfg_r),
    .io_pmp_7_addr(tlb_pmp_io_pmp_7_addr),
    .io_pmp_7_mask(tlb_pmp_io_pmp_7_mask),
    .io_addr(tlb_pmp_io_addr),
    .io_r(tlb_pmp_io_r),
    .io_w(tlb_pmp_io_w),
    .io_x(tlb_pmp_io_x)
  );
  OptimizationBarrier tlb_OptimizationBarrier_1 ( // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@177629.4]
    .io_x_ppn(tlb_OptimizationBarrier_1_io_x_ppn),
    .io_x_u(tlb_OptimizationBarrier_1_io_x_u),
    .io_x_ae(tlb_OptimizationBarrier_1_io_x_ae),
    .io_x_sw(tlb_OptimizationBarrier_1_io_x_sw),
    .io_x_sx(tlb_OptimizationBarrier_1_io_x_sx),
    .io_x_sr(tlb_OptimizationBarrier_1_io_x_sr),
    .io_x_pw(tlb_OptimizationBarrier_1_io_x_pw),
    .io_x_px(tlb_OptimizationBarrier_1_io_x_px),
    .io_x_pr(tlb_OptimizationBarrier_1_io_x_pr),
    .io_x_ppp(tlb_OptimizationBarrier_1_io_x_ppp),
    .io_x_pal(tlb_OptimizationBarrier_1_io_x_pal),
    .io_x_paa(tlb_OptimizationBarrier_1_io_x_paa),
    .io_x_eff(tlb_OptimizationBarrier_1_io_x_eff),
    .io_x_c(tlb_OptimizationBarrier_1_io_x_c),
    .io_y_ppn(tlb_OptimizationBarrier_1_io_y_ppn),
    .io_y_u(tlb_OptimizationBarrier_1_io_y_u),
    .io_y_ae(tlb_OptimizationBarrier_1_io_y_ae),
    .io_y_sw(tlb_OptimizationBarrier_1_io_y_sw),
    .io_y_sx(tlb_OptimizationBarrier_1_io_y_sx),
    .io_y_sr(tlb_OptimizationBarrier_1_io_y_sr),
    .io_y_pw(tlb_OptimizationBarrier_1_io_y_pw),
    .io_y_px(tlb_OptimizationBarrier_1_io_y_px),
    .io_y_pr(tlb_OptimizationBarrier_1_io_y_pr),
    .io_y_ppp(tlb_OptimizationBarrier_1_io_y_ppp),
    .io_y_pal(tlb_OptimizationBarrier_1_io_y_pal),
    .io_y_paa(tlb_OptimizationBarrier_1_io_y_paa),
    .io_y_eff(tlb_OptimizationBarrier_1_io_y_eff),
    .io_y_c(tlb_OptimizationBarrier_1_io_y_c)
  );
  OptimizationBarrier tlb_OptimizationBarrier_2 ( // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@177672.4]
    .io_x_ppn(tlb_OptimizationBarrier_2_io_x_ppn),
    .io_x_u(tlb_OptimizationBarrier_2_io_x_u),
    .io_x_ae(tlb_OptimizationBarrier_2_io_x_ae),
    .io_x_sw(tlb_OptimizationBarrier_2_io_x_sw),
    .io_x_sx(tlb_OptimizationBarrier_2_io_x_sx),
    .io_x_sr(tlb_OptimizationBarrier_2_io_x_sr),
    .io_x_pw(tlb_OptimizationBarrier_2_io_x_pw),
    .io_x_px(tlb_OptimizationBarrier_2_io_x_px),
    .io_x_pr(tlb_OptimizationBarrier_2_io_x_pr),
    .io_x_ppp(tlb_OptimizationBarrier_2_io_x_ppp),
    .io_x_pal(tlb_OptimizationBarrier_2_io_x_pal),
    .io_x_paa(tlb_OptimizationBarrier_2_io_x_paa),
    .io_x_eff(tlb_OptimizationBarrier_2_io_x_eff),
    .io_x_c(tlb_OptimizationBarrier_2_io_x_c),
    .io_y_ppn(tlb_OptimizationBarrier_2_io_y_ppn),
    .io_y_u(tlb_OptimizationBarrier_2_io_y_u),
    .io_y_ae(tlb_OptimizationBarrier_2_io_y_ae),
    .io_y_sw(tlb_OptimizationBarrier_2_io_y_sw),
    .io_y_sx(tlb_OptimizationBarrier_2_io_y_sx),
    .io_y_sr(tlb_OptimizationBarrier_2_io_y_sr),
    .io_y_pw(tlb_OptimizationBarrier_2_io_y_pw),
    .io_y_px(tlb_OptimizationBarrier_2_io_y_px),
    .io_y_pr(tlb_OptimizationBarrier_2_io_y_pr),
    .io_y_ppp(tlb_OptimizationBarrier_2_io_y_ppp),
    .io_y_pal(tlb_OptimizationBarrier_2_io_y_pal),
    .io_y_paa(tlb_OptimizationBarrier_2_io_y_paa),
    .io_y_eff(tlb_OptimizationBarrier_2_io_y_eff),
    .io_y_c(tlb_OptimizationBarrier_2_io_y_c)
  );
  OptimizationBarrier tlb_OptimizationBarrier_3 ( // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@177715.4]
    .io_x_ppn(tlb_OptimizationBarrier_3_io_x_ppn),
    .io_x_u(tlb_OptimizationBarrier_3_io_x_u),
    .io_x_ae(tlb_OptimizationBarrier_3_io_x_ae),
    .io_x_sw(tlb_OptimizationBarrier_3_io_x_sw),
    .io_x_sx(tlb_OptimizationBarrier_3_io_x_sx),
    .io_x_sr(tlb_OptimizationBarrier_3_io_x_sr),
    .io_x_pw(tlb_OptimizationBarrier_3_io_x_pw),
    .io_x_px(tlb_OptimizationBarrier_3_io_x_px),
    .io_x_pr(tlb_OptimizationBarrier_3_io_x_pr),
    .io_x_ppp(tlb_OptimizationBarrier_3_io_x_ppp),
    .io_x_pal(tlb_OptimizationBarrier_3_io_x_pal),
    .io_x_paa(tlb_OptimizationBarrier_3_io_x_paa),
    .io_x_eff(tlb_OptimizationBarrier_3_io_x_eff),
    .io_x_c(tlb_OptimizationBarrier_3_io_x_c),
    .io_y_ppn(tlb_OptimizationBarrier_3_io_y_ppn),
    .io_y_u(tlb_OptimizationBarrier_3_io_y_u),
    .io_y_ae(tlb_OptimizationBarrier_3_io_y_ae),
    .io_y_sw(tlb_OptimizationBarrier_3_io_y_sw),
    .io_y_sx(tlb_OptimizationBarrier_3_io_y_sx),
    .io_y_sr(tlb_OptimizationBarrier_3_io_y_sr),
    .io_y_pw(tlb_OptimizationBarrier_3_io_y_pw),
    .io_y_px(tlb_OptimizationBarrier_3_io_y_px),
    .io_y_pr(tlb_OptimizationBarrier_3_io_y_pr),
    .io_y_ppp(tlb_OptimizationBarrier_3_io_y_ppp),
    .io_y_pal(tlb_OptimizationBarrier_3_io_y_pal),
    .io_y_paa(tlb_OptimizationBarrier_3_io_y_paa),
    .io_y_eff(tlb_OptimizationBarrier_3_io_y_eff),
    .io_y_c(tlb_OptimizationBarrier_3_io_y_c)
  );
  OptimizationBarrier tlb_OptimizationBarrier_4 ( // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@177758.4]
    .io_x_ppn(tlb_OptimizationBarrier_4_io_x_ppn),
    .io_x_u(tlb_OptimizationBarrier_4_io_x_u),
    .io_x_ae(tlb_OptimizationBarrier_4_io_x_ae),
    .io_x_sw(tlb_OptimizationBarrier_4_io_x_sw),
    .io_x_sx(tlb_OptimizationBarrier_4_io_x_sx),
    .io_x_sr(tlb_OptimizationBarrier_4_io_x_sr),
    .io_x_pw(tlb_OptimizationBarrier_4_io_x_pw),
    .io_x_px(tlb_OptimizationBarrier_4_io_x_px),
    .io_x_pr(tlb_OptimizationBarrier_4_io_x_pr),
    .io_x_ppp(tlb_OptimizationBarrier_4_io_x_ppp),
    .io_x_pal(tlb_OptimizationBarrier_4_io_x_pal),
    .io_x_paa(tlb_OptimizationBarrier_4_io_x_paa),
    .io_x_eff(tlb_OptimizationBarrier_4_io_x_eff),
    .io_x_c(tlb_OptimizationBarrier_4_io_x_c),
    .io_y_ppn(tlb_OptimizationBarrier_4_io_y_ppn),
    .io_y_u(tlb_OptimizationBarrier_4_io_y_u),
    .io_y_ae(tlb_OptimizationBarrier_4_io_y_ae),
    .io_y_sw(tlb_OptimizationBarrier_4_io_y_sw),
    .io_y_sx(tlb_OptimizationBarrier_4_io_y_sx),
    .io_y_sr(tlb_OptimizationBarrier_4_io_y_sr),
    .io_y_pw(tlb_OptimizationBarrier_4_io_y_pw),
    .io_y_px(tlb_OptimizationBarrier_4_io_y_px),
    .io_y_pr(tlb_OptimizationBarrier_4_io_y_pr),
    .io_y_ppp(tlb_OptimizationBarrier_4_io_y_ppp),
    .io_y_pal(tlb_OptimizationBarrier_4_io_y_pal),
    .io_y_paa(tlb_OptimizationBarrier_4_io_y_paa),
    .io_y_eff(tlb_OptimizationBarrier_4_io_y_eff),
    .io_y_c(tlb_OptimizationBarrier_4_io_y_c)
  );
  OptimizationBarrier tlb_OptimizationBarrier_5 ( // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@177801.4]
    .io_x_ppn(tlb_OptimizationBarrier_5_io_x_ppn),
    .io_x_u(tlb_OptimizationBarrier_5_io_x_u),
    .io_x_ae(tlb_OptimizationBarrier_5_io_x_ae),
    .io_x_sw(tlb_OptimizationBarrier_5_io_x_sw),
    .io_x_sx(tlb_OptimizationBarrier_5_io_x_sx),
    .io_x_sr(tlb_OptimizationBarrier_5_io_x_sr),
    .io_x_pw(tlb_OptimizationBarrier_5_io_x_pw),
    .io_x_px(tlb_OptimizationBarrier_5_io_x_px),
    .io_x_pr(tlb_OptimizationBarrier_5_io_x_pr),
    .io_x_ppp(tlb_OptimizationBarrier_5_io_x_ppp),
    .io_x_pal(tlb_OptimizationBarrier_5_io_x_pal),
    .io_x_paa(tlb_OptimizationBarrier_5_io_x_paa),
    .io_x_eff(tlb_OptimizationBarrier_5_io_x_eff),
    .io_x_c(tlb_OptimizationBarrier_5_io_x_c),
    .io_y_ppn(tlb_OptimizationBarrier_5_io_y_ppn),
    .io_y_u(tlb_OptimizationBarrier_5_io_y_u),
    .io_y_ae(tlb_OptimizationBarrier_5_io_y_ae),
    .io_y_sw(tlb_OptimizationBarrier_5_io_y_sw),
    .io_y_sx(tlb_OptimizationBarrier_5_io_y_sx),
    .io_y_sr(tlb_OptimizationBarrier_5_io_y_sr),
    .io_y_pw(tlb_OptimizationBarrier_5_io_y_pw),
    .io_y_px(tlb_OptimizationBarrier_5_io_y_px),
    .io_y_pr(tlb_OptimizationBarrier_5_io_y_pr),
    .io_y_ppp(tlb_OptimizationBarrier_5_io_y_ppp),
    .io_y_pal(tlb_OptimizationBarrier_5_io_y_pal),
    .io_y_paa(tlb_OptimizationBarrier_5_io_y_paa),
    .io_y_eff(tlb_OptimizationBarrier_5_io_y_eff),
    .io_y_c(tlb_OptimizationBarrier_5_io_y_c)
  );
  OptimizationBarrier tlb_OptimizationBarrier_6 ( // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@177844.4]
    .io_x_ppn(tlb_OptimizationBarrier_6_io_x_ppn),
    .io_x_u(tlb_OptimizationBarrier_6_io_x_u),
    .io_x_ae(tlb_OptimizationBarrier_6_io_x_ae),
    .io_x_sw(tlb_OptimizationBarrier_6_io_x_sw),
    .io_x_sx(tlb_OptimizationBarrier_6_io_x_sx),
    .io_x_sr(tlb_OptimizationBarrier_6_io_x_sr),
    .io_x_pw(tlb_OptimizationBarrier_6_io_x_pw),
    .io_x_px(tlb_OptimizationBarrier_6_io_x_px),
    .io_x_pr(tlb_OptimizationBarrier_6_io_x_pr),
    .io_x_ppp(tlb_OptimizationBarrier_6_io_x_ppp),
    .io_x_pal(tlb_OptimizationBarrier_6_io_x_pal),
    .io_x_paa(tlb_OptimizationBarrier_6_io_x_paa),
    .io_x_eff(tlb_OptimizationBarrier_6_io_x_eff),
    .io_x_c(tlb_OptimizationBarrier_6_io_x_c),
    .io_y_ppn(tlb_OptimizationBarrier_6_io_y_ppn),
    .io_y_u(tlb_OptimizationBarrier_6_io_y_u),
    .io_y_ae(tlb_OptimizationBarrier_6_io_y_ae),
    .io_y_sw(tlb_OptimizationBarrier_6_io_y_sw),
    .io_y_sx(tlb_OptimizationBarrier_6_io_y_sx),
    .io_y_sr(tlb_OptimizationBarrier_6_io_y_sr),
    .io_y_pw(tlb_OptimizationBarrier_6_io_y_pw),
    .io_y_px(tlb_OptimizationBarrier_6_io_y_px),
    .io_y_pr(tlb_OptimizationBarrier_6_io_y_pr),
    .io_y_ppp(tlb_OptimizationBarrier_6_io_y_ppp),
    .io_y_pal(tlb_OptimizationBarrier_6_io_y_pal),
    .io_y_paa(tlb_OptimizationBarrier_6_io_y_paa),
    .io_y_eff(tlb_OptimizationBarrier_6_io_y_eff),
    .io_y_c(tlb_OptimizationBarrier_6_io_y_c)
  );
  OptimizationBarrier tlb_OptimizationBarrier_7 ( // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@177887.4]
    .io_x_ppn(tlb_OptimizationBarrier_7_io_x_ppn),
    .io_x_u(tlb_OptimizationBarrier_7_io_x_u),
    .io_x_ae(tlb_OptimizationBarrier_7_io_x_ae),
    .io_x_sw(tlb_OptimizationBarrier_7_io_x_sw),
    .io_x_sx(tlb_OptimizationBarrier_7_io_x_sx),
    .io_x_sr(tlb_OptimizationBarrier_7_io_x_sr),
    .io_x_pw(tlb_OptimizationBarrier_7_io_x_pw),
    .io_x_px(tlb_OptimizationBarrier_7_io_x_px),
    .io_x_pr(tlb_OptimizationBarrier_7_io_x_pr),
    .io_x_ppp(tlb_OptimizationBarrier_7_io_x_ppp),
    .io_x_pal(tlb_OptimizationBarrier_7_io_x_pal),
    .io_x_paa(tlb_OptimizationBarrier_7_io_x_paa),
    .io_x_eff(tlb_OptimizationBarrier_7_io_x_eff),
    .io_x_c(tlb_OptimizationBarrier_7_io_x_c),
    .io_y_ppn(tlb_OptimizationBarrier_7_io_y_ppn),
    .io_y_u(tlb_OptimizationBarrier_7_io_y_u),
    .io_y_ae(tlb_OptimizationBarrier_7_io_y_ae),
    .io_y_sw(tlb_OptimizationBarrier_7_io_y_sw),
    .io_y_sx(tlb_OptimizationBarrier_7_io_y_sx),
    .io_y_sr(tlb_OptimizationBarrier_7_io_y_sr),
    .io_y_pw(tlb_OptimizationBarrier_7_io_y_pw),
    .io_y_px(tlb_OptimizationBarrier_7_io_y_px),
    .io_y_pr(tlb_OptimizationBarrier_7_io_y_pr),
    .io_y_ppp(tlb_OptimizationBarrier_7_io_y_ppp),
    .io_y_pal(tlb_OptimizationBarrier_7_io_y_pal),
    .io_y_paa(tlb_OptimizationBarrier_7_io_y_paa),
    .io_y_eff(tlb_OptimizationBarrier_7_io_y_eff),
    .io_y_c(tlb_OptimizationBarrier_7_io_y_c)
  );
  OptimizationBarrier tlb_OptimizationBarrier_8 ( // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@177930.4]
    .io_x_ppn(tlb_OptimizationBarrier_8_io_x_ppn),
    .io_x_u(tlb_OptimizationBarrier_8_io_x_u),
    .io_x_ae(tlb_OptimizationBarrier_8_io_x_ae),
    .io_x_sw(tlb_OptimizationBarrier_8_io_x_sw),
    .io_x_sx(tlb_OptimizationBarrier_8_io_x_sx),
    .io_x_sr(tlb_OptimizationBarrier_8_io_x_sr),
    .io_x_pw(tlb_OptimizationBarrier_8_io_x_pw),
    .io_x_px(tlb_OptimizationBarrier_8_io_x_px),
    .io_x_pr(tlb_OptimizationBarrier_8_io_x_pr),
    .io_x_ppp(tlb_OptimizationBarrier_8_io_x_ppp),
    .io_x_pal(tlb_OptimizationBarrier_8_io_x_pal),
    .io_x_paa(tlb_OptimizationBarrier_8_io_x_paa),
    .io_x_eff(tlb_OptimizationBarrier_8_io_x_eff),
    .io_x_c(tlb_OptimizationBarrier_8_io_x_c),
    .io_y_ppn(tlb_OptimizationBarrier_8_io_y_ppn),
    .io_y_u(tlb_OptimizationBarrier_8_io_y_u),
    .io_y_ae(tlb_OptimizationBarrier_8_io_y_ae),
    .io_y_sw(tlb_OptimizationBarrier_8_io_y_sw),
    .io_y_sx(tlb_OptimizationBarrier_8_io_y_sx),
    .io_y_sr(tlb_OptimizationBarrier_8_io_y_sr),
    .io_y_pw(tlb_OptimizationBarrier_8_io_y_pw),
    .io_y_px(tlb_OptimizationBarrier_8_io_y_px),
    .io_y_pr(tlb_OptimizationBarrier_8_io_y_pr),
    .io_y_ppp(tlb_OptimizationBarrier_8_io_y_ppp),
    .io_y_pal(tlb_OptimizationBarrier_8_io_y_pal),
    .io_y_paa(tlb_OptimizationBarrier_8_io_y_paa),
    .io_y_eff(tlb_OptimizationBarrier_8_io_y_eff),
    .io_y_c(tlb_OptimizationBarrier_8_io_y_c)
  );
  OptimizationBarrier tlb_OptimizationBarrier_9 ( // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@177972.4]
    .io_x_ppn(tlb_OptimizationBarrier_9_io_x_ppn),
    .io_x_u(tlb_OptimizationBarrier_9_io_x_u),
    .io_x_ae(tlb_OptimizationBarrier_9_io_x_ae),
    .io_x_sw(tlb_OptimizationBarrier_9_io_x_sw),
    .io_x_sx(tlb_OptimizationBarrier_9_io_x_sx),
    .io_x_sr(tlb_OptimizationBarrier_9_io_x_sr),
    .io_x_pw(tlb_OptimizationBarrier_9_io_x_pw),
    .io_x_px(tlb_OptimizationBarrier_9_io_x_px),
    .io_x_pr(tlb_OptimizationBarrier_9_io_x_pr),
    .io_x_ppp(tlb_OptimizationBarrier_9_io_x_ppp),
    .io_x_pal(tlb_OptimizationBarrier_9_io_x_pal),
    .io_x_paa(tlb_OptimizationBarrier_9_io_x_paa),
    .io_x_eff(tlb_OptimizationBarrier_9_io_x_eff),
    .io_x_c(tlb_OptimizationBarrier_9_io_x_c),
    .io_y_ppn(tlb_OptimizationBarrier_9_io_y_ppn),
    .io_y_u(tlb_OptimizationBarrier_9_io_y_u),
    .io_y_ae(tlb_OptimizationBarrier_9_io_y_ae),
    .io_y_sw(tlb_OptimizationBarrier_9_io_y_sw),
    .io_y_sx(tlb_OptimizationBarrier_9_io_y_sx),
    .io_y_sr(tlb_OptimizationBarrier_9_io_y_sr),
    .io_y_pw(tlb_OptimizationBarrier_9_io_y_pw),
    .io_y_px(tlb_OptimizationBarrier_9_io_y_px),
    .io_y_pr(tlb_OptimizationBarrier_9_io_y_pr),
    .io_y_ppp(tlb_OptimizationBarrier_9_io_y_ppp),
    .io_y_pal(tlb_OptimizationBarrier_9_io_y_pal),
    .io_y_paa(tlb_OptimizationBarrier_9_io_y_paa),
    .io_y_eff(tlb_OptimizationBarrier_9_io_y_eff),
    .io_y_c(tlb_OptimizationBarrier_9_io_y_c)
  );
  OptimizationBarrier tlb_OptimizationBarrier_10 ( // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178021.4]
    .io_x_ppn(tlb_OptimizationBarrier_10_io_x_ppn),
    .io_x_u(tlb_OptimizationBarrier_10_io_x_u),
    .io_x_ae(tlb_OptimizationBarrier_10_io_x_ae),
    .io_x_sw(tlb_OptimizationBarrier_10_io_x_sw),
    .io_x_sx(tlb_OptimizationBarrier_10_io_x_sx),
    .io_x_sr(tlb_OptimizationBarrier_10_io_x_sr),
    .io_x_pw(tlb_OptimizationBarrier_10_io_x_pw),
    .io_x_px(tlb_OptimizationBarrier_10_io_x_px),
    .io_x_pr(tlb_OptimizationBarrier_10_io_x_pr),
    .io_x_ppp(tlb_OptimizationBarrier_10_io_x_ppp),
    .io_x_pal(tlb_OptimizationBarrier_10_io_x_pal),
    .io_x_paa(tlb_OptimizationBarrier_10_io_x_paa),
    .io_x_eff(tlb_OptimizationBarrier_10_io_x_eff),
    .io_x_c(tlb_OptimizationBarrier_10_io_x_c),
    .io_y_ppn(tlb_OptimizationBarrier_10_io_y_ppn),
    .io_y_u(tlb_OptimizationBarrier_10_io_y_u),
    .io_y_ae(tlb_OptimizationBarrier_10_io_y_ae),
    .io_y_sw(tlb_OptimizationBarrier_10_io_y_sw),
    .io_y_sx(tlb_OptimizationBarrier_10_io_y_sx),
    .io_y_sr(tlb_OptimizationBarrier_10_io_y_sr),
    .io_y_pw(tlb_OptimizationBarrier_10_io_y_pw),
    .io_y_px(tlb_OptimizationBarrier_10_io_y_px),
    .io_y_pr(tlb_OptimizationBarrier_10_io_y_pr),
    .io_y_ppp(tlb_OptimizationBarrier_10_io_y_ppp),
    .io_y_pal(tlb_OptimizationBarrier_10_io_y_pal),
    .io_y_paa(tlb_OptimizationBarrier_10_io_y_paa),
    .io_y_eff(tlb_OptimizationBarrier_10_io_y_eff),
    .io_y_c(tlb_OptimizationBarrier_10_io_y_c)
  );
  OptimizationBarrier tlb_OptimizationBarrier_11 ( // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178070.4]
    .io_x_ppn(tlb_OptimizationBarrier_11_io_x_ppn),
    .io_x_u(tlb_OptimizationBarrier_11_io_x_u),
    .io_x_ae(tlb_OptimizationBarrier_11_io_x_ae),
    .io_x_sw(tlb_OptimizationBarrier_11_io_x_sw),
    .io_x_sx(tlb_OptimizationBarrier_11_io_x_sx),
    .io_x_sr(tlb_OptimizationBarrier_11_io_x_sr),
    .io_x_pw(tlb_OptimizationBarrier_11_io_x_pw),
    .io_x_px(tlb_OptimizationBarrier_11_io_x_px),
    .io_x_pr(tlb_OptimizationBarrier_11_io_x_pr),
    .io_x_ppp(tlb_OptimizationBarrier_11_io_x_ppp),
    .io_x_pal(tlb_OptimizationBarrier_11_io_x_pal),
    .io_x_paa(tlb_OptimizationBarrier_11_io_x_paa),
    .io_x_eff(tlb_OptimizationBarrier_11_io_x_eff),
    .io_x_c(tlb_OptimizationBarrier_11_io_x_c),
    .io_y_ppn(tlb_OptimizationBarrier_11_io_y_ppn),
    .io_y_u(tlb_OptimizationBarrier_11_io_y_u),
    .io_y_ae(tlb_OptimizationBarrier_11_io_y_ae),
    .io_y_sw(tlb_OptimizationBarrier_11_io_y_sw),
    .io_y_sx(tlb_OptimizationBarrier_11_io_y_sx),
    .io_y_sr(tlb_OptimizationBarrier_11_io_y_sr),
    .io_y_pw(tlb_OptimizationBarrier_11_io_y_pw),
    .io_y_px(tlb_OptimizationBarrier_11_io_y_px),
    .io_y_pr(tlb_OptimizationBarrier_11_io_y_pr),
    .io_y_ppp(tlb_OptimizationBarrier_11_io_y_ppp),
    .io_y_pal(tlb_OptimizationBarrier_11_io_y_pal),
    .io_y_paa(tlb_OptimizationBarrier_11_io_y_paa),
    .io_y_eff(tlb_OptimizationBarrier_11_io_y_eff),
    .io_y_c(tlb_OptimizationBarrier_11_io_y_c)
  );
  OptimizationBarrier tlb_OptimizationBarrier_12 ( // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178119.4]
    .io_x_ppn(tlb_OptimizationBarrier_12_io_x_ppn),
    .io_x_u(tlb_OptimizationBarrier_12_io_x_u),
    .io_x_ae(tlb_OptimizationBarrier_12_io_x_ae),
    .io_x_sw(tlb_OptimizationBarrier_12_io_x_sw),
    .io_x_sx(tlb_OptimizationBarrier_12_io_x_sx),
    .io_x_sr(tlb_OptimizationBarrier_12_io_x_sr),
    .io_x_pw(tlb_OptimizationBarrier_12_io_x_pw),
    .io_x_px(tlb_OptimizationBarrier_12_io_x_px),
    .io_x_pr(tlb_OptimizationBarrier_12_io_x_pr),
    .io_x_ppp(tlb_OptimizationBarrier_12_io_x_ppp),
    .io_x_pal(tlb_OptimizationBarrier_12_io_x_pal),
    .io_x_paa(tlb_OptimizationBarrier_12_io_x_paa),
    .io_x_eff(tlb_OptimizationBarrier_12_io_x_eff),
    .io_x_c(tlb_OptimizationBarrier_12_io_x_c),
    .io_y_ppn(tlb_OptimizationBarrier_12_io_y_ppn),
    .io_y_u(tlb_OptimizationBarrier_12_io_y_u),
    .io_y_ae(tlb_OptimizationBarrier_12_io_y_ae),
    .io_y_sw(tlb_OptimizationBarrier_12_io_y_sw),
    .io_y_sx(tlb_OptimizationBarrier_12_io_y_sx),
    .io_y_sr(tlb_OptimizationBarrier_12_io_y_sr),
    .io_y_pw(tlb_OptimizationBarrier_12_io_y_pw),
    .io_y_px(tlb_OptimizationBarrier_12_io_y_px),
    .io_y_pr(tlb_OptimizationBarrier_12_io_y_pr),
    .io_y_ppp(tlb_OptimizationBarrier_12_io_y_ppp),
    .io_y_pal(tlb_OptimizationBarrier_12_io_y_pal),
    .io_y_paa(tlb_OptimizationBarrier_12_io_y_paa),
    .io_y_eff(tlb_OptimizationBarrier_12_io_y_eff),
    .io_y_c(tlb_OptimizationBarrier_12_io_y_c)
  );
  OptimizationBarrier tlb_OptimizationBarrier_13 ( // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178168.4]
    .io_x_ppn(tlb_OptimizationBarrier_13_io_x_ppn),
    .io_x_u(tlb_OptimizationBarrier_13_io_x_u),
    .io_x_ae(tlb_OptimizationBarrier_13_io_x_ae),
    .io_x_sw(tlb_OptimizationBarrier_13_io_x_sw),
    .io_x_sx(tlb_OptimizationBarrier_13_io_x_sx),
    .io_x_sr(tlb_OptimizationBarrier_13_io_x_sr),
    .io_x_pw(tlb_OptimizationBarrier_13_io_x_pw),
    .io_x_px(tlb_OptimizationBarrier_13_io_x_px),
    .io_x_pr(tlb_OptimizationBarrier_13_io_x_pr),
    .io_x_ppp(tlb_OptimizationBarrier_13_io_x_ppp),
    .io_x_pal(tlb_OptimizationBarrier_13_io_x_pal),
    .io_x_paa(tlb_OptimizationBarrier_13_io_x_paa),
    .io_x_eff(tlb_OptimizationBarrier_13_io_x_eff),
    .io_x_c(tlb_OptimizationBarrier_13_io_x_c),
    .io_y_ppn(tlb_OptimizationBarrier_13_io_y_ppn),
    .io_y_u(tlb_OptimizationBarrier_13_io_y_u),
    .io_y_ae(tlb_OptimizationBarrier_13_io_y_ae),
    .io_y_sw(tlb_OptimizationBarrier_13_io_y_sw),
    .io_y_sx(tlb_OptimizationBarrier_13_io_y_sx),
    .io_y_sr(tlb_OptimizationBarrier_13_io_y_sr),
    .io_y_pw(tlb_OptimizationBarrier_13_io_y_pw),
    .io_y_px(tlb_OptimizationBarrier_13_io_y_px),
    .io_y_pr(tlb_OptimizationBarrier_13_io_y_pr),
    .io_y_ppp(tlb_OptimizationBarrier_13_io_y_ppp),
    .io_y_pal(tlb_OptimizationBarrier_13_io_y_pal),
    .io_y_paa(tlb_OptimizationBarrier_13_io_y_paa),
    .io_y_eff(tlb_OptimizationBarrier_13_io_y_eff),
    .io_y_c(tlb_OptimizationBarrier_13_io_y_c)
  );
  OptimizationBarrier tlb_OptimizationBarrier_14 ( // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178649.4]
    .io_x_ppn(tlb_OptimizationBarrier_14_io_x_ppn),
    .io_x_u(tlb_OptimizationBarrier_14_io_x_u),
    .io_x_ae(tlb_OptimizationBarrier_14_io_x_ae),
    .io_x_sw(tlb_OptimizationBarrier_14_io_x_sw),
    .io_x_sx(tlb_OptimizationBarrier_14_io_x_sx),
    .io_x_sr(tlb_OptimizationBarrier_14_io_x_sr),
    .io_x_pw(tlb_OptimizationBarrier_14_io_x_pw),
    .io_x_px(tlb_OptimizationBarrier_14_io_x_px),
    .io_x_pr(tlb_OptimizationBarrier_14_io_x_pr),
    .io_x_ppp(tlb_OptimizationBarrier_14_io_x_ppp),
    .io_x_pal(tlb_OptimizationBarrier_14_io_x_pal),
    .io_x_paa(tlb_OptimizationBarrier_14_io_x_paa),
    .io_x_eff(tlb_OptimizationBarrier_14_io_x_eff),
    .io_x_c(tlb_OptimizationBarrier_14_io_x_c),
    .io_y_ppn(tlb_OptimizationBarrier_14_io_y_ppn),
    .io_y_u(tlb_OptimizationBarrier_14_io_y_u),
    .io_y_ae(tlb_OptimizationBarrier_14_io_y_ae),
    .io_y_sw(tlb_OptimizationBarrier_14_io_y_sw),
    .io_y_sx(tlb_OptimizationBarrier_14_io_y_sx),
    .io_y_sr(tlb_OptimizationBarrier_14_io_y_sr),
    .io_y_pw(tlb_OptimizationBarrier_14_io_y_pw),
    .io_y_px(tlb_OptimizationBarrier_14_io_y_px),
    .io_y_pr(tlb_OptimizationBarrier_14_io_y_pr),
    .io_y_ppp(tlb_OptimizationBarrier_14_io_y_ppp),
    .io_y_pal(tlb_OptimizationBarrier_14_io_y_pal),
    .io_y_paa(tlb_OptimizationBarrier_14_io_y_paa),
    .io_y_eff(tlb_OptimizationBarrier_14_io_y_eff),
    .io_y_c(tlb_OptimizationBarrier_14_io_y_c)
  );
  OptimizationBarrier tlb_OptimizationBarrier_15 ( // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178692.4]
    .io_x_ppn(tlb_OptimizationBarrier_15_io_x_ppn),
    .io_x_u(tlb_OptimizationBarrier_15_io_x_u),
    .io_x_ae(tlb_OptimizationBarrier_15_io_x_ae),
    .io_x_sw(tlb_OptimizationBarrier_15_io_x_sw),
    .io_x_sx(tlb_OptimizationBarrier_15_io_x_sx),
    .io_x_sr(tlb_OptimizationBarrier_15_io_x_sr),
    .io_x_pw(tlb_OptimizationBarrier_15_io_x_pw),
    .io_x_px(tlb_OptimizationBarrier_15_io_x_px),
    .io_x_pr(tlb_OptimizationBarrier_15_io_x_pr),
    .io_x_ppp(tlb_OptimizationBarrier_15_io_x_ppp),
    .io_x_pal(tlb_OptimizationBarrier_15_io_x_pal),
    .io_x_paa(tlb_OptimizationBarrier_15_io_x_paa),
    .io_x_eff(tlb_OptimizationBarrier_15_io_x_eff),
    .io_x_c(tlb_OptimizationBarrier_15_io_x_c),
    .io_y_ppn(tlb_OptimizationBarrier_15_io_y_ppn),
    .io_y_u(tlb_OptimizationBarrier_15_io_y_u),
    .io_y_ae(tlb_OptimizationBarrier_15_io_y_ae),
    .io_y_sw(tlb_OptimizationBarrier_15_io_y_sw),
    .io_y_sx(tlb_OptimizationBarrier_15_io_y_sx),
    .io_y_sr(tlb_OptimizationBarrier_15_io_y_sr),
    .io_y_pw(tlb_OptimizationBarrier_15_io_y_pw),
    .io_y_px(tlb_OptimizationBarrier_15_io_y_px),
    .io_y_pr(tlb_OptimizationBarrier_15_io_y_pr),
    .io_y_ppp(tlb_OptimizationBarrier_15_io_y_ppp),
    .io_y_pal(tlb_OptimizationBarrier_15_io_y_pal),
    .io_y_paa(tlb_OptimizationBarrier_15_io_y_paa),
    .io_y_eff(tlb_OptimizationBarrier_15_io_y_eff),
    .io_y_c(tlb_OptimizationBarrier_15_io_y_c)
  );
  OptimizationBarrier tlb_OptimizationBarrier_16 ( // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178735.4]
    .io_x_ppn(tlb_OptimizationBarrier_16_io_x_ppn),
    .io_x_u(tlb_OptimizationBarrier_16_io_x_u),
    .io_x_ae(tlb_OptimizationBarrier_16_io_x_ae),
    .io_x_sw(tlb_OptimizationBarrier_16_io_x_sw),
    .io_x_sx(tlb_OptimizationBarrier_16_io_x_sx),
    .io_x_sr(tlb_OptimizationBarrier_16_io_x_sr),
    .io_x_pw(tlb_OptimizationBarrier_16_io_x_pw),
    .io_x_px(tlb_OptimizationBarrier_16_io_x_px),
    .io_x_pr(tlb_OptimizationBarrier_16_io_x_pr),
    .io_x_ppp(tlb_OptimizationBarrier_16_io_x_ppp),
    .io_x_pal(tlb_OptimizationBarrier_16_io_x_pal),
    .io_x_paa(tlb_OptimizationBarrier_16_io_x_paa),
    .io_x_eff(tlb_OptimizationBarrier_16_io_x_eff),
    .io_x_c(tlb_OptimizationBarrier_16_io_x_c),
    .io_y_ppn(tlb_OptimizationBarrier_16_io_y_ppn),
    .io_y_u(tlb_OptimizationBarrier_16_io_y_u),
    .io_y_ae(tlb_OptimizationBarrier_16_io_y_ae),
    .io_y_sw(tlb_OptimizationBarrier_16_io_y_sw),
    .io_y_sx(tlb_OptimizationBarrier_16_io_y_sx),
    .io_y_sr(tlb_OptimizationBarrier_16_io_y_sr),
    .io_y_pw(tlb_OptimizationBarrier_16_io_y_pw),
    .io_y_px(tlb_OptimizationBarrier_16_io_y_px),
    .io_y_pr(tlb_OptimizationBarrier_16_io_y_pr),
    .io_y_ppp(tlb_OptimizationBarrier_16_io_y_ppp),
    .io_y_pal(tlb_OptimizationBarrier_16_io_y_pal),
    .io_y_paa(tlb_OptimizationBarrier_16_io_y_paa),
    .io_y_eff(tlb_OptimizationBarrier_16_io_y_eff),
    .io_y_c(tlb_OptimizationBarrier_16_io_y_c)
  );
  OptimizationBarrier tlb_OptimizationBarrier_17 ( // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178778.4]
    .io_x_ppn(tlb_OptimizationBarrier_17_io_x_ppn),
    .io_x_u(tlb_OptimizationBarrier_17_io_x_u),
    .io_x_ae(tlb_OptimizationBarrier_17_io_x_ae),
    .io_x_sw(tlb_OptimizationBarrier_17_io_x_sw),
    .io_x_sx(tlb_OptimizationBarrier_17_io_x_sx),
    .io_x_sr(tlb_OptimizationBarrier_17_io_x_sr),
    .io_x_pw(tlb_OptimizationBarrier_17_io_x_pw),
    .io_x_px(tlb_OptimizationBarrier_17_io_x_px),
    .io_x_pr(tlb_OptimizationBarrier_17_io_x_pr),
    .io_x_ppp(tlb_OptimizationBarrier_17_io_x_ppp),
    .io_x_pal(tlb_OptimizationBarrier_17_io_x_pal),
    .io_x_paa(tlb_OptimizationBarrier_17_io_x_paa),
    .io_x_eff(tlb_OptimizationBarrier_17_io_x_eff),
    .io_x_c(tlb_OptimizationBarrier_17_io_x_c),
    .io_y_ppn(tlb_OptimizationBarrier_17_io_y_ppn),
    .io_y_u(tlb_OptimizationBarrier_17_io_y_u),
    .io_y_ae(tlb_OptimizationBarrier_17_io_y_ae),
    .io_y_sw(tlb_OptimizationBarrier_17_io_y_sw),
    .io_y_sx(tlb_OptimizationBarrier_17_io_y_sx),
    .io_y_sr(tlb_OptimizationBarrier_17_io_y_sr),
    .io_y_pw(tlb_OptimizationBarrier_17_io_y_pw),
    .io_y_px(tlb_OptimizationBarrier_17_io_y_px),
    .io_y_pr(tlb_OptimizationBarrier_17_io_y_pr),
    .io_y_ppp(tlb_OptimizationBarrier_17_io_y_ppp),
    .io_y_pal(tlb_OptimizationBarrier_17_io_y_pal),
    .io_y_paa(tlb_OptimizationBarrier_17_io_y_paa),
    .io_y_eff(tlb_OptimizationBarrier_17_io_y_eff),
    .io_y_c(tlb_OptimizationBarrier_17_io_y_c)
  );
  OptimizationBarrier tlb_OptimizationBarrier_18 ( // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178821.4]
    .io_x_ppn(tlb_OptimizationBarrier_18_io_x_ppn),
    .io_x_u(tlb_OptimizationBarrier_18_io_x_u),
    .io_x_ae(tlb_OptimizationBarrier_18_io_x_ae),
    .io_x_sw(tlb_OptimizationBarrier_18_io_x_sw),
    .io_x_sx(tlb_OptimizationBarrier_18_io_x_sx),
    .io_x_sr(tlb_OptimizationBarrier_18_io_x_sr),
    .io_x_pw(tlb_OptimizationBarrier_18_io_x_pw),
    .io_x_px(tlb_OptimizationBarrier_18_io_x_px),
    .io_x_pr(tlb_OptimizationBarrier_18_io_x_pr),
    .io_x_ppp(tlb_OptimizationBarrier_18_io_x_ppp),
    .io_x_pal(tlb_OptimizationBarrier_18_io_x_pal),
    .io_x_paa(tlb_OptimizationBarrier_18_io_x_paa),
    .io_x_eff(tlb_OptimizationBarrier_18_io_x_eff),
    .io_x_c(tlb_OptimizationBarrier_18_io_x_c),
    .io_y_ppn(tlb_OptimizationBarrier_18_io_y_ppn),
    .io_y_u(tlb_OptimizationBarrier_18_io_y_u),
    .io_y_ae(tlb_OptimizationBarrier_18_io_y_ae),
    .io_y_sw(tlb_OptimizationBarrier_18_io_y_sw),
    .io_y_sx(tlb_OptimizationBarrier_18_io_y_sx),
    .io_y_sr(tlb_OptimizationBarrier_18_io_y_sr),
    .io_y_pw(tlb_OptimizationBarrier_18_io_y_pw),
    .io_y_px(tlb_OptimizationBarrier_18_io_y_px),
    .io_y_pr(tlb_OptimizationBarrier_18_io_y_pr),
    .io_y_ppp(tlb_OptimizationBarrier_18_io_y_ppp),
    .io_y_pal(tlb_OptimizationBarrier_18_io_y_pal),
    .io_y_paa(tlb_OptimizationBarrier_18_io_y_paa),
    .io_y_eff(tlb_OptimizationBarrier_18_io_y_eff),
    .io_y_c(tlb_OptimizationBarrier_18_io_y_c)
  );
  OptimizationBarrier tlb_OptimizationBarrier_19 ( // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178864.4]
    .io_x_ppn(tlb_OptimizationBarrier_19_io_x_ppn),
    .io_x_u(tlb_OptimizationBarrier_19_io_x_u),
    .io_x_ae(tlb_OptimizationBarrier_19_io_x_ae),
    .io_x_sw(tlb_OptimizationBarrier_19_io_x_sw),
    .io_x_sx(tlb_OptimizationBarrier_19_io_x_sx),
    .io_x_sr(tlb_OptimizationBarrier_19_io_x_sr),
    .io_x_pw(tlb_OptimizationBarrier_19_io_x_pw),
    .io_x_px(tlb_OptimizationBarrier_19_io_x_px),
    .io_x_pr(tlb_OptimizationBarrier_19_io_x_pr),
    .io_x_ppp(tlb_OptimizationBarrier_19_io_x_ppp),
    .io_x_pal(tlb_OptimizationBarrier_19_io_x_pal),
    .io_x_paa(tlb_OptimizationBarrier_19_io_x_paa),
    .io_x_eff(tlb_OptimizationBarrier_19_io_x_eff),
    .io_x_c(tlb_OptimizationBarrier_19_io_x_c),
    .io_y_ppn(tlb_OptimizationBarrier_19_io_y_ppn),
    .io_y_u(tlb_OptimizationBarrier_19_io_y_u),
    .io_y_ae(tlb_OptimizationBarrier_19_io_y_ae),
    .io_y_sw(tlb_OptimizationBarrier_19_io_y_sw),
    .io_y_sx(tlb_OptimizationBarrier_19_io_y_sx),
    .io_y_sr(tlb_OptimizationBarrier_19_io_y_sr),
    .io_y_pw(tlb_OptimizationBarrier_19_io_y_pw),
    .io_y_px(tlb_OptimizationBarrier_19_io_y_px),
    .io_y_pr(tlb_OptimizationBarrier_19_io_y_pr),
    .io_y_ppp(tlb_OptimizationBarrier_19_io_y_ppp),
    .io_y_pal(tlb_OptimizationBarrier_19_io_y_pal),
    .io_y_paa(tlb_OptimizationBarrier_19_io_y_paa),
    .io_y_eff(tlb_OptimizationBarrier_19_io_y_eff),
    .io_y_c(tlb_OptimizationBarrier_19_io_y_c)
  );
  OptimizationBarrier tlb_OptimizationBarrier_20 ( // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178907.4]
    .io_x_ppn(tlb_OptimizationBarrier_20_io_x_ppn),
    .io_x_u(tlb_OptimizationBarrier_20_io_x_u),
    .io_x_ae(tlb_OptimizationBarrier_20_io_x_ae),
    .io_x_sw(tlb_OptimizationBarrier_20_io_x_sw),
    .io_x_sx(tlb_OptimizationBarrier_20_io_x_sx),
    .io_x_sr(tlb_OptimizationBarrier_20_io_x_sr),
    .io_x_pw(tlb_OptimizationBarrier_20_io_x_pw),
    .io_x_px(tlb_OptimizationBarrier_20_io_x_px),
    .io_x_pr(tlb_OptimizationBarrier_20_io_x_pr),
    .io_x_ppp(tlb_OptimizationBarrier_20_io_x_ppp),
    .io_x_pal(tlb_OptimizationBarrier_20_io_x_pal),
    .io_x_paa(tlb_OptimizationBarrier_20_io_x_paa),
    .io_x_eff(tlb_OptimizationBarrier_20_io_x_eff),
    .io_x_c(tlb_OptimizationBarrier_20_io_x_c),
    .io_y_ppn(tlb_OptimizationBarrier_20_io_y_ppn),
    .io_y_u(tlb_OptimizationBarrier_20_io_y_u),
    .io_y_ae(tlb_OptimizationBarrier_20_io_y_ae),
    .io_y_sw(tlb_OptimizationBarrier_20_io_y_sw),
    .io_y_sx(tlb_OptimizationBarrier_20_io_y_sx),
    .io_y_sr(tlb_OptimizationBarrier_20_io_y_sr),
    .io_y_pw(tlb_OptimizationBarrier_20_io_y_pw),
    .io_y_px(tlb_OptimizationBarrier_20_io_y_px),
    .io_y_pr(tlb_OptimizationBarrier_20_io_y_pr),
    .io_y_ppp(tlb_OptimizationBarrier_20_io_y_ppp),
    .io_y_pal(tlb_OptimizationBarrier_20_io_y_pal),
    .io_y_paa(tlb_OptimizationBarrier_20_io_y_paa),
    .io_y_eff(tlb_OptimizationBarrier_20_io_y_eff),
    .io_y_c(tlb_OptimizationBarrier_20_io_y_c)
  );
  OptimizationBarrier tlb_OptimizationBarrier_21 ( // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178950.4]
    .io_x_ppn(tlb_OptimizationBarrier_21_io_x_ppn),
    .io_x_u(tlb_OptimizationBarrier_21_io_x_u),
    .io_x_ae(tlb_OptimizationBarrier_21_io_x_ae),
    .io_x_sw(tlb_OptimizationBarrier_21_io_x_sw),
    .io_x_sx(tlb_OptimizationBarrier_21_io_x_sx),
    .io_x_sr(tlb_OptimizationBarrier_21_io_x_sr),
    .io_x_pw(tlb_OptimizationBarrier_21_io_x_pw),
    .io_x_px(tlb_OptimizationBarrier_21_io_x_px),
    .io_x_pr(tlb_OptimizationBarrier_21_io_x_pr),
    .io_x_ppp(tlb_OptimizationBarrier_21_io_x_ppp),
    .io_x_pal(tlb_OptimizationBarrier_21_io_x_pal),
    .io_x_paa(tlb_OptimizationBarrier_21_io_x_paa),
    .io_x_eff(tlb_OptimizationBarrier_21_io_x_eff),
    .io_x_c(tlb_OptimizationBarrier_21_io_x_c),
    .io_y_ppn(tlb_OptimizationBarrier_21_io_y_ppn),
    .io_y_u(tlb_OptimizationBarrier_21_io_y_u),
    .io_y_ae(tlb_OptimizationBarrier_21_io_y_ae),
    .io_y_sw(tlb_OptimizationBarrier_21_io_y_sw),
    .io_y_sx(tlb_OptimizationBarrier_21_io_y_sx),
    .io_y_sr(tlb_OptimizationBarrier_21_io_y_sr),
    .io_y_pw(tlb_OptimizationBarrier_21_io_y_pw),
    .io_y_px(tlb_OptimizationBarrier_21_io_y_px),
    .io_y_pr(tlb_OptimizationBarrier_21_io_y_pr),
    .io_y_ppp(tlb_OptimizationBarrier_21_io_y_ppp),
    .io_y_pal(tlb_OptimizationBarrier_21_io_y_pal),
    .io_y_paa(tlb_OptimizationBarrier_21_io_y_paa),
    .io_y_eff(tlb_OptimizationBarrier_21_io_y_eff),
    .io_y_c(tlb_OptimizationBarrier_21_io_y_c)
  );
  OptimizationBarrier tlb_OptimizationBarrier_22 ( // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178992.4]
    .io_x_ppn(tlb_OptimizationBarrier_22_io_x_ppn),
    .io_x_u(tlb_OptimizationBarrier_22_io_x_u),
    .io_x_ae(tlb_OptimizationBarrier_22_io_x_ae),
    .io_x_sw(tlb_OptimizationBarrier_22_io_x_sw),
    .io_x_sx(tlb_OptimizationBarrier_22_io_x_sx),
    .io_x_sr(tlb_OptimizationBarrier_22_io_x_sr),
    .io_x_pw(tlb_OptimizationBarrier_22_io_x_pw),
    .io_x_px(tlb_OptimizationBarrier_22_io_x_px),
    .io_x_pr(tlb_OptimizationBarrier_22_io_x_pr),
    .io_x_ppp(tlb_OptimizationBarrier_22_io_x_ppp),
    .io_x_pal(tlb_OptimizationBarrier_22_io_x_pal),
    .io_x_paa(tlb_OptimizationBarrier_22_io_x_paa),
    .io_x_eff(tlb_OptimizationBarrier_22_io_x_eff),
    .io_x_c(tlb_OptimizationBarrier_22_io_x_c),
    .io_y_ppn(tlb_OptimizationBarrier_22_io_y_ppn),
    .io_y_u(tlb_OptimizationBarrier_22_io_y_u),
    .io_y_ae(tlb_OptimizationBarrier_22_io_y_ae),
    .io_y_sw(tlb_OptimizationBarrier_22_io_y_sw),
    .io_y_sx(tlb_OptimizationBarrier_22_io_y_sx),
    .io_y_sr(tlb_OptimizationBarrier_22_io_y_sr),
    .io_y_pw(tlb_OptimizationBarrier_22_io_y_pw),
    .io_y_px(tlb_OptimizationBarrier_22_io_y_px),
    .io_y_pr(tlb_OptimizationBarrier_22_io_y_pr),
    .io_y_ppp(tlb_OptimizationBarrier_22_io_y_ppp),
    .io_y_pal(tlb_OptimizationBarrier_22_io_y_pal),
    .io_y_paa(tlb_OptimizationBarrier_22_io_y_paa),
    .io_y_eff(tlb_OptimizationBarrier_22_io_y_eff),
    .io_y_c(tlb_OptimizationBarrier_22_io_y_c)
  );
  OptimizationBarrier tlb_OptimizationBarrier_23 ( // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179034.4]
    .io_x_ppn(tlb_OptimizationBarrier_23_io_x_ppn),
    .io_x_u(tlb_OptimizationBarrier_23_io_x_u),
    .io_x_ae(tlb_OptimizationBarrier_23_io_x_ae),
    .io_x_sw(tlb_OptimizationBarrier_23_io_x_sw),
    .io_x_sx(tlb_OptimizationBarrier_23_io_x_sx),
    .io_x_sr(tlb_OptimizationBarrier_23_io_x_sr),
    .io_x_pw(tlb_OptimizationBarrier_23_io_x_pw),
    .io_x_px(tlb_OptimizationBarrier_23_io_x_px),
    .io_x_pr(tlb_OptimizationBarrier_23_io_x_pr),
    .io_x_ppp(tlb_OptimizationBarrier_23_io_x_ppp),
    .io_x_pal(tlb_OptimizationBarrier_23_io_x_pal),
    .io_x_paa(tlb_OptimizationBarrier_23_io_x_paa),
    .io_x_eff(tlb_OptimizationBarrier_23_io_x_eff),
    .io_x_c(tlb_OptimizationBarrier_23_io_x_c),
    .io_y_ppn(tlb_OptimizationBarrier_23_io_y_ppn),
    .io_y_u(tlb_OptimizationBarrier_23_io_y_u),
    .io_y_ae(tlb_OptimizationBarrier_23_io_y_ae),
    .io_y_sw(tlb_OptimizationBarrier_23_io_y_sw),
    .io_y_sx(tlb_OptimizationBarrier_23_io_y_sx),
    .io_y_sr(tlb_OptimizationBarrier_23_io_y_sr),
    .io_y_pw(tlb_OptimizationBarrier_23_io_y_pw),
    .io_y_px(tlb_OptimizationBarrier_23_io_y_px),
    .io_y_pr(tlb_OptimizationBarrier_23_io_y_pr),
    .io_y_ppp(tlb_OptimizationBarrier_23_io_y_ppp),
    .io_y_pal(tlb_OptimizationBarrier_23_io_y_pal),
    .io_y_paa(tlb_OptimizationBarrier_23_io_y_paa),
    .io_y_eff(tlb_OptimizationBarrier_23_io_y_eff),
    .io_y_c(tlb_OptimizationBarrier_23_io_y_c)
  );
  OptimizationBarrier tlb_OptimizationBarrier_24 ( // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179076.4]
    .io_x_ppn(tlb_OptimizationBarrier_24_io_x_ppn),
    .io_x_u(tlb_OptimizationBarrier_24_io_x_u),
    .io_x_ae(tlb_OptimizationBarrier_24_io_x_ae),
    .io_x_sw(tlb_OptimizationBarrier_24_io_x_sw),
    .io_x_sx(tlb_OptimizationBarrier_24_io_x_sx),
    .io_x_sr(tlb_OptimizationBarrier_24_io_x_sr),
    .io_x_pw(tlb_OptimizationBarrier_24_io_x_pw),
    .io_x_px(tlb_OptimizationBarrier_24_io_x_px),
    .io_x_pr(tlb_OptimizationBarrier_24_io_x_pr),
    .io_x_ppp(tlb_OptimizationBarrier_24_io_x_ppp),
    .io_x_pal(tlb_OptimizationBarrier_24_io_x_pal),
    .io_x_paa(tlb_OptimizationBarrier_24_io_x_paa),
    .io_x_eff(tlb_OptimizationBarrier_24_io_x_eff),
    .io_x_c(tlb_OptimizationBarrier_24_io_x_c),
    .io_y_ppn(tlb_OptimizationBarrier_24_io_y_ppn),
    .io_y_u(tlb_OptimizationBarrier_24_io_y_u),
    .io_y_ae(tlb_OptimizationBarrier_24_io_y_ae),
    .io_y_sw(tlb_OptimizationBarrier_24_io_y_sw),
    .io_y_sx(tlb_OptimizationBarrier_24_io_y_sx),
    .io_y_sr(tlb_OptimizationBarrier_24_io_y_sr),
    .io_y_pw(tlb_OptimizationBarrier_24_io_y_pw),
    .io_y_px(tlb_OptimizationBarrier_24_io_y_px),
    .io_y_pr(tlb_OptimizationBarrier_24_io_y_pr),
    .io_y_ppp(tlb_OptimizationBarrier_24_io_y_ppp),
    .io_y_pal(tlb_OptimizationBarrier_24_io_y_pal),
    .io_y_paa(tlb_OptimizationBarrier_24_io_y_paa),
    .io_y_eff(tlb_OptimizationBarrier_24_io_y_eff),
    .io_y_c(tlb_OptimizationBarrier_24_io_y_c)
  );
  OptimizationBarrier tlb_OptimizationBarrier_25 ( // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179118.4]
    .io_x_ppn(tlb_OptimizationBarrier_25_io_x_ppn),
    .io_x_u(tlb_OptimizationBarrier_25_io_x_u),
    .io_x_ae(tlb_OptimizationBarrier_25_io_x_ae),
    .io_x_sw(tlb_OptimizationBarrier_25_io_x_sw),
    .io_x_sx(tlb_OptimizationBarrier_25_io_x_sx),
    .io_x_sr(tlb_OptimizationBarrier_25_io_x_sr),
    .io_x_pw(tlb_OptimizationBarrier_25_io_x_pw),
    .io_x_px(tlb_OptimizationBarrier_25_io_x_px),
    .io_x_pr(tlb_OptimizationBarrier_25_io_x_pr),
    .io_x_ppp(tlb_OptimizationBarrier_25_io_x_ppp),
    .io_x_pal(tlb_OptimizationBarrier_25_io_x_pal),
    .io_x_paa(tlb_OptimizationBarrier_25_io_x_paa),
    .io_x_eff(tlb_OptimizationBarrier_25_io_x_eff),
    .io_x_c(tlb_OptimizationBarrier_25_io_x_c),
    .io_y_ppn(tlb_OptimizationBarrier_25_io_y_ppn),
    .io_y_u(tlb_OptimizationBarrier_25_io_y_u),
    .io_y_ae(tlb_OptimizationBarrier_25_io_y_ae),
    .io_y_sw(tlb_OptimizationBarrier_25_io_y_sw),
    .io_y_sx(tlb_OptimizationBarrier_25_io_y_sx),
    .io_y_sr(tlb_OptimizationBarrier_25_io_y_sr),
    .io_y_pw(tlb_OptimizationBarrier_25_io_y_pw),
    .io_y_px(tlb_OptimizationBarrier_25_io_y_px),
    .io_y_pr(tlb_OptimizationBarrier_25_io_y_pr),
    .io_y_ppp(tlb_OptimizationBarrier_25_io_y_ppp),
    .io_y_pal(tlb_OptimizationBarrier_25_io_y_pal),
    .io_y_paa(tlb_OptimizationBarrier_25_io_y_paa),
    .io_y_eff(tlb_OptimizationBarrier_25_io_y_eff),
    .io_y_c(tlb_OptimizationBarrier_25_io_y_c)
  );
  OptimizationBarrier tlb_OptimizationBarrier_26 ( // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179160.4]
    .io_x_ppn(tlb_OptimizationBarrier_26_io_x_ppn),
    .io_x_u(tlb_OptimizationBarrier_26_io_x_u),
    .io_x_ae(tlb_OptimizationBarrier_26_io_x_ae),
    .io_x_sw(tlb_OptimizationBarrier_26_io_x_sw),
    .io_x_sx(tlb_OptimizationBarrier_26_io_x_sx),
    .io_x_sr(tlb_OptimizationBarrier_26_io_x_sr),
    .io_x_pw(tlb_OptimizationBarrier_26_io_x_pw),
    .io_x_px(tlb_OptimizationBarrier_26_io_x_px),
    .io_x_pr(tlb_OptimizationBarrier_26_io_x_pr),
    .io_x_ppp(tlb_OptimizationBarrier_26_io_x_ppp),
    .io_x_pal(tlb_OptimizationBarrier_26_io_x_pal),
    .io_x_paa(tlb_OptimizationBarrier_26_io_x_paa),
    .io_x_eff(tlb_OptimizationBarrier_26_io_x_eff),
    .io_x_c(tlb_OptimizationBarrier_26_io_x_c),
    .io_y_ppn(tlb_OptimizationBarrier_26_io_y_ppn),
    .io_y_u(tlb_OptimizationBarrier_26_io_y_u),
    .io_y_ae(tlb_OptimizationBarrier_26_io_y_ae),
    .io_y_sw(tlb_OptimizationBarrier_26_io_y_sw),
    .io_y_sx(tlb_OptimizationBarrier_26_io_y_sx),
    .io_y_sr(tlb_OptimizationBarrier_26_io_y_sr),
    .io_y_pw(tlb_OptimizationBarrier_26_io_y_pw),
    .io_y_px(tlb_OptimizationBarrier_26_io_y_px),
    .io_y_pr(tlb_OptimizationBarrier_26_io_y_pr),
    .io_y_ppp(tlb_OptimizationBarrier_26_io_y_ppp),
    .io_y_pal(tlb_OptimizationBarrier_26_io_y_pal),
    .io_y_paa(tlb_OptimizationBarrier_26_io_y_paa),
    .io_y_eff(tlb_OptimizationBarrier_26_io_y_eff),
    .io_y_c(tlb_OptimizationBarrier_26_io_y_c)
  );
  OptimizationBarrier tlb_OptimizationBarrier_27 ( // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179203.4]
    .io_x_ppn(tlb_OptimizationBarrier_27_io_x_ppn),
    .io_x_u(tlb_OptimizationBarrier_27_io_x_u),
    .io_x_ae(tlb_OptimizationBarrier_27_io_x_ae),
    .io_x_sw(tlb_OptimizationBarrier_27_io_x_sw),
    .io_x_sx(tlb_OptimizationBarrier_27_io_x_sx),
    .io_x_sr(tlb_OptimizationBarrier_27_io_x_sr),
    .io_x_pw(tlb_OptimizationBarrier_27_io_x_pw),
    .io_x_px(tlb_OptimizationBarrier_27_io_x_px),
    .io_x_pr(tlb_OptimizationBarrier_27_io_x_pr),
    .io_x_ppp(tlb_OptimizationBarrier_27_io_x_ppp),
    .io_x_pal(tlb_OptimizationBarrier_27_io_x_pal),
    .io_x_paa(tlb_OptimizationBarrier_27_io_x_paa),
    .io_x_eff(tlb_OptimizationBarrier_27_io_x_eff),
    .io_x_c(tlb_OptimizationBarrier_27_io_x_c),
    .io_y_ppn(tlb_OptimizationBarrier_27_io_y_ppn),
    .io_y_u(tlb_OptimizationBarrier_27_io_y_u),
    .io_y_ae(tlb_OptimizationBarrier_27_io_y_ae),
    .io_y_sw(tlb_OptimizationBarrier_27_io_y_sw),
    .io_y_sx(tlb_OptimizationBarrier_27_io_y_sx),
    .io_y_sr(tlb_OptimizationBarrier_27_io_y_sr),
    .io_y_pw(tlb_OptimizationBarrier_27_io_y_pw),
    .io_y_px(tlb_OptimizationBarrier_27_io_y_px),
    .io_y_pr(tlb_OptimizationBarrier_27_io_y_pr),
    .io_y_ppp(tlb_OptimizationBarrier_27_io_y_ppp),
    .io_y_pal(tlb_OptimizationBarrier_27_io_y_pal),
    .io_y_paa(tlb_OptimizationBarrier_27_io_y_paa),
    .io_y_eff(tlb_OptimizationBarrier_27_io_y_eff),
    .io_y_c(tlb_OptimizationBarrier_27_io_y_c)
  );
  OptimizationBarrier tlb_OptimizationBarrier_28 ( // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179246.4]
    .io_x_ppn(tlb_OptimizationBarrier_28_io_x_ppn),
    .io_x_u(tlb_OptimizationBarrier_28_io_x_u),
    .io_x_ae(tlb_OptimizationBarrier_28_io_x_ae),
    .io_x_sw(tlb_OptimizationBarrier_28_io_x_sw),
    .io_x_sx(tlb_OptimizationBarrier_28_io_x_sx),
    .io_x_sr(tlb_OptimizationBarrier_28_io_x_sr),
    .io_x_pw(tlb_OptimizationBarrier_28_io_x_pw),
    .io_x_px(tlb_OptimizationBarrier_28_io_x_px),
    .io_x_pr(tlb_OptimizationBarrier_28_io_x_pr),
    .io_x_ppp(tlb_OptimizationBarrier_28_io_x_ppp),
    .io_x_pal(tlb_OptimizationBarrier_28_io_x_pal),
    .io_x_paa(tlb_OptimizationBarrier_28_io_x_paa),
    .io_x_eff(tlb_OptimizationBarrier_28_io_x_eff),
    .io_x_c(tlb_OptimizationBarrier_28_io_x_c),
    .io_y_ppn(tlb_OptimizationBarrier_28_io_y_ppn),
    .io_y_u(tlb_OptimizationBarrier_28_io_y_u),
    .io_y_ae(tlb_OptimizationBarrier_28_io_y_ae),
    .io_y_sw(tlb_OptimizationBarrier_28_io_y_sw),
    .io_y_sx(tlb_OptimizationBarrier_28_io_y_sx),
    .io_y_sr(tlb_OptimizationBarrier_28_io_y_sr),
    .io_y_pw(tlb_OptimizationBarrier_28_io_y_pw),
    .io_y_px(tlb_OptimizationBarrier_28_io_y_px),
    .io_y_pr(tlb_OptimizationBarrier_28_io_y_pr),
    .io_y_ppp(tlb_OptimizationBarrier_28_io_y_ppp),
    .io_y_pal(tlb_OptimizationBarrier_28_io_y_pal),
    .io_y_paa(tlb_OptimizationBarrier_28_io_y_paa),
    .io_y_eff(tlb_OptimizationBarrier_28_io_y_eff),
    .io_y_c(tlb_OptimizationBarrier_28_io_y_c)
  );
  OptimizationBarrier tlb_OptimizationBarrier_29 ( // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179289.4]
    .io_x_ppn(tlb_OptimizationBarrier_29_io_x_ppn),
    .io_x_u(tlb_OptimizationBarrier_29_io_x_u),
    .io_x_ae(tlb_OptimizationBarrier_29_io_x_ae),
    .io_x_sw(tlb_OptimizationBarrier_29_io_x_sw),
    .io_x_sx(tlb_OptimizationBarrier_29_io_x_sx),
    .io_x_sr(tlb_OptimizationBarrier_29_io_x_sr),
    .io_x_pw(tlb_OptimizationBarrier_29_io_x_pw),
    .io_x_px(tlb_OptimizationBarrier_29_io_x_px),
    .io_x_pr(tlb_OptimizationBarrier_29_io_x_pr),
    .io_x_ppp(tlb_OptimizationBarrier_29_io_x_ppp),
    .io_x_pal(tlb_OptimizationBarrier_29_io_x_pal),
    .io_x_paa(tlb_OptimizationBarrier_29_io_x_paa),
    .io_x_eff(tlb_OptimizationBarrier_29_io_x_eff),
    .io_x_c(tlb_OptimizationBarrier_29_io_x_c),
    .io_y_ppn(tlb_OptimizationBarrier_29_io_y_ppn),
    .io_y_u(tlb_OptimizationBarrier_29_io_y_u),
    .io_y_ae(tlb_OptimizationBarrier_29_io_y_ae),
    .io_y_sw(tlb_OptimizationBarrier_29_io_y_sw),
    .io_y_sx(tlb_OptimizationBarrier_29_io_y_sx),
    .io_y_sr(tlb_OptimizationBarrier_29_io_y_sr),
    .io_y_pw(tlb_OptimizationBarrier_29_io_y_pw),
    .io_y_px(tlb_OptimizationBarrier_29_io_y_px),
    .io_y_pr(tlb_OptimizationBarrier_29_io_y_pr),
    .io_y_ppp(tlb_OptimizationBarrier_29_io_y_ppp),
    .io_y_pal(tlb_OptimizationBarrier_29_io_y_pal),
    .io_y_paa(tlb_OptimizationBarrier_29_io_y_paa),
    .io_y_eff(tlb_OptimizationBarrier_29_io_y_eff),
    .io_y_c(tlb_OptimizationBarrier_29_io_y_c)
  );
  OptimizationBarrier tlb_OptimizationBarrier_30 ( // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179332.4]
    .io_x_ppn(tlb_OptimizationBarrier_30_io_x_ppn),
    .io_x_u(tlb_OptimizationBarrier_30_io_x_u),
    .io_x_ae(tlb_OptimizationBarrier_30_io_x_ae),
    .io_x_sw(tlb_OptimizationBarrier_30_io_x_sw),
    .io_x_sx(tlb_OptimizationBarrier_30_io_x_sx),
    .io_x_sr(tlb_OptimizationBarrier_30_io_x_sr),
    .io_x_pw(tlb_OptimizationBarrier_30_io_x_pw),
    .io_x_px(tlb_OptimizationBarrier_30_io_x_px),
    .io_x_pr(tlb_OptimizationBarrier_30_io_x_pr),
    .io_x_ppp(tlb_OptimizationBarrier_30_io_x_ppp),
    .io_x_pal(tlb_OptimizationBarrier_30_io_x_pal),
    .io_x_paa(tlb_OptimizationBarrier_30_io_x_paa),
    .io_x_eff(tlb_OptimizationBarrier_30_io_x_eff),
    .io_x_c(tlb_OptimizationBarrier_30_io_x_c),
    .io_y_ppn(tlb_OptimizationBarrier_30_io_y_ppn),
    .io_y_u(tlb_OptimizationBarrier_30_io_y_u),
    .io_y_ae(tlb_OptimizationBarrier_30_io_y_ae),
    .io_y_sw(tlb_OptimizationBarrier_30_io_y_sw),
    .io_y_sx(tlb_OptimizationBarrier_30_io_y_sx),
    .io_y_sr(tlb_OptimizationBarrier_30_io_y_sr),
    .io_y_pw(tlb_OptimizationBarrier_30_io_y_pw),
    .io_y_px(tlb_OptimizationBarrier_30_io_y_px),
    .io_y_pr(tlb_OptimizationBarrier_30_io_y_pr),
    .io_y_ppp(tlb_OptimizationBarrier_30_io_y_ppp),
    .io_y_pal(tlb_OptimizationBarrier_30_io_y_pal),
    .io_y_paa(tlb_OptimizationBarrier_30_io_y_paa),
    .io_y_eff(tlb_OptimizationBarrier_30_io_y_eff),
    .io_y_c(tlb_OptimizationBarrier_30_io_y_c)
  );
  OptimizationBarrier tlb_OptimizationBarrier_31 ( // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179375.4]
    .io_x_ppn(tlb_OptimizationBarrier_31_io_x_ppn),
    .io_x_u(tlb_OptimizationBarrier_31_io_x_u),
    .io_x_ae(tlb_OptimizationBarrier_31_io_x_ae),
    .io_x_sw(tlb_OptimizationBarrier_31_io_x_sw),
    .io_x_sx(tlb_OptimizationBarrier_31_io_x_sx),
    .io_x_sr(tlb_OptimizationBarrier_31_io_x_sr),
    .io_x_pw(tlb_OptimizationBarrier_31_io_x_pw),
    .io_x_px(tlb_OptimizationBarrier_31_io_x_px),
    .io_x_pr(tlb_OptimizationBarrier_31_io_x_pr),
    .io_x_ppp(tlb_OptimizationBarrier_31_io_x_ppp),
    .io_x_pal(tlb_OptimizationBarrier_31_io_x_pal),
    .io_x_paa(tlb_OptimizationBarrier_31_io_x_paa),
    .io_x_eff(tlb_OptimizationBarrier_31_io_x_eff),
    .io_x_c(tlb_OptimizationBarrier_31_io_x_c),
    .io_y_ppn(tlb_OptimizationBarrier_31_io_y_ppn),
    .io_y_u(tlb_OptimizationBarrier_31_io_y_u),
    .io_y_ae(tlb_OptimizationBarrier_31_io_y_ae),
    .io_y_sw(tlb_OptimizationBarrier_31_io_y_sw),
    .io_y_sx(tlb_OptimizationBarrier_31_io_y_sx),
    .io_y_sr(tlb_OptimizationBarrier_31_io_y_sr),
    .io_y_pw(tlb_OptimizationBarrier_31_io_y_pw),
    .io_y_px(tlb_OptimizationBarrier_31_io_y_px),
    .io_y_pr(tlb_OptimizationBarrier_31_io_y_pr),
    .io_y_ppp(tlb_OptimizationBarrier_31_io_y_ppp),
    .io_y_pal(tlb_OptimizationBarrier_31_io_y_pal),
    .io_y_paa(tlb_OptimizationBarrier_31_io_y_paa),
    .io_y_eff(tlb_OptimizationBarrier_31_io_y_eff),
    .io_y_c(tlb_OptimizationBarrier_31_io_y_c)
  );
  OptimizationBarrier tlb_OptimizationBarrier_32 ( // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179418.4]
    .io_x_ppn(tlb_OptimizationBarrier_32_io_x_ppn),
    .io_x_u(tlb_OptimizationBarrier_32_io_x_u),
    .io_x_ae(tlb_OptimizationBarrier_32_io_x_ae),
    .io_x_sw(tlb_OptimizationBarrier_32_io_x_sw),
    .io_x_sx(tlb_OptimizationBarrier_32_io_x_sx),
    .io_x_sr(tlb_OptimizationBarrier_32_io_x_sr),
    .io_x_pw(tlb_OptimizationBarrier_32_io_x_pw),
    .io_x_px(tlb_OptimizationBarrier_32_io_x_px),
    .io_x_pr(tlb_OptimizationBarrier_32_io_x_pr),
    .io_x_ppp(tlb_OptimizationBarrier_32_io_x_ppp),
    .io_x_pal(tlb_OptimizationBarrier_32_io_x_pal),
    .io_x_paa(tlb_OptimizationBarrier_32_io_x_paa),
    .io_x_eff(tlb_OptimizationBarrier_32_io_x_eff),
    .io_x_c(tlb_OptimizationBarrier_32_io_x_c),
    .io_y_ppn(tlb_OptimizationBarrier_32_io_y_ppn),
    .io_y_u(tlb_OptimizationBarrier_32_io_y_u),
    .io_y_ae(tlb_OptimizationBarrier_32_io_y_ae),
    .io_y_sw(tlb_OptimizationBarrier_32_io_y_sw),
    .io_y_sx(tlb_OptimizationBarrier_32_io_y_sx),
    .io_y_sr(tlb_OptimizationBarrier_32_io_y_sr),
    .io_y_pw(tlb_OptimizationBarrier_32_io_y_pw),
    .io_y_px(tlb_OptimizationBarrier_32_io_y_px),
    .io_y_pr(tlb_OptimizationBarrier_32_io_y_pr),
    .io_y_ppp(tlb_OptimizationBarrier_32_io_y_ppp),
    .io_y_pal(tlb_OptimizationBarrier_32_io_y_pal),
    .io_y_paa(tlb_OptimizationBarrier_32_io_y_paa),
    .io_y_eff(tlb_OptimizationBarrier_32_io_y_eff),
    .io_y_c(tlb_OptimizationBarrier_32_io_y_c)
  );
  OptimizationBarrier tlb_OptimizationBarrier_33 ( // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179461.4]
    .io_x_ppn(tlb_OptimizationBarrier_33_io_x_ppn),
    .io_x_u(tlb_OptimizationBarrier_33_io_x_u),
    .io_x_ae(tlb_OptimizationBarrier_33_io_x_ae),
    .io_x_sw(tlb_OptimizationBarrier_33_io_x_sw),
    .io_x_sx(tlb_OptimizationBarrier_33_io_x_sx),
    .io_x_sr(tlb_OptimizationBarrier_33_io_x_sr),
    .io_x_pw(tlb_OptimizationBarrier_33_io_x_pw),
    .io_x_px(tlb_OptimizationBarrier_33_io_x_px),
    .io_x_pr(tlb_OptimizationBarrier_33_io_x_pr),
    .io_x_ppp(tlb_OptimizationBarrier_33_io_x_ppp),
    .io_x_pal(tlb_OptimizationBarrier_33_io_x_pal),
    .io_x_paa(tlb_OptimizationBarrier_33_io_x_paa),
    .io_x_eff(tlb_OptimizationBarrier_33_io_x_eff),
    .io_x_c(tlb_OptimizationBarrier_33_io_x_c),
    .io_y_ppn(tlb_OptimizationBarrier_33_io_y_ppn),
    .io_y_u(tlb_OptimizationBarrier_33_io_y_u),
    .io_y_ae(tlb_OptimizationBarrier_33_io_y_ae),
    .io_y_sw(tlb_OptimizationBarrier_33_io_y_sw),
    .io_y_sx(tlb_OptimizationBarrier_33_io_y_sx),
    .io_y_sr(tlb_OptimizationBarrier_33_io_y_sr),
    .io_y_pw(tlb_OptimizationBarrier_33_io_y_pw),
    .io_y_px(tlb_OptimizationBarrier_33_io_y_px),
    .io_y_pr(tlb_OptimizationBarrier_33_io_y_pr),
    .io_y_ppp(tlb_OptimizationBarrier_33_io_y_ppp),
    .io_y_pal(tlb_OptimizationBarrier_33_io_y_pal),
    .io_y_paa(tlb_OptimizationBarrier_33_io_y_paa),
    .io_y_eff(tlb_OptimizationBarrier_33_io_y_eff),
    .io_y_c(tlb_OptimizationBarrier_33_io_y_c)
  );
  OptimizationBarrier tlb_OptimizationBarrier_34 ( // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179504.4]
    .io_x_ppn(tlb_OptimizationBarrier_34_io_x_ppn),
    .io_x_u(tlb_OptimizationBarrier_34_io_x_u),
    .io_x_ae(tlb_OptimizationBarrier_34_io_x_ae),
    .io_x_sw(tlb_OptimizationBarrier_34_io_x_sw),
    .io_x_sx(tlb_OptimizationBarrier_34_io_x_sx),
    .io_x_sr(tlb_OptimizationBarrier_34_io_x_sr),
    .io_x_pw(tlb_OptimizationBarrier_34_io_x_pw),
    .io_x_px(tlb_OptimizationBarrier_34_io_x_px),
    .io_x_pr(tlb_OptimizationBarrier_34_io_x_pr),
    .io_x_ppp(tlb_OptimizationBarrier_34_io_x_ppp),
    .io_x_pal(tlb_OptimizationBarrier_34_io_x_pal),
    .io_x_paa(tlb_OptimizationBarrier_34_io_x_paa),
    .io_x_eff(tlb_OptimizationBarrier_34_io_x_eff),
    .io_x_c(tlb_OptimizationBarrier_34_io_x_c),
    .io_y_ppn(tlb_OptimizationBarrier_34_io_y_ppn),
    .io_y_u(tlb_OptimizationBarrier_34_io_y_u),
    .io_y_ae(tlb_OptimizationBarrier_34_io_y_ae),
    .io_y_sw(tlb_OptimizationBarrier_34_io_y_sw),
    .io_y_sx(tlb_OptimizationBarrier_34_io_y_sx),
    .io_y_sr(tlb_OptimizationBarrier_34_io_y_sr),
    .io_y_pw(tlb_OptimizationBarrier_34_io_y_pw),
    .io_y_px(tlb_OptimizationBarrier_34_io_y_px),
    .io_y_pr(tlb_OptimizationBarrier_34_io_y_pr),
    .io_y_ppp(tlb_OptimizationBarrier_34_io_y_ppp),
    .io_y_pal(tlb_OptimizationBarrier_34_io_y_pal),
    .io_y_paa(tlb_OptimizationBarrier_34_io_y_paa),
    .io_y_eff(tlb_OptimizationBarrier_34_io_y_eff),
    .io_y_c(tlb_OptimizationBarrier_34_io_y_c)
  );
  OptimizationBarrier tlb_OptimizationBarrier_35 ( // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179546.4]
    .io_x_ppn(tlb_OptimizationBarrier_35_io_x_ppn),
    .io_x_u(tlb_OptimizationBarrier_35_io_x_u),
    .io_x_ae(tlb_OptimizationBarrier_35_io_x_ae),
    .io_x_sw(tlb_OptimizationBarrier_35_io_x_sw),
    .io_x_sx(tlb_OptimizationBarrier_35_io_x_sx),
    .io_x_sr(tlb_OptimizationBarrier_35_io_x_sr),
    .io_x_pw(tlb_OptimizationBarrier_35_io_x_pw),
    .io_x_px(tlb_OptimizationBarrier_35_io_x_px),
    .io_x_pr(tlb_OptimizationBarrier_35_io_x_pr),
    .io_x_ppp(tlb_OptimizationBarrier_35_io_x_ppp),
    .io_x_pal(tlb_OptimizationBarrier_35_io_x_pal),
    .io_x_paa(tlb_OptimizationBarrier_35_io_x_paa),
    .io_x_eff(tlb_OptimizationBarrier_35_io_x_eff),
    .io_x_c(tlb_OptimizationBarrier_35_io_x_c),
    .io_y_ppn(tlb_OptimizationBarrier_35_io_y_ppn),
    .io_y_u(tlb_OptimizationBarrier_35_io_y_u),
    .io_y_ae(tlb_OptimizationBarrier_35_io_y_ae),
    .io_y_sw(tlb_OptimizationBarrier_35_io_y_sw),
    .io_y_sx(tlb_OptimizationBarrier_35_io_y_sx),
    .io_y_sr(tlb_OptimizationBarrier_35_io_y_sr),
    .io_y_pw(tlb_OptimizationBarrier_35_io_y_pw),
    .io_y_px(tlb_OptimizationBarrier_35_io_y_px),
    .io_y_pr(tlb_OptimizationBarrier_35_io_y_pr),
    .io_y_ppp(tlb_OptimizationBarrier_35_io_y_ppp),
    .io_y_pal(tlb_OptimizationBarrier_35_io_y_pal),
    .io_y_paa(tlb_OptimizationBarrier_35_io_y_paa),
    .io_y_eff(tlb_OptimizationBarrier_35_io_y_eff),
    .io_y_c(tlb_OptimizationBarrier_35_io_y_c)
  );
  OptimizationBarrier tlb_OptimizationBarrier_36 ( // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179588.4]
    .io_x_ppn(tlb_OptimizationBarrier_36_io_x_ppn),
    .io_x_u(tlb_OptimizationBarrier_36_io_x_u),
    .io_x_ae(tlb_OptimizationBarrier_36_io_x_ae),
    .io_x_sw(tlb_OptimizationBarrier_36_io_x_sw),
    .io_x_sx(tlb_OptimizationBarrier_36_io_x_sx),
    .io_x_sr(tlb_OptimizationBarrier_36_io_x_sr),
    .io_x_pw(tlb_OptimizationBarrier_36_io_x_pw),
    .io_x_px(tlb_OptimizationBarrier_36_io_x_px),
    .io_x_pr(tlb_OptimizationBarrier_36_io_x_pr),
    .io_x_ppp(tlb_OptimizationBarrier_36_io_x_ppp),
    .io_x_pal(tlb_OptimizationBarrier_36_io_x_pal),
    .io_x_paa(tlb_OptimizationBarrier_36_io_x_paa),
    .io_x_eff(tlb_OptimizationBarrier_36_io_x_eff),
    .io_x_c(tlb_OptimizationBarrier_36_io_x_c),
    .io_y_ppn(tlb_OptimizationBarrier_36_io_y_ppn),
    .io_y_u(tlb_OptimizationBarrier_36_io_y_u),
    .io_y_ae(tlb_OptimizationBarrier_36_io_y_ae),
    .io_y_sw(tlb_OptimizationBarrier_36_io_y_sw),
    .io_y_sx(tlb_OptimizationBarrier_36_io_y_sx),
    .io_y_sr(tlb_OptimizationBarrier_36_io_y_sr),
    .io_y_pw(tlb_OptimizationBarrier_36_io_y_pw),
    .io_y_px(tlb_OptimizationBarrier_36_io_y_px),
    .io_y_pr(tlb_OptimizationBarrier_36_io_y_pr),
    .io_y_ppp(tlb_OptimizationBarrier_36_io_y_ppp),
    .io_y_pal(tlb_OptimizationBarrier_36_io_y_pal),
    .io_y_paa(tlb_OptimizationBarrier_36_io_y_paa),
    .io_y_eff(tlb_OptimizationBarrier_36_io_y_eff),
    .io_y_c(tlb_OptimizationBarrier_36_io_y_c)
  );
  OptimizationBarrier tlb_OptimizationBarrier_37 ( // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179630.4]
    .io_x_ppn(tlb_OptimizationBarrier_37_io_x_ppn),
    .io_x_u(tlb_OptimizationBarrier_37_io_x_u),
    .io_x_ae(tlb_OptimizationBarrier_37_io_x_ae),
    .io_x_sw(tlb_OptimizationBarrier_37_io_x_sw),
    .io_x_sx(tlb_OptimizationBarrier_37_io_x_sx),
    .io_x_sr(tlb_OptimizationBarrier_37_io_x_sr),
    .io_x_pw(tlb_OptimizationBarrier_37_io_x_pw),
    .io_x_px(tlb_OptimizationBarrier_37_io_x_px),
    .io_x_pr(tlb_OptimizationBarrier_37_io_x_pr),
    .io_x_ppp(tlb_OptimizationBarrier_37_io_x_ppp),
    .io_x_pal(tlb_OptimizationBarrier_37_io_x_pal),
    .io_x_paa(tlb_OptimizationBarrier_37_io_x_paa),
    .io_x_eff(tlb_OptimizationBarrier_37_io_x_eff),
    .io_x_c(tlb_OptimizationBarrier_37_io_x_c),
    .io_y_ppn(tlb_OptimizationBarrier_37_io_y_ppn),
    .io_y_u(tlb_OptimizationBarrier_37_io_y_u),
    .io_y_ae(tlb_OptimizationBarrier_37_io_y_ae),
    .io_y_sw(tlb_OptimizationBarrier_37_io_y_sw),
    .io_y_sx(tlb_OptimizationBarrier_37_io_y_sx),
    .io_y_sr(tlb_OptimizationBarrier_37_io_y_sr),
    .io_y_pw(tlb_OptimizationBarrier_37_io_y_pw),
    .io_y_px(tlb_OptimizationBarrier_37_io_y_px),
    .io_y_pr(tlb_OptimizationBarrier_37_io_y_pr),
    .io_y_ppp(tlb_OptimizationBarrier_37_io_y_ppp),
    .io_y_pal(tlb_OptimizationBarrier_37_io_y_pal),
    .io_y_paa(tlb_OptimizationBarrier_37_io_y_paa),
    .io_y_eff(tlb_OptimizationBarrier_37_io_y_eff),
    .io_y_c(tlb_OptimizationBarrier_37_io_y_c)
  );
  OptimizationBarrier tlb_OptimizationBarrier_38 ( // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179672.4]
    .io_x_ppn(tlb_OptimizationBarrier_38_io_x_ppn),
    .io_x_u(tlb_OptimizationBarrier_38_io_x_u),
    .io_x_ae(tlb_OptimizationBarrier_38_io_x_ae),
    .io_x_sw(tlb_OptimizationBarrier_38_io_x_sw),
    .io_x_sx(tlb_OptimizationBarrier_38_io_x_sx),
    .io_x_sr(tlb_OptimizationBarrier_38_io_x_sr),
    .io_x_pw(tlb_OptimizationBarrier_38_io_x_pw),
    .io_x_px(tlb_OptimizationBarrier_38_io_x_px),
    .io_x_pr(tlb_OptimizationBarrier_38_io_x_pr),
    .io_x_ppp(tlb_OptimizationBarrier_38_io_x_ppp),
    .io_x_pal(tlb_OptimizationBarrier_38_io_x_pal),
    .io_x_paa(tlb_OptimizationBarrier_38_io_x_paa),
    .io_x_eff(tlb_OptimizationBarrier_38_io_x_eff),
    .io_x_c(tlb_OptimizationBarrier_38_io_x_c),
    .io_y_ppn(tlb_OptimizationBarrier_38_io_y_ppn),
    .io_y_u(tlb_OptimizationBarrier_38_io_y_u),
    .io_y_ae(tlb_OptimizationBarrier_38_io_y_ae),
    .io_y_sw(tlb_OptimizationBarrier_38_io_y_sw),
    .io_y_sx(tlb_OptimizationBarrier_38_io_y_sx),
    .io_y_sr(tlb_OptimizationBarrier_38_io_y_sr),
    .io_y_pw(tlb_OptimizationBarrier_38_io_y_pw),
    .io_y_px(tlb_OptimizationBarrier_38_io_y_px),
    .io_y_pr(tlb_OptimizationBarrier_38_io_y_pr),
    .io_y_ppp(tlb_OptimizationBarrier_38_io_y_ppp),
    .io_y_pal(tlb_OptimizationBarrier_38_io_y_pal),
    .io_y_paa(tlb_OptimizationBarrier_38_io_y_paa),
    .io_y_eff(tlb_OptimizationBarrier_38_io_y_eff),
    .io_y_c(tlb_OptimizationBarrier_38_io_y_c)
  );
  OptimizationBarrier pma_checker_OptimizationBarrier ( // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@176907.4]
    .io_x_ppn(pma_checker_OptimizationBarrier_io_x_ppn),
    .io_x_u(pma_checker_OptimizationBarrier_io_x_u),
    .io_x_ae(pma_checker_OptimizationBarrier_io_x_ae),
    .io_x_sw(pma_checker_OptimizationBarrier_io_x_sw),
    .io_x_sx(pma_checker_OptimizationBarrier_io_x_sx),
    .io_x_sr(pma_checker_OptimizationBarrier_io_x_sr),
    .io_x_pw(pma_checker_OptimizationBarrier_io_x_pw),
    .io_x_px(pma_checker_OptimizationBarrier_io_x_px),
    .io_x_pr(pma_checker_OptimizationBarrier_io_x_pr),
    .io_x_ppp(pma_checker_OptimizationBarrier_io_x_ppp),
    .io_x_pal(pma_checker_OptimizationBarrier_io_x_pal),
    .io_x_paa(pma_checker_OptimizationBarrier_io_x_paa),
    .io_x_eff(pma_checker_OptimizationBarrier_io_x_eff),
    .io_x_c(pma_checker_OptimizationBarrier_io_x_c),
    .io_y_ppn(pma_checker_OptimizationBarrier_io_y_ppn),
    .io_y_u(pma_checker_OptimizationBarrier_io_y_u),
    .io_y_ae(pma_checker_OptimizationBarrier_io_y_ae),
    .io_y_sw(pma_checker_OptimizationBarrier_io_y_sw),
    .io_y_sx(pma_checker_OptimizationBarrier_io_y_sx),
    .io_y_sr(pma_checker_OptimizationBarrier_io_y_sr),
    .io_y_pw(pma_checker_OptimizationBarrier_io_y_pw),
    .io_y_px(pma_checker_OptimizationBarrier_io_y_px),
    .io_y_pr(pma_checker_OptimizationBarrier_io_y_pr),
    .io_y_ppp(pma_checker_OptimizationBarrier_io_y_ppp),
    .io_y_pal(pma_checker_OptimizationBarrier_io_y_pal),
    .io_y_paa(pma_checker_OptimizationBarrier_io_y_paa),
    .io_y_eff(pma_checker_OptimizationBarrier_io_y_eff),
    .io_y_c(pma_checker_OptimizationBarrier_io_y_c)
  );
  PMPChecker pma_checker_pmp ( // @[TLB.scala 190:19:freechips.rocketchip.system.DefaultRV32Config.fir@176928.4]
    .io_prv(pma_checker_pmp_io_prv),
    .io_pmp_0_cfg_l(pma_checker_pmp_io_pmp_0_cfg_l),
    .io_pmp_0_cfg_a(pma_checker_pmp_io_pmp_0_cfg_a),
    .io_pmp_0_cfg_x(pma_checker_pmp_io_pmp_0_cfg_x),
    .io_pmp_0_cfg_w(pma_checker_pmp_io_pmp_0_cfg_w),
    .io_pmp_0_cfg_r(pma_checker_pmp_io_pmp_0_cfg_r),
    .io_pmp_0_addr(pma_checker_pmp_io_pmp_0_addr),
    .io_pmp_0_mask(pma_checker_pmp_io_pmp_0_mask),
    .io_pmp_1_cfg_l(pma_checker_pmp_io_pmp_1_cfg_l),
    .io_pmp_1_cfg_a(pma_checker_pmp_io_pmp_1_cfg_a),
    .io_pmp_1_cfg_x(pma_checker_pmp_io_pmp_1_cfg_x),
    .io_pmp_1_cfg_w(pma_checker_pmp_io_pmp_1_cfg_w),
    .io_pmp_1_cfg_r(pma_checker_pmp_io_pmp_1_cfg_r),
    .io_pmp_1_addr(pma_checker_pmp_io_pmp_1_addr),
    .io_pmp_1_mask(pma_checker_pmp_io_pmp_1_mask),
    .io_pmp_2_cfg_l(pma_checker_pmp_io_pmp_2_cfg_l),
    .io_pmp_2_cfg_a(pma_checker_pmp_io_pmp_2_cfg_a),
    .io_pmp_2_cfg_x(pma_checker_pmp_io_pmp_2_cfg_x),
    .io_pmp_2_cfg_w(pma_checker_pmp_io_pmp_2_cfg_w),
    .io_pmp_2_cfg_r(pma_checker_pmp_io_pmp_2_cfg_r),
    .io_pmp_2_addr(pma_checker_pmp_io_pmp_2_addr),
    .io_pmp_2_mask(pma_checker_pmp_io_pmp_2_mask),
    .io_pmp_3_cfg_l(pma_checker_pmp_io_pmp_3_cfg_l),
    .io_pmp_3_cfg_a(pma_checker_pmp_io_pmp_3_cfg_a),
    .io_pmp_3_cfg_x(pma_checker_pmp_io_pmp_3_cfg_x),
    .io_pmp_3_cfg_w(pma_checker_pmp_io_pmp_3_cfg_w),
    .io_pmp_3_cfg_r(pma_checker_pmp_io_pmp_3_cfg_r),
    .io_pmp_3_addr(pma_checker_pmp_io_pmp_3_addr),
    .io_pmp_3_mask(pma_checker_pmp_io_pmp_3_mask),
    .io_pmp_4_cfg_l(pma_checker_pmp_io_pmp_4_cfg_l),
    .io_pmp_4_cfg_a(pma_checker_pmp_io_pmp_4_cfg_a),
    .io_pmp_4_cfg_x(pma_checker_pmp_io_pmp_4_cfg_x),
    .io_pmp_4_cfg_w(pma_checker_pmp_io_pmp_4_cfg_w),
    .io_pmp_4_cfg_r(pma_checker_pmp_io_pmp_4_cfg_r),
    .io_pmp_4_addr(pma_checker_pmp_io_pmp_4_addr),
    .io_pmp_4_mask(pma_checker_pmp_io_pmp_4_mask),
    .io_pmp_5_cfg_l(pma_checker_pmp_io_pmp_5_cfg_l),
    .io_pmp_5_cfg_a(pma_checker_pmp_io_pmp_5_cfg_a),
    .io_pmp_5_cfg_x(pma_checker_pmp_io_pmp_5_cfg_x),
    .io_pmp_5_cfg_w(pma_checker_pmp_io_pmp_5_cfg_w),
    .io_pmp_5_cfg_r(pma_checker_pmp_io_pmp_5_cfg_r),
    .io_pmp_5_addr(pma_checker_pmp_io_pmp_5_addr),
    .io_pmp_5_mask(pma_checker_pmp_io_pmp_5_mask),
    .io_pmp_6_cfg_l(pma_checker_pmp_io_pmp_6_cfg_l),
    .io_pmp_6_cfg_a(pma_checker_pmp_io_pmp_6_cfg_a),
    .io_pmp_6_cfg_x(pma_checker_pmp_io_pmp_6_cfg_x),
    .io_pmp_6_cfg_w(pma_checker_pmp_io_pmp_6_cfg_w),
    .io_pmp_6_cfg_r(pma_checker_pmp_io_pmp_6_cfg_r),
    .io_pmp_6_addr(pma_checker_pmp_io_pmp_6_addr),
    .io_pmp_6_mask(pma_checker_pmp_io_pmp_6_mask),
    .io_pmp_7_cfg_l(pma_checker_pmp_io_pmp_7_cfg_l),
    .io_pmp_7_cfg_a(pma_checker_pmp_io_pmp_7_cfg_a),
    .io_pmp_7_cfg_x(pma_checker_pmp_io_pmp_7_cfg_x),
    .io_pmp_7_cfg_w(pma_checker_pmp_io_pmp_7_cfg_w),
    .io_pmp_7_cfg_r(pma_checker_pmp_io_pmp_7_cfg_r),
    .io_pmp_7_addr(pma_checker_pmp_io_pmp_7_addr),
    .io_pmp_7_mask(pma_checker_pmp_io_pmp_7_mask),
    .io_addr(pma_checker_pmp_io_addr),
    .io_r(pma_checker_pmp_io_r),
    .io_w(pma_checker_pmp_io_w),
    .io_x(pma_checker_pmp_io_x)
  );
  OptimizationBarrier pma_checker_OptimizationBarrier_1 ( // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@177629.4]
    .io_x_ppn(pma_checker_OptimizationBarrier_1_io_x_ppn),
    .io_x_u(pma_checker_OptimizationBarrier_1_io_x_u),
    .io_x_ae(pma_checker_OptimizationBarrier_1_io_x_ae),
    .io_x_sw(pma_checker_OptimizationBarrier_1_io_x_sw),
    .io_x_sx(pma_checker_OptimizationBarrier_1_io_x_sx),
    .io_x_sr(pma_checker_OptimizationBarrier_1_io_x_sr),
    .io_x_pw(pma_checker_OptimizationBarrier_1_io_x_pw),
    .io_x_px(pma_checker_OptimizationBarrier_1_io_x_px),
    .io_x_pr(pma_checker_OptimizationBarrier_1_io_x_pr),
    .io_x_ppp(pma_checker_OptimizationBarrier_1_io_x_ppp),
    .io_x_pal(pma_checker_OptimizationBarrier_1_io_x_pal),
    .io_x_paa(pma_checker_OptimizationBarrier_1_io_x_paa),
    .io_x_eff(pma_checker_OptimizationBarrier_1_io_x_eff),
    .io_x_c(pma_checker_OptimizationBarrier_1_io_x_c),
    .io_y_ppn(pma_checker_OptimizationBarrier_1_io_y_ppn),
    .io_y_u(pma_checker_OptimizationBarrier_1_io_y_u),
    .io_y_ae(pma_checker_OptimizationBarrier_1_io_y_ae),
    .io_y_sw(pma_checker_OptimizationBarrier_1_io_y_sw),
    .io_y_sx(pma_checker_OptimizationBarrier_1_io_y_sx),
    .io_y_sr(pma_checker_OptimizationBarrier_1_io_y_sr),
    .io_y_pw(pma_checker_OptimizationBarrier_1_io_y_pw),
    .io_y_px(pma_checker_OptimizationBarrier_1_io_y_px),
    .io_y_pr(pma_checker_OptimizationBarrier_1_io_y_pr),
    .io_y_ppp(pma_checker_OptimizationBarrier_1_io_y_ppp),
    .io_y_pal(pma_checker_OptimizationBarrier_1_io_y_pal),
    .io_y_paa(pma_checker_OptimizationBarrier_1_io_y_paa),
    .io_y_eff(pma_checker_OptimizationBarrier_1_io_y_eff),
    .io_y_c(pma_checker_OptimizationBarrier_1_io_y_c)
  );
  OptimizationBarrier pma_checker_OptimizationBarrier_2 ( // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@177672.4]
    .io_x_ppn(pma_checker_OptimizationBarrier_2_io_x_ppn),
    .io_x_u(pma_checker_OptimizationBarrier_2_io_x_u),
    .io_x_ae(pma_checker_OptimizationBarrier_2_io_x_ae),
    .io_x_sw(pma_checker_OptimizationBarrier_2_io_x_sw),
    .io_x_sx(pma_checker_OptimizationBarrier_2_io_x_sx),
    .io_x_sr(pma_checker_OptimizationBarrier_2_io_x_sr),
    .io_x_pw(pma_checker_OptimizationBarrier_2_io_x_pw),
    .io_x_px(pma_checker_OptimizationBarrier_2_io_x_px),
    .io_x_pr(pma_checker_OptimizationBarrier_2_io_x_pr),
    .io_x_ppp(pma_checker_OptimizationBarrier_2_io_x_ppp),
    .io_x_pal(pma_checker_OptimizationBarrier_2_io_x_pal),
    .io_x_paa(pma_checker_OptimizationBarrier_2_io_x_paa),
    .io_x_eff(pma_checker_OptimizationBarrier_2_io_x_eff),
    .io_x_c(pma_checker_OptimizationBarrier_2_io_x_c),
    .io_y_ppn(pma_checker_OptimizationBarrier_2_io_y_ppn),
    .io_y_u(pma_checker_OptimizationBarrier_2_io_y_u),
    .io_y_ae(pma_checker_OptimizationBarrier_2_io_y_ae),
    .io_y_sw(pma_checker_OptimizationBarrier_2_io_y_sw),
    .io_y_sx(pma_checker_OptimizationBarrier_2_io_y_sx),
    .io_y_sr(pma_checker_OptimizationBarrier_2_io_y_sr),
    .io_y_pw(pma_checker_OptimizationBarrier_2_io_y_pw),
    .io_y_px(pma_checker_OptimizationBarrier_2_io_y_px),
    .io_y_pr(pma_checker_OptimizationBarrier_2_io_y_pr),
    .io_y_ppp(pma_checker_OptimizationBarrier_2_io_y_ppp),
    .io_y_pal(pma_checker_OptimizationBarrier_2_io_y_pal),
    .io_y_paa(pma_checker_OptimizationBarrier_2_io_y_paa),
    .io_y_eff(pma_checker_OptimizationBarrier_2_io_y_eff),
    .io_y_c(pma_checker_OptimizationBarrier_2_io_y_c)
  );
  OptimizationBarrier pma_checker_OptimizationBarrier_3 ( // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@177715.4]
    .io_x_ppn(pma_checker_OptimizationBarrier_3_io_x_ppn),
    .io_x_u(pma_checker_OptimizationBarrier_3_io_x_u),
    .io_x_ae(pma_checker_OptimizationBarrier_3_io_x_ae),
    .io_x_sw(pma_checker_OptimizationBarrier_3_io_x_sw),
    .io_x_sx(pma_checker_OptimizationBarrier_3_io_x_sx),
    .io_x_sr(pma_checker_OptimizationBarrier_3_io_x_sr),
    .io_x_pw(pma_checker_OptimizationBarrier_3_io_x_pw),
    .io_x_px(pma_checker_OptimizationBarrier_3_io_x_px),
    .io_x_pr(pma_checker_OptimizationBarrier_3_io_x_pr),
    .io_x_ppp(pma_checker_OptimizationBarrier_3_io_x_ppp),
    .io_x_pal(pma_checker_OptimizationBarrier_3_io_x_pal),
    .io_x_paa(pma_checker_OptimizationBarrier_3_io_x_paa),
    .io_x_eff(pma_checker_OptimizationBarrier_3_io_x_eff),
    .io_x_c(pma_checker_OptimizationBarrier_3_io_x_c),
    .io_y_ppn(pma_checker_OptimizationBarrier_3_io_y_ppn),
    .io_y_u(pma_checker_OptimizationBarrier_3_io_y_u),
    .io_y_ae(pma_checker_OptimizationBarrier_3_io_y_ae),
    .io_y_sw(pma_checker_OptimizationBarrier_3_io_y_sw),
    .io_y_sx(pma_checker_OptimizationBarrier_3_io_y_sx),
    .io_y_sr(pma_checker_OptimizationBarrier_3_io_y_sr),
    .io_y_pw(pma_checker_OptimizationBarrier_3_io_y_pw),
    .io_y_px(pma_checker_OptimizationBarrier_3_io_y_px),
    .io_y_pr(pma_checker_OptimizationBarrier_3_io_y_pr),
    .io_y_ppp(pma_checker_OptimizationBarrier_3_io_y_ppp),
    .io_y_pal(pma_checker_OptimizationBarrier_3_io_y_pal),
    .io_y_paa(pma_checker_OptimizationBarrier_3_io_y_paa),
    .io_y_eff(pma_checker_OptimizationBarrier_3_io_y_eff),
    .io_y_c(pma_checker_OptimizationBarrier_3_io_y_c)
  );
  OptimizationBarrier pma_checker_OptimizationBarrier_4 ( // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@177758.4]
    .io_x_ppn(pma_checker_OptimizationBarrier_4_io_x_ppn),
    .io_x_u(pma_checker_OptimizationBarrier_4_io_x_u),
    .io_x_ae(pma_checker_OptimizationBarrier_4_io_x_ae),
    .io_x_sw(pma_checker_OptimizationBarrier_4_io_x_sw),
    .io_x_sx(pma_checker_OptimizationBarrier_4_io_x_sx),
    .io_x_sr(pma_checker_OptimizationBarrier_4_io_x_sr),
    .io_x_pw(pma_checker_OptimizationBarrier_4_io_x_pw),
    .io_x_px(pma_checker_OptimizationBarrier_4_io_x_px),
    .io_x_pr(pma_checker_OptimizationBarrier_4_io_x_pr),
    .io_x_ppp(pma_checker_OptimizationBarrier_4_io_x_ppp),
    .io_x_pal(pma_checker_OptimizationBarrier_4_io_x_pal),
    .io_x_paa(pma_checker_OptimizationBarrier_4_io_x_paa),
    .io_x_eff(pma_checker_OptimizationBarrier_4_io_x_eff),
    .io_x_c(pma_checker_OptimizationBarrier_4_io_x_c),
    .io_y_ppn(pma_checker_OptimizationBarrier_4_io_y_ppn),
    .io_y_u(pma_checker_OptimizationBarrier_4_io_y_u),
    .io_y_ae(pma_checker_OptimizationBarrier_4_io_y_ae),
    .io_y_sw(pma_checker_OptimizationBarrier_4_io_y_sw),
    .io_y_sx(pma_checker_OptimizationBarrier_4_io_y_sx),
    .io_y_sr(pma_checker_OptimizationBarrier_4_io_y_sr),
    .io_y_pw(pma_checker_OptimizationBarrier_4_io_y_pw),
    .io_y_px(pma_checker_OptimizationBarrier_4_io_y_px),
    .io_y_pr(pma_checker_OptimizationBarrier_4_io_y_pr),
    .io_y_ppp(pma_checker_OptimizationBarrier_4_io_y_ppp),
    .io_y_pal(pma_checker_OptimizationBarrier_4_io_y_pal),
    .io_y_paa(pma_checker_OptimizationBarrier_4_io_y_paa),
    .io_y_eff(pma_checker_OptimizationBarrier_4_io_y_eff),
    .io_y_c(pma_checker_OptimizationBarrier_4_io_y_c)
  );
  OptimizationBarrier pma_checker_OptimizationBarrier_5 ( // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@177801.4]
    .io_x_ppn(pma_checker_OptimizationBarrier_5_io_x_ppn),
    .io_x_u(pma_checker_OptimizationBarrier_5_io_x_u),
    .io_x_ae(pma_checker_OptimizationBarrier_5_io_x_ae),
    .io_x_sw(pma_checker_OptimizationBarrier_5_io_x_sw),
    .io_x_sx(pma_checker_OptimizationBarrier_5_io_x_sx),
    .io_x_sr(pma_checker_OptimizationBarrier_5_io_x_sr),
    .io_x_pw(pma_checker_OptimizationBarrier_5_io_x_pw),
    .io_x_px(pma_checker_OptimizationBarrier_5_io_x_px),
    .io_x_pr(pma_checker_OptimizationBarrier_5_io_x_pr),
    .io_x_ppp(pma_checker_OptimizationBarrier_5_io_x_ppp),
    .io_x_pal(pma_checker_OptimizationBarrier_5_io_x_pal),
    .io_x_paa(pma_checker_OptimizationBarrier_5_io_x_paa),
    .io_x_eff(pma_checker_OptimizationBarrier_5_io_x_eff),
    .io_x_c(pma_checker_OptimizationBarrier_5_io_x_c),
    .io_y_ppn(pma_checker_OptimizationBarrier_5_io_y_ppn),
    .io_y_u(pma_checker_OptimizationBarrier_5_io_y_u),
    .io_y_ae(pma_checker_OptimizationBarrier_5_io_y_ae),
    .io_y_sw(pma_checker_OptimizationBarrier_5_io_y_sw),
    .io_y_sx(pma_checker_OptimizationBarrier_5_io_y_sx),
    .io_y_sr(pma_checker_OptimizationBarrier_5_io_y_sr),
    .io_y_pw(pma_checker_OptimizationBarrier_5_io_y_pw),
    .io_y_px(pma_checker_OptimizationBarrier_5_io_y_px),
    .io_y_pr(pma_checker_OptimizationBarrier_5_io_y_pr),
    .io_y_ppp(pma_checker_OptimizationBarrier_5_io_y_ppp),
    .io_y_pal(pma_checker_OptimizationBarrier_5_io_y_pal),
    .io_y_paa(pma_checker_OptimizationBarrier_5_io_y_paa),
    .io_y_eff(pma_checker_OptimizationBarrier_5_io_y_eff),
    .io_y_c(pma_checker_OptimizationBarrier_5_io_y_c)
  );
  OptimizationBarrier pma_checker_OptimizationBarrier_6 ( // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@177844.4]
    .io_x_ppn(pma_checker_OptimizationBarrier_6_io_x_ppn),
    .io_x_u(pma_checker_OptimizationBarrier_6_io_x_u),
    .io_x_ae(pma_checker_OptimizationBarrier_6_io_x_ae),
    .io_x_sw(pma_checker_OptimizationBarrier_6_io_x_sw),
    .io_x_sx(pma_checker_OptimizationBarrier_6_io_x_sx),
    .io_x_sr(pma_checker_OptimizationBarrier_6_io_x_sr),
    .io_x_pw(pma_checker_OptimizationBarrier_6_io_x_pw),
    .io_x_px(pma_checker_OptimizationBarrier_6_io_x_px),
    .io_x_pr(pma_checker_OptimizationBarrier_6_io_x_pr),
    .io_x_ppp(pma_checker_OptimizationBarrier_6_io_x_ppp),
    .io_x_pal(pma_checker_OptimizationBarrier_6_io_x_pal),
    .io_x_paa(pma_checker_OptimizationBarrier_6_io_x_paa),
    .io_x_eff(pma_checker_OptimizationBarrier_6_io_x_eff),
    .io_x_c(pma_checker_OptimizationBarrier_6_io_x_c),
    .io_y_ppn(pma_checker_OptimizationBarrier_6_io_y_ppn),
    .io_y_u(pma_checker_OptimizationBarrier_6_io_y_u),
    .io_y_ae(pma_checker_OptimizationBarrier_6_io_y_ae),
    .io_y_sw(pma_checker_OptimizationBarrier_6_io_y_sw),
    .io_y_sx(pma_checker_OptimizationBarrier_6_io_y_sx),
    .io_y_sr(pma_checker_OptimizationBarrier_6_io_y_sr),
    .io_y_pw(pma_checker_OptimizationBarrier_6_io_y_pw),
    .io_y_px(pma_checker_OptimizationBarrier_6_io_y_px),
    .io_y_pr(pma_checker_OptimizationBarrier_6_io_y_pr),
    .io_y_ppp(pma_checker_OptimizationBarrier_6_io_y_ppp),
    .io_y_pal(pma_checker_OptimizationBarrier_6_io_y_pal),
    .io_y_paa(pma_checker_OptimizationBarrier_6_io_y_paa),
    .io_y_eff(pma_checker_OptimizationBarrier_6_io_y_eff),
    .io_y_c(pma_checker_OptimizationBarrier_6_io_y_c)
  );
  OptimizationBarrier pma_checker_OptimizationBarrier_7 ( // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@177887.4]
    .io_x_ppn(pma_checker_OptimizationBarrier_7_io_x_ppn),
    .io_x_u(pma_checker_OptimizationBarrier_7_io_x_u),
    .io_x_ae(pma_checker_OptimizationBarrier_7_io_x_ae),
    .io_x_sw(pma_checker_OptimizationBarrier_7_io_x_sw),
    .io_x_sx(pma_checker_OptimizationBarrier_7_io_x_sx),
    .io_x_sr(pma_checker_OptimizationBarrier_7_io_x_sr),
    .io_x_pw(pma_checker_OptimizationBarrier_7_io_x_pw),
    .io_x_px(pma_checker_OptimizationBarrier_7_io_x_px),
    .io_x_pr(pma_checker_OptimizationBarrier_7_io_x_pr),
    .io_x_ppp(pma_checker_OptimizationBarrier_7_io_x_ppp),
    .io_x_pal(pma_checker_OptimizationBarrier_7_io_x_pal),
    .io_x_paa(pma_checker_OptimizationBarrier_7_io_x_paa),
    .io_x_eff(pma_checker_OptimizationBarrier_7_io_x_eff),
    .io_x_c(pma_checker_OptimizationBarrier_7_io_x_c),
    .io_y_ppn(pma_checker_OptimizationBarrier_7_io_y_ppn),
    .io_y_u(pma_checker_OptimizationBarrier_7_io_y_u),
    .io_y_ae(pma_checker_OptimizationBarrier_7_io_y_ae),
    .io_y_sw(pma_checker_OptimizationBarrier_7_io_y_sw),
    .io_y_sx(pma_checker_OptimizationBarrier_7_io_y_sx),
    .io_y_sr(pma_checker_OptimizationBarrier_7_io_y_sr),
    .io_y_pw(pma_checker_OptimizationBarrier_7_io_y_pw),
    .io_y_px(pma_checker_OptimizationBarrier_7_io_y_px),
    .io_y_pr(pma_checker_OptimizationBarrier_7_io_y_pr),
    .io_y_ppp(pma_checker_OptimizationBarrier_7_io_y_ppp),
    .io_y_pal(pma_checker_OptimizationBarrier_7_io_y_pal),
    .io_y_paa(pma_checker_OptimizationBarrier_7_io_y_paa),
    .io_y_eff(pma_checker_OptimizationBarrier_7_io_y_eff),
    .io_y_c(pma_checker_OptimizationBarrier_7_io_y_c)
  );
  OptimizationBarrier pma_checker_OptimizationBarrier_8 ( // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@177930.4]
    .io_x_ppn(pma_checker_OptimizationBarrier_8_io_x_ppn),
    .io_x_u(pma_checker_OptimizationBarrier_8_io_x_u),
    .io_x_ae(pma_checker_OptimizationBarrier_8_io_x_ae),
    .io_x_sw(pma_checker_OptimizationBarrier_8_io_x_sw),
    .io_x_sx(pma_checker_OptimizationBarrier_8_io_x_sx),
    .io_x_sr(pma_checker_OptimizationBarrier_8_io_x_sr),
    .io_x_pw(pma_checker_OptimizationBarrier_8_io_x_pw),
    .io_x_px(pma_checker_OptimizationBarrier_8_io_x_px),
    .io_x_pr(pma_checker_OptimizationBarrier_8_io_x_pr),
    .io_x_ppp(pma_checker_OptimizationBarrier_8_io_x_ppp),
    .io_x_pal(pma_checker_OptimizationBarrier_8_io_x_pal),
    .io_x_paa(pma_checker_OptimizationBarrier_8_io_x_paa),
    .io_x_eff(pma_checker_OptimizationBarrier_8_io_x_eff),
    .io_x_c(pma_checker_OptimizationBarrier_8_io_x_c),
    .io_y_ppn(pma_checker_OptimizationBarrier_8_io_y_ppn),
    .io_y_u(pma_checker_OptimizationBarrier_8_io_y_u),
    .io_y_ae(pma_checker_OptimizationBarrier_8_io_y_ae),
    .io_y_sw(pma_checker_OptimizationBarrier_8_io_y_sw),
    .io_y_sx(pma_checker_OptimizationBarrier_8_io_y_sx),
    .io_y_sr(pma_checker_OptimizationBarrier_8_io_y_sr),
    .io_y_pw(pma_checker_OptimizationBarrier_8_io_y_pw),
    .io_y_px(pma_checker_OptimizationBarrier_8_io_y_px),
    .io_y_pr(pma_checker_OptimizationBarrier_8_io_y_pr),
    .io_y_ppp(pma_checker_OptimizationBarrier_8_io_y_ppp),
    .io_y_pal(pma_checker_OptimizationBarrier_8_io_y_pal),
    .io_y_paa(pma_checker_OptimizationBarrier_8_io_y_paa),
    .io_y_eff(pma_checker_OptimizationBarrier_8_io_y_eff),
    .io_y_c(pma_checker_OptimizationBarrier_8_io_y_c)
  );
  OptimizationBarrier pma_checker_OptimizationBarrier_9 ( // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@177972.4]
    .io_x_ppn(pma_checker_OptimizationBarrier_9_io_x_ppn),
    .io_x_u(pma_checker_OptimizationBarrier_9_io_x_u),
    .io_x_ae(pma_checker_OptimizationBarrier_9_io_x_ae),
    .io_x_sw(pma_checker_OptimizationBarrier_9_io_x_sw),
    .io_x_sx(pma_checker_OptimizationBarrier_9_io_x_sx),
    .io_x_sr(pma_checker_OptimizationBarrier_9_io_x_sr),
    .io_x_pw(pma_checker_OptimizationBarrier_9_io_x_pw),
    .io_x_px(pma_checker_OptimizationBarrier_9_io_x_px),
    .io_x_pr(pma_checker_OptimizationBarrier_9_io_x_pr),
    .io_x_ppp(pma_checker_OptimizationBarrier_9_io_x_ppp),
    .io_x_pal(pma_checker_OptimizationBarrier_9_io_x_pal),
    .io_x_paa(pma_checker_OptimizationBarrier_9_io_x_paa),
    .io_x_eff(pma_checker_OptimizationBarrier_9_io_x_eff),
    .io_x_c(pma_checker_OptimizationBarrier_9_io_x_c),
    .io_y_ppn(pma_checker_OptimizationBarrier_9_io_y_ppn),
    .io_y_u(pma_checker_OptimizationBarrier_9_io_y_u),
    .io_y_ae(pma_checker_OptimizationBarrier_9_io_y_ae),
    .io_y_sw(pma_checker_OptimizationBarrier_9_io_y_sw),
    .io_y_sx(pma_checker_OptimizationBarrier_9_io_y_sx),
    .io_y_sr(pma_checker_OptimizationBarrier_9_io_y_sr),
    .io_y_pw(pma_checker_OptimizationBarrier_9_io_y_pw),
    .io_y_px(pma_checker_OptimizationBarrier_9_io_y_px),
    .io_y_pr(pma_checker_OptimizationBarrier_9_io_y_pr),
    .io_y_ppp(pma_checker_OptimizationBarrier_9_io_y_ppp),
    .io_y_pal(pma_checker_OptimizationBarrier_9_io_y_pal),
    .io_y_paa(pma_checker_OptimizationBarrier_9_io_y_paa),
    .io_y_eff(pma_checker_OptimizationBarrier_9_io_y_eff),
    .io_y_c(pma_checker_OptimizationBarrier_9_io_y_c)
  );
  OptimizationBarrier pma_checker_OptimizationBarrier_10 ( // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178021.4]
    .io_x_ppn(pma_checker_OptimizationBarrier_10_io_x_ppn),
    .io_x_u(pma_checker_OptimizationBarrier_10_io_x_u),
    .io_x_ae(pma_checker_OptimizationBarrier_10_io_x_ae),
    .io_x_sw(pma_checker_OptimizationBarrier_10_io_x_sw),
    .io_x_sx(pma_checker_OptimizationBarrier_10_io_x_sx),
    .io_x_sr(pma_checker_OptimizationBarrier_10_io_x_sr),
    .io_x_pw(pma_checker_OptimizationBarrier_10_io_x_pw),
    .io_x_px(pma_checker_OptimizationBarrier_10_io_x_px),
    .io_x_pr(pma_checker_OptimizationBarrier_10_io_x_pr),
    .io_x_ppp(pma_checker_OptimizationBarrier_10_io_x_ppp),
    .io_x_pal(pma_checker_OptimizationBarrier_10_io_x_pal),
    .io_x_paa(pma_checker_OptimizationBarrier_10_io_x_paa),
    .io_x_eff(pma_checker_OptimizationBarrier_10_io_x_eff),
    .io_x_c(pma_checker_OptimizationBarrier_10_io_x_c),
    .io_y_ppn(pma_checker_OptimizationBarrier_10_io_y_ppn),
    .io_y_u(pma_checker_OptimizationBarrier_10_io_y_u),
    .io_y_ae(pma_checker_OptimizationBarrier_10_io_y_ae),
    .io_y_sw(pma_checker_OptimizationBarrier_10_io_y_sw),
    .io_y_sx(pma_checker_OptimizationBarrier_10_io_y_sx),
    .io_y_sr(pma_checker_OptimizationBarrier_10_io_y_sr),
    .io_y_pw(pma_checker_OptimizationBarrier_10_io_y_pw),
    .io_y_px(pma_checker_OptimizationBarrier_10_io_y_px),
    .io_y_pr(pma_checker_OptimizationBarrier_10_io_y_pr),
    .io_y_ppp(pma_checker_OptimizationBarrier_10_io_y_ppp),
    .io_y_pal(pma_checker_OptimizationBarrier_10_io_y_pal),
    .io_y_paa(pma_checker_OptimizationBarrier_10_io_y_paa),
    .io_y_eff(pma_checker_OptimizationBarrier_10_io_y_eff),
    .io_y_c(pma_checker_OptimizationBarrier_10_io_y_c)
  );
  OptimizationBarrier pma_checker_OptimizationBarrier_11 ( // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178070.4]
    .io_x_ppn(pma_checker_OptimizationBarrier_11_io_x_ppn),
    .io_x_u(pma_checker_OptimizationBarrier_11_io_x_u),
    .io_x_ae(pma_checker_OptimizationBarrier_11_io_x_ae),
    .io_x_sw(pma_checker_OptimizationBarrier_11_io_x_sw),
    .io_x_sx(pma_checker_OptimizationBarrier_11_io_x_sx),
    .io_x_sr(pma_checker_OptimizationBarrier_11_io_x_sr),
    .io_x_pw(pma_checker_OptimizationBarrier_11_io_x_pw),
    .io_x_px(pma_checker_OptimizationBarrier_11_io_x_px),
    .io_x_pr(pma_checker_OptimizationBarrier_11_io_x_pr),
    .io_x_ppp(pma_checker_OptimizationBarrier_11_io_x_ppp),
    .io_x_pal(pma_checker_OptimizationBarrier_11_io_x_pal),
    .io_x_paa(pma_checker_OptimizationBarrier_11_io_x_paa),
    .io_x_eff(pma_checker_OptimizationBarrier_11_io_x_eff),
    .io_x_c(pma_checker_OptimizationBarrier_11_io_x_c),
    .io_y_ppn(pma_checker_OptimizationBarrier_11_io_y_ppn),
    .io_y_u(pma_checker_OptimizationBarrier_11_io_y_u),
    .io_y_ae(pma_checker_OptimizationBarrier_11_io_y_ae),
    .io_y_sw(pma_checker_OptimizationBarrier_11_io_y_sw),
    .io_y_sx(pma_checker_OptimizationBarrier_11_io_y_sx),
    .io_y_sr(pma_checker_OptimizationBarrier_11_io_y_sr),
    .io_y_pw(pma_checker_OptimizationBarrier_11_io_y_pw),
    .io_y_px(pma_checker_OptimizationBarrier_11_io_y_px),
    .io_y_pr(pma_checker_OptimizationBarrier_11_io_y_pr),
    .io_y_ppp(pma_checker_OptimizationBarrier_11_io_y_ppp),
    .io_y_pal(pma_checker_OptimizationBarrier_11_io_y_pal),
    .io_y_paa(pma_checker_OptimizationBarrier_11_io_y_paa),
    .io_y_eff(pma_checker_OptimizationBarrier_11_io_y_eff),
    .io_y_c(pma_checker_OptimizationBarrier_11_io_y_c)
  );
  OptimizationBarrier pma_checker_OptimizationBarrier_12 ( // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178119.4]
    .io_x_ppn(pma_checker_OptimizationBarrier_12_io_x_ppn),
    .io_x_u(pma_checker_OptimizationBarrier_12_io_x_u),
    .io_x_ae(pma_checker_OptimizationBarrier_12_io_x_ae),
    .io_x_sw(pma_checker_OptimizationBarrier_12_io_x_sw),
    .io_x_sx(pma_checker_OptimizationBarrier_12_io_x_sx),
    .io_x_sr(pma_checker_OptimizationBarrier_12_io_x_sr),
    .io_x_pw(pma_checker_OptimizationBarrier_12_io_x_pw),
    .io_x_px(pma_checker_OptimizationBarrier_12_io_x_px),
    .io_x_pr(pma_checker_OptimizationBarrier_12_io_x_pr),
    .io_x_ppp(pma_checker_OptimizationBarrier_12_io_x_ppp),
    .io_x_pal(pma_checker_OptimizationBarrier_12_io_x_pal),
    .io_x_paa(pma_checker_OptimizationBarrier_12_io_x_paa),
    .io_x_eff(pma_checker_OptimizationBarrier_12_io_x_eff),
    .io_x_c(pma_checker_OptimizationBarrier_12_io_x_c),
    .io_y_ppn(pma_checker_OptimizationBarrier_12_io_y_ppn),
    .io_y_u(pma_checker_OptimizationBarrier_12_io_y_u),
    .io_y_ae(pma_checker_OptimizationBarrier_12_io_y_ae),
    .io_y_sw(pma_checker_OptimizationBarrier_12_io_y_sw),
    .io_y_sx(pma_checker_OptimizationBarrier_12_io_y_sx),
    .io_y_sr(pma_checker_OptimizationBarrier_12_io_y_sr),
    .io_y_pw(pma_checker_OptimizationBarrier_12_io_y_pw),
    .io_y_px(pma_checker_OptimizationBarrier_12_io_y_px),
    .io_y_pr(pma_checker_OptimizationBarrier_12_io_y_pr),
    .io_y_ppp(pma_checker_OptimizationBarrier_12_io_y_ppp),
    .io_y_pal(pma_checker_OptimizationBarrier_12_io_y_pal),
    .io_y_paa(pma_checker_OptimizationBarrier_12_io_y_paa),
    .io_y_eff(pma_checker_OptimizationBarrier_12_io_y_eff),
    .io_y_c(pma_checker_OptimizationBarrier_12_io_y_c)
  );
  OptimizationBarrier pma_checker_OptimizationBarrier_13 ( // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178168.4]
    .io_x_ppn(pma_checker_OptimizationBarrier_13_io_x_ppn),
    .io_x_u(pma_checker_OptimizationBarrier_13_io_x_u),
    .io_x_ae(pma_checker_OptimizationBarrier_13_io_x_ae),
    .io_x_sw(pma_checker_OptimizationBarrier_13_io_x_sw),
    .io_x_sx(pma_checker_OptimizationBarrier_13_io_x_sx),
    .io_x_sr(pma_checker_OptimizationBarrier_13_io_x_sr),
    .io_x_pw(pma_checker_OptimizationBarrier_13_io_x_pw),
    .io_x_px(pma_checker_OptimizationBarrier_13_io_x_px),
    .io_x_pr(pma_checker_OptimizationBarrier_13_io_x_pr),
    .io_x_ppp(pma_checker_OptimizationBarrier_13_io_x_ppp),
    .io_x_pal(pma_checker_OptimizationBarrier_13_io_x_pal),
    .io_x_paa(pma_checker_OptimizationBarrier_13_io_x_paa),
    .io_x_eff(pma_checker_OptimizationBarrier_13_io_x_eff),
    .io_x_c(pma_checker_OptimizationBarrier_13_io_x_c),
    .io_y_ppn(pma_checker_OptimizationBarrier_13_io_y_ppn),
    .io_y_u(pma_checker_OptimizationBarrier_13_io_y_u),
    .io_y_ae(pma_checker_OptimizationBarrier_13_io_y_ae),
    .io_y_sw(pma_checker_OptimizationBarrier_13_io_y_sw),
    .io_y_sx(pma_checker_OptimizationBarrier_13_io_y_sx),
    .io_y_sr(pma_checker_OptimizationBarrier_13_io_y_sr),
    .io_y_pw(pma_checker_OptimizationBarrier_13_io_y_pw),
    .io_y_px(pma_checker_OptimizationBarrier_13_io_y_px),
    .io_y_pr(pma_checker_OptimizationBarrier_13_io_y_pr),
    .io_y_ppp(pma_checker_OptimizationBarrier_13_io_y_ppp),
    .io_y_pal(pma_checker_OptimizationBarrier_13_io_y_pal),
    .io_y_paa(pma_checker_OptimizationBarrier_13_io_y_paa),
    .io_y_eff(pma_checker_OptimizationBarrier_13_io_y_eff),
    .io_y_c(pma_checker_OptimizationBarrier_13_io_y_c)
  );
  OptimizationBarrier pma_checker_OptimizationBarrier_14 ( // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178649.4]
    .io_x_ppn(pma_checker_OptimizationBarrier_14_io_x_ppn),
    .io_x_u(pma_checker_OptimizationBarrier_14_io_x_u),
    .io_x_ae(pma_checker_OptimizationBarrier_14_io_x_ae),
    .io_x_sw(pma_checker_OptimizationBarrier_14_io_x_sw),
    .io_x_sx(pma_checker_OptimizationBarrier_14_io_x_sx),
    .io_x_sr(pma_checker_OptimizationBarrier_14_io_x_sr),
    .io_x_pw(pma_checker_OptimizationBarrier_14_io_x_pw),
    .io_x_px(pma_checker_OptimizationBarrier_14_io_x_px),
    .io_x_pr(pma_checker_OptimizationBarrier_14_io_x_pr),
    .io_x_ppp(pma_checker_OptimizationBarrier_14_io_x_ppp),
    .io_x_pal(pma_checker_OptimizationBarrier_14_io_x_pal),
    .io_x_paa(pma_checker_OptimizationBarrier_14_io_x_paa),
    .io_x_eff(pma_checker_OptimizationBarrier_14_io_x_eff),
    .io_x_c(pma_checker_OptimizationBarrier_14_io_x_c),
    .io_y_ppn(pma_checker_OptimizationBarrier_14_io_y_ppn),
    .io_y_u(pma_checker_OptimizationBarrier_14_io_y_u),
    .io_y_ae(pma_checker_OptimizationBarrier_14_io_y_ae),
    .io_y_sw(pma_checker_OptimizationBarrier_14_io_y_sw),
    .io_y_sx(pma_checker_OptimizationBarrier_14_io_y_sx),
    .io_y_sr(pma_checker_OptimizationBarrier_14_io_y_sr),
    .io_y_pw(pma_checker_OptimizationBarrier_14_io_y_pw),
    .io_y_px(pma_checker_OptimizationBarrier_14_io_y_px),
    .io_y_pr(pma_checker_OptimizationBarrier_14_io_y_pr),
    .io_y_ppp(pma_checker_OptimizationBarrier_14_io_y_ppp),
    .io_y_pal(pma_checker_OptimizationBarrier_14_io_y_pal),
    .io_y_paa(pma_checker_OptimizationBarrier_14_io_y_paa),
    .io_y_eff(pma_checker_OptimizationBarrier_14_io_y_eff),
    .io_y_c(pma_checker_OptimizationBarrier_14_io_y_c)
  );
  OptimizationBarrier pma_checker_OptimizationBarrier_15 ( // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178692.4]
    .io_x_ppn(pma_checker_OptimizationBarrier_15_io_x_ppn),
    .io_x_u(pma_checker_OptimizationBarrier_15_io_x_u),
    .io_x_ae(pma_checker_OptimizationBarrier_15_io_x_ae),
    .io_x_sw(pma_checker_OptimizationBarrier_15_io_x_sw),
    .io_x_sx(pma_checker_OptimizationBarrier_15_io_x_sx),
    .io_x_sr(pma_checker_OptimizationBarrier_15_io_x_sr),
    .io_x_pw(pma_checker_OptimizationBarrier_15_io_x_pw),
    .io_x_px(pma_checker_OptimizationBarrier_15_io_x_px),
    .io_x_pr(pma_checker_OptimizationBarrier_15_io_x_pr),
    .io_x_ppp(pma_checker_OptimizationBarrier_15_io_x_ppp),
    .io_x_pal(pma_checker_OptimizationBarrier_15_io_x_pal),
    .io_x_paa(pma_checker_OptimizationBarrier_15_io_x_paa),
    .io_x_eff(pma_checker_OptimizationBarrier_15_io_x_eff),
    .io_x_c(pma_checker_OptimizationBarrier_15_io_x_c),
    .io_y_ppn(pma_checker_OptimizationBarrier_15_io_y_ppn),
    .io_y_u(pma_checker_OptimizationBarrier_15_io_y_u),
    .io_y_ae(pma_checker_OptimizationBarrier_15_io_y_ae),
    .io_y_sw(pma_checker_OptimizationBarrier_15_io_y_sw),
    .io_y_sx(pma_checker_OptimizationBarrier_15_io_y_sx),
    .io_y_sr(pma_checker_OptimizationBarrier_15_io_y_sr),
    .io_y_pw(pma_checker_OptimizationBarrier_15_io_y_pw),
    .io_y_px(pma_checker_OptimizationBarrier_15_io_y_px),
    .io_y_pr(pma_checker_OptimizationBarrier_15_io_y_pr),
    .io_y_ppp(pma_checker_OptimizationBarrier_15_io_y_ppp),
    .io_y_pal(pma_checker_OptimizationBarrier_15_io_y_pal),
    .io_y_paa(pma_checker_OptimizationBarrier_15_io_y_paa),
    .io_y_eff(pma_checker_OptimizationBarrier_15_io_y_eff),
    .io_y_c(pma_checker_OptimizationBarrier_15_io_y_c)
  );
  OptimizationBarrier pma_checker_OptimizationBarrier_16 ( // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178735.4]
    .io_x_ppn(pma_checker_OptimizationBarrier_16_io_x_ppn),
    .io_x_u(pma_checker_OptimizationBarrier_16_io_x_u),
    .io_x_ae(pma_checker_OptimizationBarrier_16_io_x_ae),
    .io_x_sw(pma_checker_OptimizationBarrier_16_io_x_sw),
    .io_x_sx(pma_checker_OptimizationBarrier_16_io_x_sx),
    .io_x_sr(pma_checker_OptimizationBarrier_16_io_x_sr),
    .io_x_pw(pma_checker_OptimizationBarrier_16_io_x_pw),
    .io_x_px(pma_checker_OptimizationBarrier_16_io_x_px),
    .io_x_pr(pma_checker_OptimizationBarrier_16_io_x_pr),
    .io_x_ppp(pma_checker_OptimizationBarrier_16_io_x_ppp),
    .io_x_pal(pma_checker_OptimizationBarrier_16_io_x_pal),
    .io_x_paa(pma_checker_OptimizationBarrier_16_io_x_paa),
    .io_x_eff(pma_checker_OptimizationBarrier_16_io_x_eff),
    .io_x_c(pma_checker_OptimizationBarrier_16_io_x_c),
    .io_y_ppn(pma_checker_OptimizationBarrier_16_io_y_ppn),
    .io_y_u(pma_checker_OptimizationBarrier_16_io_y_u),
    .io_y_ae(pma_checker_OptimizationBarrier_16_io_y_ae),
    .io_y_sw(pma_checker_OptimizationBarrier_16_io_y_sw),
    .io_y_sx(pma_checker_OptimizationBarrier_16_io_y_sx),
    .io_y_sr(pma_checker_OptimizationBarrier_16_io_y_sr),
    .io_y_pw(pma_checker_OptimizationBarrier_16_io_y_pw),
    .io_y_px(pma_checker_OptimizationBarrier_16_io_y_px),
    .io_y_pr(pma_checker_OptimizationBarrier_16_io_y_pr),
    .io_y_ppp(pma_checker_OptimizationBarrier_16_io_y_ppp),
    .io_y_pal(pma_checker_OptimizationBarrier_16_io_y_pal),
    .io_y_paa(pma_checker_OptimizationBarrier_16_io_y_paa),
    .io_y_eff(pma_checker_OptimizationBarrier_16_io_y_eff),
    .io_y_c(pma_checker_OptimizationBarrier_16_io_y_c)
  );
  OptimizationBarrier pma_checker_OptimizationBarrier_17 ( // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178778.4]
    .io_x_ppn(pma_checker_OptimizationBarrier_17_io_x_ppn),
    .io_x_u(pma_checker_OptimizationBarrier_17_io_x_u),
    .io_x_ae(pma_checker_OptimizationBarrier_17_io_x_ae),
    .io_x_sw(pma_checker_OptimizationBarrier_17_io_x_sw),
    .io_x_sx(pma_checker_OptimizationBarrier_17_io_x_sx),
    .io_x_sr(pma_checker_OptimizationBarrier_17_io_x_sr),
    .io_x_pw(pma_checker_OptimizationBarrier_17_io_x_pw),
    .io_x_px(pma_checker_OptimizationBarrier_17_io_x_px),
    .io_x_pr(pma_checker_OptimizationBarrier_17_io_x_pr),
    .io_x_ppp(pma_checker_OptimizationBarrier_17_io_x_ppp),
    .io_x_pal(pma_checker_OptimizationBarrier_17_io_x_pal),
    .io_x_paa(pma_checker_OptimizationBarrier_17_io_x_paa),
    .io_x_eff(pma_checker_OptimizationBarrier_17_io_x_eff),
    .io_x_c(pma_checker_OptimizationBarrier_17_io_x_c),
    .io_y_ppn(pma_checker_OptimizationBarrier_17_io_y_ppn),
    .io_y_u(pma_checker_OptimizationBarrier_17_io_y_u),
    .io_y_ae(pma_checker_OptimizationBarrier_17_io_y_ae),
    .io_y_sw(pma_checker_OptimizationBarrier_17_io_y_sw),
    .io_y_sx(pma_checker_OptimizationBarrier_17_io_y_sx),
    .io_y_sr(pma_checker_OptimizationBarrier_17_io_y_sr),
    .io_y_pw(pma_checker_OptimizationBarrier_17_io_y_pw),
    .io_y_px(pma_checker_OptimizationBarrier_17_io_y_px),
    .io_y_pr(pma_checker_OptimizationBarrier_17_io_y_pr),
    .io_y_ppp(pma_checker_OptimizationBarrier_17_io_y_ppp),
    .io_y_pal(pma_checker_OptimizationBarrier_17_io_y_pal),
    .io_y_paa(pma_checker_OptimizationBarrier_17_io_y_paa),
    .io_y_eff(pma_checker_OptimizationBarrier_17_io_y_eff),
    .io_y_c(pma_checker_OptimizationBarrier_17_io_y_c)
  );
  OptimizationBarrier pma_checker_OptimizationBarrier_18 ( // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178821.4]
    .io_x_ppn(pma_checker_OptimizationBarrier_18_io_x_ppn),
    .io_x_u(pma_checker_OptimizationBarrier_18_io_x_u),
    .io_x_ae(pma_checker_OptimizationBarrier_18_io_x_ae),
    .io_x_sw(pma_checker_OptimizationBarrier_18_io_x_sw),
    .io_x_sx(pma_checker_OptimizationBarrier_18_io_x_sx),
    .io_x_sr(pma_checker_OptimizationBarrier_18_io_x_sr),
    .io_x_pw(pma_checker_OptimizationBarrier_18_io_x_pw),
    .io_x_px(pma_checker_OptimizationBarrier_18_io_x_px),
    .io_x_pr(pma_checker_OptimizationBarrier_18_io_x_pr),
    .io_x_ppp(pma_checker_OptimizationBarrier_18_io_x_ppp),
    .io_x_pal(pma_checker_OptimizationBarrier_18_io_x_pal),
    .io_x_paa(pma_checker_OptimizationBarrier_18_io_x_paa),
    .io_x_eff(pma_checker_OptimizationBarrier_18_io_x_eff),
    .io_x_c(pma_checker_OptimizationBarrier_18_io_x_c),
    .io_y_ppn(pma_checker_OptimizationBarrier_18_io_y_ppn),
    .io_y_u(pma_checker_OptimizationBarrier_18_io_y_u),
    .io_y_ae(pma_checker_OptimizationBarrier_18_io_y_ae),
    .io_y_sw(pma_checker_OptimizationBarrier_18_io_y_sw),
    .io_y_sx(pma_checker_OptimizationBarrier_18_io_y_sx),
    .io_y_sr(pma_checker_OptimizationBarrier_18_io_y_sr),
    .io_y_pw(pma_checker_OptimizationBarrier_18_io_y_pw),
    .io_y_px(pma_checker_OptimizationBarrier_18_io_y_px),
    .io_y_pr(pma_checker_OptimizationBarrier_18_io_y_pr),
    .io_y_ppp(pma_checker_OptimizationBarrier_18_io_y_ppp),
    .io_y_pal(pma_checker_OptimizationBarrier_18_io_y_pal),
    .io_y_paa(pma_checker_OptimizationBarrier_18_io_y_paa),
    .io_y_eff(pma_checker_OptimizationBarrier_18_io_y_eff),
    .io_y_c(pma_checker_OptimizationBarrier_18_io_y_c)
  );
  OptimizationBarrier pma_checker_OptimizationBarrier_19 ( // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178864.4]
    .io_x_ppn(pma_checker_OptimizationBarrier_19_io_x_ppn),
    .io_x_u(pma_checker_OptimizationBarrier_19_io_x_u),
    .io_x_ae(pma_checker_OptimizationBarrier_19_io_x_ae),
    .io_x_sw(pma_checker_OptimizationBarrier_19_io_x_sw),
    .io_x_sx(pma_checker_OptimizationBarrier_19_io_x_sx),
    .io_x_sr(pma_checker_OptimizationBarrier_19_io_x_sr),
    .io_x_pw(pma_checker_OptimizationBarrier_19_io_x_pw),
    .io_x_px(pma_checker_OptimizationBarrier_19_io_x_px),
    .io_x_pr(pma_checker_OptimizationBarrier_19_io_x_pr),
    .io_x_ppp(pma_checker_OptimizationBarrier_19_io_x_ppp),
    .io_x_pal(pma_checker_OptimizationBarrier_19_io_x_pal),
    .io_x_paa(pma_checker_OptimizationBarrier_19_io_x_paa),
    .io_x_eff(pma_checker_OptimizationBarrier_19_io_x_eff),
    .io_x_c(pma_checker_OptimizationBarrier_19_io_x_c),
    .io_y_ppn(pma_checker_OptimizationBarrier_19_io_y_ppn),
    .io_y_u(pma_checker_OptimizationBarrier_19_io_y_u),
    .io_y_ae(pma_checker_OptimizationBarrier_19_io_y_ae),
    .io_y_sw(pma_checker_OptimizationBarrier_19_io_y_sw),
    .io_y_sx(pma_checker_OptimizationBarrier_19_io_y_sx),
    .io_y_sr(pma_checker_OptimizationBarrier_19_io_y_sr),
    .io_y_pw(pma_checker_OptimizationBarrier_19_io_y_pw),
    .io_y_px(pma_checker_OptimizationBarrier_19_io_y_px),
    .io_y_pr(pma_checker_OptimizationBarrier_19_io_y_pr),
    .io_y_ppp(pma_checker_OptimizationBarrier_19_io_y_ppp),
    .io_y_pal(pma_checker_OptimizationBarrier_19_io_y_pal),
    .io_y_paa(pma_checker_OptimizationBarrier_19_io_y_paa),
    .io_y_eff(pma_checker_OptimizationBarrier_19_io_y_eff),
    .io_y_c(pma_checker_OptimizationBarrier_19_io_y_c)
  );
  OptimizationBarrier pma_checker_OptimizationBarrier_20 ( // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178907.4]
    .io_x_ppn(pma_checker_OptimizationBarrier_20_io_x_ppn),
    .io_x_u(pma_checker_OptimizationBarrier_20_io_x_u),
    .io_x_ae(pma_checker_OptimizationBarrier_20_io_x_ae),
    .io_x_sw(pma_checker_OptimizationBarrier_20_io_x_sw),
    .io_x_sx(pma_checker_OptimizationBarrier_20_io_x_sx),
    .io_x_sr(pma_checker_OptimizationBarrier_20_io_x_sr),
    .io_x_pw(pma_checker_OptimizationBarrier_20_io_x_pw),
    .io_x_px(pma_checker_OptimizationBarrier_20_io_x_px),
    .io_x_pr(pma_checker_OptimizationBarrier_20_io_x_pr),
    .io_x_ppp(pma_checker_OptimizationBarrier_20_io_x_ppp),
    .io_x_pal(pma_checker_OptimizationBarrier_20_io_x_pal),
    .io_x_paa(pma_checker_OptimizationBarrier_20_io_x_paa),
    .io_x_eff(pma_checker_OptimizationBarrier_20_io_x_eff),
    .io_x_c(pma_checker_OptimizationBarrier_20_io_x_c),
    .io_y_ppn(pma_checker_OptimizationBarrier_20_io_y_ppn),
    .io_y_u(pma_checker_OptimizationBarrier_20_io_y_u),
    .io_y_ae(pma_checker_OptimizationBarrier_20_io_y_ae),
    .io_y_sw(pma_checker_OptimizationBarrier_20_io_y_sw),
    .io_y_sx(pma_checker_OptimizationBarrier_20_io_y_sx),
    .io_y_sr(pma_checker_OptimizationBarrier_20_io_y_sr),
    .io_y_pw(pma_checker_OptimizationBarrier_20_io_y_pw),
    .io_y_px(pma_checker_OptimizationBarrier_20_io_y_px),
    .io_y_pr(pma_checker_OptimizationBarrier_20_io_y_pr),
    .io_y_ppp(pma_checker_OptimizationBarrier_20_io_y_ppp),
    .io_y_pal(pma_checker_OptimizationBarrier_20_io_y_pal),
    .io_y_paa(pma_checker_OptimizationBarrier_20_io_y_paa),
    .io_y_eff(pma_checker_OptimizationBarrier_20_io_y_eff),
    .io_y_c(pma_checker_OptimizationBarrier_20_io_y_c)
  );
  OptimizationBarrier pma_checker_OptimizationBarrier_21 ( // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178950.4]
    .io_x_ppn(pma_checker_OptimizationBarrier_21_io_x_ppn),
    .io_x_u(pma_checker_OptimizationBarrier_21_io_x_u),
    .io_x_ae(pma_checker_OptimizationBarrier_21_io_x_ae),
    .io_x_sw(pma_checker_OptimizationBarrier_21_io_x_sw),
    .io_x_sx(pma_checker_OptimizationBarrier_21_io_x_sx),
    .io_x_sr(pma_checker_OptimizationBarrier_21_io_x_sr),
    .io_x_pw(pma_checker_OptimizationBarrier_21_io_x_pw),
    .io_x_px(pma_checker_OptimizationBarrier_21_io_x_px),
    .io_x_pr(pma_checker_OptimizationBarrier_21_io_x_pr),
    .io_x_ppp(pma_checker_OptimizationBarrier_21_io_x_ppp),
    .io_x_pal(pma_checker_OptimizationBarrier_21_io_x_pal),
    .io_x_paa(pma_checker_OptimizationBarrier_21_io_x_paa),
    .io_x_eff(pma_checker_OptimizationBarrier_21_io_x_eff),
    .io_x_c(pma_checker_OptimizationBarrier_21_io_x_c),
    .io_y_ppn(pma_checker_OptimizationBarrier_21_io_y_ppn),
    .io_y_u(pma_checker_OptimizationBarrier_21_io_y_u),
    .io_y_ae(pma_checker_OptimizationBarrier_21_io_y_ae),
    .io_y_sw(pma_checker_OptimizationBarrier_21_io_y_sw),
    .io_y_sx(pma_checker_OptimizationBarrier_21_io_y_sx),
    .io_y_sr(pma_checker_OptimizationBarrier_21_io_y_sr),
    .io_y_pw(pma_checker_OptimizationBarrier_21_io_y_pw),
    .io_y_px(pma_checker_OptimizationBarrier_21_io_y_px),
    .io_y_pr(pma_checker_OptimizationBarrier_21_io_y_pr),
    .io_y_ppp(pma_checker_OptimizationBarrier_21_io_y_ppp),
    .io_y_pal(pma_checker_OptimizationBarrier_21_io_y_pal),
    .io_y_paa(pma_checker_OptimizationBarrier_21_io_y_paa),
    .io_y_eff(pma_checker_OptimizationBarrier_21_io_y_eff),
    .io_y_c(pma_checker_OptimizationBarrier_21_io_y_c)
  );
  OptimizationBarrier pma_checker_OptimizationBarrier_22 ( // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@178992.4]
    .io_x_ppn(pma_checker_OptimizationBarrier_22_io_x_ppn),
    .io_x_u(pma_checker_OptimizationBarrier_22_io_x_u),
    .io_x_ae(pma_checker_OptimizationBarrier_22_io_x_ae),
    .io_x_sw(pma_checker_OptimizationBarrier_22_io_x_sw),
    .io_x_sx(pma_checker_OptimizationBarrier_22_io_x_sx),
    .io_x_sr(pma_checker_OptimizationBarrier_22_io_x_sr),
    .io_x_pw(pma_checker_OptimizationBarrier_22_io_x_pw),
    .io_x_px(pma_checker_OptimizationBarrier_22_io_x_px),
    .io_x_pr(pma_checker_OptimizationBarrier_22_io_x_pr),
    .io_x_ppp(pma_checker_OptimizationBarrier_22_io_x_ppp),
    .io_x_pal(pma_checker_OptimizationBarrier_22_io_x_pal),
    .io_x_paa(pma_checker_OptimizationBarrier_22_io_x_paa),
    .io_x_eff(pma_checker_OptimizationBarrier_22_io_x_eff),
    .io_x_c(pma_checker_OptimizationBarrier_22_io_x_c),
    .io_y_ppn(pma_checker_OptimizationBarrier_22_io_y_ppn),
    .io_y_u(pma_checker_OptimizationBarrier_22_io_y_u),
    .io_y_ae(pma_checker_OptimizationBarrier_22_io_y_ae),
    .io_y_sw(pma_checker_OptimizationBarrier_22_io_y_sw),
    .io_y_sx(pma_checker_OptimizationBarrier_22_io_y_sx),
    .io_y_sr(pma_checker_OptimizationBarrier_22_io_y_sr),
    .io_y_pw(pma_checker_OptimizationBarrier_22_io_y_pw),
    .io_y_px(pma_checker_OptimizationBarrier_22_io_y_px),
    .io_y_pr(pma_checker_OptimizationBarrier_22_io_y_pr),
    .io_y_ppp(pma_checker_OptimizationBarrier_22_io_y_ppp),
    .io_y_pal(pma_checker_OptimizationBarrier_22_io_y_pal),
    .io_y_paa(pma_checker_OptimizationBarrier_22_io_y_paa),
    .io_y_eff(pma_checker_OptimizationBarrier_22_io_y_eff),
    .io_y_c(pma_checker_OptimizationBarrier_22_io_y_c)
  );
  OptimizationBarrier pma_checker_OptimizationBarrier_23 ( // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179034.4]
    .io_x_ppn(pma_checker_OptimizationBarrier_23_io_x_ppn),
    .io_x_u(pma_checker_OptimizationBarrier_23_io_x_u),
    .io_x_ae(pma_checker_OptimizationBarrier_23_io_x_ae),
    .io_x_sw(pma_checker_OptimizationBarrier_23_io_x_sw),
    .io_x_sx(pma_checker_OptimizationBarrier_23_io_x_sx),
    .io_x_sr(pma_checker_OptimizationBarrier_23_io_x_sr),
    .io_x_pw(pma_checker_OptimizationBarrier_23_io_x_pw),
    .io_x_px(pma_checker_OptimizationBarrier_23_io_x_px),
    .io_x_pr(pma_checker_OptimizationBarrier_23_io_x_pr),
    .io_x_ppp(pma_checker_OptimizationBarrier_23_io_x_ppp),
    .io_x_pal(pma_checker_OptimizationBarrier_23_io_x_pal),
    .io_x_paa(pma_checker_OptimizationBarrier_23_io_x_paa),
    .io_x_eff(pma_checker_OptimizationBarrier_23_io_x_eff),
    .io_x_c(pma_checker_OptimizationBarrier_23_io_x_c),
    .io_y_ppn(pma_checker_OptimizationBarrier_23_io_y_ppn),
    .io_y_u(pma_checker_OptimizationBarrier_23_io_y_u),
    .io_y_ae(pma_checker_OptimizationBarrier_23_io_y_ae),
    .io_y_sw(pma_checker_OptimizationBarrier_23_io_y_sw),
    .io_y_sx(pma_checker_OptimizationBarrier_23_io_y_sx),
    .io_y_sr(pma_checker_OptimizationBarrier_23_io_y_sr),
    .io_y_pw(pma_checker_OptimizationBarrier_23_io_y_pw),
    .io_y_px(pma_checker_OptimizationBarrier_23_io_y_px),
    .io_y_pr(pma_checker_OptimizationBarrier_23_io_y_pr),
    .io_y_ppp(pma_checker_OptimizationBarrier_23_io_y_ppp),
    .io_y_pal(pma_checker_OptimizationBarrier_23_io_y_pal),
    .io_y_paa(pma_checker_OptimizationBarrier_23_io_y_paa),
    .io_y_eff(pma_checker_OptimizationBarrier_23_io_y_eff),
    .io_y_c(pma_checker_OptimizationBarrier_23_io_y_c)
  );
  OptimizationBarrier pma_checker_OptimizationBarrier_24 ( // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179076.4]
    .io_x_ppn(pma_checker_OptimizationBarrier_24_io_x_ppn),
    .io_x_u(pma_checker_OptimizationBarrier_24_io_x_u),
    .io_x_ae(pma_checker_OptimizationBarrier_24_io_x_ae),
    .io_x_sw(pma_checker_OptimizationBarrier_24_io_x_sw),
    .io_x_sx(pma_checker_OptimizationBarrier_24_io_x_sx),
    .io_x_sr(pma_checker_OptimizationBarrier_24_io_x_sr),
    .io_x_pw(pma_checker_OptimizationBarrier_24_io_x_pw),
    .io_x_px(pma_checker_OptimizationBarrier_24_io_x_px),
    .io_x_pr(pma_checker_OptimizationBarrier_24_io_x_pr),
    .io_x_ppp(pma_checker_OptimizationBarrier_24_io_x_ppp),
    .io_x_pal(pma_checker_OptimizationBarrier_24_io_x_pal),
    .io_x_paa(pma_checker_OptimizationBarrier_24_io_x_paa),
    .io_x_eff(pma_checker_OptimizationBarrier_24_io_x_eff),
    .io_x_c(pma_checker_OptimizationBarrier_24_io_x_c),
    .io_y_ppn(pma_checker_OptimizationBarrier_24_io_y_ppn),
    .io_y_u(pma_checker_OptimizationBarrier_24_io_y_u),
    .io_y_ae(pma_checker_OptimizationBarrier_24_io_y_ae),
    .io_y_sw(pma_checker_OptimizationBarrier_24_io_y_sw),
    .io_y_sx(pma_checker_OptimizationBarrier_24_io_y_sx),
    .io_y_sr(pma_checker_OptimizationBarrier_24_io_y_sr),
    .io_y_pw(pma_checker_OptimizationBarrier_24_io_y_pw),
    .io_y_px(pma_checker_OptimizationBarrier_24_io_y_px),
    .io_y_pr(pma_checker_OptimizationBarrier_24_io_y_pr),
    .io_y_ppp(pma_checker_OptimizationBarrier_24_io_y_ppp),
    .io_y_pal(pma_checker_OptimizationBarrier_24_io_y_pal),
    .io_y_paa(pma_checker_OptimizationBarrier_24_io_y_paa),
    .io_y_eff(pma_checker_OptimizationBarrier_24_io_y_eff),
    .io_y_c(pma_checker_OptimizationBarrier_24_io_y_c)
  );
  OptimizationBarrier pma_checker_OptimizationBarrier_25 ( // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179118.4]
    .io_x_ppn(pma_checker_OptimizationBarrier_25_io_x_ppn),
    .io_x_u(pma_checker_OptimizationBarrier_25_io_x_u),
    .io_x_ae(pma_checker_OptimizationBarrier_25_io_x_ae),
    .io_x_sw(pma_checker_OptimizationBarrier_25_io_x_sw),
    .io_x_sx(pma_checker_OptimizationBarrier_25_io_x_sx),
    .io_x_sr(pma_checker_OptimizationBarrier_25_io_x_sr),
    .io_x_pw(pma_checker_OptimizationBarrier_25_io_x_pw),
    .io_x_px(pma_checker_OptimizationBarrier_25_io_x_px),
    .io_x_pr(pma_checker_OptimizationBarrier_25_io_x_pr),
    .io_x_ppp(pma_checker_OptimizationBarrier_25_io_x_ppp),
    .io_x_pal(pma_checker_OptimizationBarrier_25_io_x_pal),
    .io_x_paa(pma_checker_OptimizationBarrier_25_io_x_paa),
    .io_x_eff(pma_checker_OptimizationBarrier_25_io_x_eff),
    .io_x_c(pma_checker_OptimizationBarrier_25_io_x_c),
    .io_y_ppn(pma_checker_OptimizationBarrier_25_io_y_ppn),
    .io_y_u(pma_checker_OptimizationBarrier_25_io_y_u),
    .io_y_ae(pma_checker_OptimizationBarrier_25_io_y_ae),
    .io_y_sw(pma_checker_OptimizationBarrier_25_io_y_sw),
    .io_y_sx(pma_checker_OptimizationBarrier_25_io_y_sx),
    .io_y_sr(pma_checker_OptimizationBarrier_25_io_y_sr),
    .io_y_pw(pma_checker_OptimizationBarrier_25_io_y_pw),
    .io_y_px(pma_checker_OptimizationBarrier_25_io_y_px),
    .io_y_pr(pma_checker_OptimizationBarrier_25_io_y_pr),
    .io_y_ppp(pma_checker_OptimizationBarrier_25_io_y_ppp),
    .io_y_pal(pma_checker_OptimizationBarrier_25_io_y_pal),
    .io_y_paa(pma_checker_OptimizationBarrier_25_io_y_paa),
    .io_y_eff(pma_checker_OptimizationBarrier_25_io_y_eff),
    .io_y_c(pma_checker_OptimizationBarrier_25_io_y_c)
  );
  OptimizationBarrier pma_checker_OptimizationBarrier_26 ( // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179160.4]
    .io_x_ppn(pma_checker_OptimizationBarrier_26_io_x_ppn),
    .io_x_u(pma_checker_OptimizationBarrier_26_io_x_u),
    .io_x_ae(pma_checker_OptimizationBarrier_26_io_x_ae),
    .io_x_sw(pma_checker_OptimizationBarrier_26_io_x_sw),
    .io_x_sx(pma_checker_OptimizationBarrier_26_io_x_sx),
    .io_x_sr(pma_checker_OptimizationBarrier_26_io_x_sr),
    .io_x_pw(pma_checker_OptimizationBarrier_26_io_x_pw),
    .io_x_px(pma_checker_OptimizationBarrier_26_io_x_px),
    .io_x_pr(pma_checker_OptimizationBarrier_26_io_x_pr),
    .io_x_ppp(pma_checker_OptimizationBarrier_26_io_x_ppp),
    .io_x_pal(pma_checker_OptimizationBarrier_26_io_x_pal),
    .io_x_paa(pma_checker_OptimizationBarrier_26_io_x_paa),
    .io_x_eff(pma_checker_OptimizationBarrier_26_io_x_eff),
    .io_x_c(pma_checker_OptimizationBarrier_26_io_x_c),
    .io_y_ppn(pma_checker_OptimizationBarrier_26_io_y_ppn),
    .io_y_u(pma_checker_OptimizationBarrier_26_io_y_u),
    .io_y_ae(pma_checker_OptimizationBarrier_26_io_y_ae),
    .io_y_sw(pma_checker_OptimizationBarrier_26_io_y_sw),
    .io_y_sx(pma_checker_OptimizationBarrier_26_io_y_sx),
    .io_y_sr(pma_checker_OptimizationBarrier_26_io_y_sr),
    .io_y_pw(pma_checker_OptimizationBarrier_26_io_y_pw),
    .io_y_px(pma_checker_OptimizationBarrier_26_io_y_px),
    .io_y_pr(pma_checker_OptimizationBarrier_26_io_y_pr),
    .io_y_ppp(pma_checker_OptimizationBarrier_26_io_y_ppp),
    .io_y_pal(pma_checker_OptimizationBarrier_26_io_y_pal),
    .io_y_paa(pma_checker_OptimizationBarrier_26_io_y_paa),
    .io_y_eff(pma_checker_OptimizationBarrier_26_io_y_eff),
    .io_y_c(pma_checker_OptimizationBarrier_26_io_y_c)
  );
  OptimizationBarrier pma_checker_OptimizationBarrier_27 ( // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179203.4]
    .io_x_ppn(pma_checker_OptimizationBarrier_27_io_x_ppn),
    .io_x_u(pma_checker_OptimizationBarrier_27_io_x_u),
    .io_x_ae(pma_checker_OptimizationBarrier_27_io_x_ae),
    .io_x_sw(pma_checker_OptimizationBarrier_27_io_x_sw),
    .io_x_sx(pma_checker_OptimizationBarrier_27_io_x_sx),
    .io_x_sr(pma_checker_OptimizationBarrier_27_io_x_sr),
    .io_x_pw(pma_checker_OptimizationBarrier_27_io_x_pw),
    .io_x_px(pma_checker_OptimizationBarrier_27_io_x_px),
    .io_x_pr(pma_checker_OptimizationBarrier_27_io_x_pr),
    .io_x_ppp(pma_checker_OptimizationBarrier_27_io_x_ppp),
    .io_x_pal(pma_checker_OptimizationBarrier_27_io_x_pal),
    .io_x_paa(pma_checker_OptimizationBarrier_27_io_x_paa),
    .io_x_eff(pma_checker_OptimizationBarrier_27_io_x_eff),
    .io_x_c(pma_checker_OptimizationBarrier_27_io_x_c),
    .io_y_ppn(pma_checker_OptimizationBarrier_27_io_y_ppn),
    .io_y_u(pma_checker_OptimizationBarrier_27_io_y_u),
    .io_y_ae(pma_checker_OptimizationBarrier_27_io_y_ae),
    .io_y_sw(pma_checker_OptimizationBarrier_27_io_y_sw),
    .io_y_sx(pma_checker_OptimizationBarrier_27_io_y_sx),
    .io_y_sr(pma_checker_OptimizationBarrier_27_io_y_sr),
    .io_y_pw(pma_checker_OptimizationBarrier_27_io_y_pw),
    .io_y_px(pma_checker_OptimizationBarrier_27_io_y_px),
    .io_y_pr(pma_checker_OptimizationBarrier_27_io_y_pr),
    .io_y_ppp(pma_checker_OptimizationBarrier_27_io_y_ppp),
    .io_y_pal(pma_checker_OptimizationBarrier_27_io_y_pal),
    .io_y_paa(pma_checker_OptimizationBarrier_27_io_y_paa),
    .io_y_eff(pma_checker_OptimizationBarrier_27_io_y_eff),
    .io_y_c(pma_checker_OptimizationBarrier_27_io_y_c)
  );
  OptimizationBarrier pma_checker_OptimizationBarrier_28 ( // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179246.4]
    .io_x_ppn(pma_checker_OptimizationBarrier_28_io_x_ppn),
    .io_x_u(pma_checker_OptimizationBarrier_28_io_x_u),
    .io_x_ae(pma_checker_OptimizationBarrier_28_io_x_ae),
    .io_x_sw(pma_checker_OptimizationBarrier_28_io_x_sw),
    .io_x_sx(pma_checker_OptimizationBarrier_28_io_x_sx),
    .io_x_sr(pma_checker_OptimizationBarrier_28_io_x_sr),
    .io_x_pw(pma_checker_OptimizationBarrier_28_io_x_pw),
    .io_x_px(pma_checker_OptimizationBarrier_28_io_x_px),
    .io_x_pr(pma_checker_OptimizationBarrier_28_io_x_pr),
    .io_x_ppp(pma_checker_OptimizationBarrier_28_io_x_ppp),
    .io_x_pal(pma_checker_OptimizationBarrier_28_io_x_pal),
    .io_x_paa(pma_checker_OptimizationBarrier_28_io_x_paa),
    .io_x_eff(pma_checker_OptimizationBarrier_28_io_x_eff),
    .io_x_c(pma_checker_OptimizationBarrier_28_io_x_c),
    .io_y_ppn(pma_checker_OptimizationBarrier_28_io_y_ppn),
    .io_y_u(pma_checker_OptimizationBarrier_28_io_y_u),
    .io_y_ae(pma_checker_OptimizationBarrier_28_io_y_ae),
    .io_y_sw(pma_checker_OptimizationBarrier_28_io_y_sw),
    .io_y_sx(pma_checker_OptimizationBarrier_28_io_y_sx),
    .io_y_sr(pma_checker_OptimizationBarrier_28_io_y_sr),
    .io_y_pw(pma_checker_OptimizationBarrier_28_io_y_pw),
    .io_y_px(pma_checker_OptimizationBarrier_28_io_y_px),
    .io_y_pr(pma_checker_OptimizationBarrier_28_io_y_pr),
    .io_y_ppp(pma_checker_OptimizationBarrier_28_io_y_ppp),
    .io_y_pal(pma_checker_OptimizationBarrier_28_io_y_pal),
    .io_y_paa(pma_checker_OptimizationBarrier_28_io_y_paa),
    .io_y_eff(pma_checker_OptimizationBarrier_28_io_y_eff),
    .io_y_c(pma_checker_OptimizationBarrier_28_io_y_c)
  );
  OptimizationBarrier pma_checker_OptimizationBarrier_29 ( // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179289.4]
    .io_x_ppn(pma_checker_OptimizationBarrier_29_io_x_ppn),
    .io_x_u(pma_checker_OptimizationBarrier_29_io_x_u),
    .io_x_ae(pma_checker_OptimizationBarrier_29_io_x_ae),
    .io_x_sw(pma_checker_OptimizationBarrier_29_io_x_sw),
    .io_x_sx(pma_checker_OptimizationBarrier_29_io_x_sx),
    .io_x_sr(pma_checker_OptimizationBarrier_29_io_x_sr),
    .io_x_pw(pma_checker_OptimizationBarrier_29_io_x_pw),
    .io_x_px(pma_checker_OptimizationBarrier_29_io_x_px),
    .io_x_pr(pma_checker_OptimizationBarrier_29_io_x_pr),
    .io_x_ppp(pma_checker_OptimizationBarrier_29_io_x_ppp),
    .io_x_pal(pma_checker_OptimizationBarrier_29_io_x_pal),
    .io_x_paa(pma_checker_OptimizationBarrier_29_io_x_paa),
    .io_x_eff(pma_checker_OptimizationBarrier_29_io_x_eff),
    .io_x_c(pma_checker_OptimizationBarrier_29_io_x_c),
    .io_y_ppn(pma_checker_OptimizationBarrier_29_io_y_ppn),
    .io_y_u(pma_checker_OptimizationBarrier_29_io_y_u),
    .io_y_ae(pma_checker_OptimizationBarrier_29_io_y_ae),
    .io_y_sw(pma_checker_OptimizationBarrier_29_io_y_sw),
    .io_y_sx(pma_checker_OptimizationBarrier_29_io_y_sx),
    .io_y_sr(pma_checker_OptimizationBarrier_29_io_y_sr),
    .io_y_pw(pma_checker_OptimizationBarrier_29_io_y_pw),
    .io_y_px(pma_checker_OptimizationBarrier_29_io_y_px),
    .io_y_pr(pma_checker_OptimizationBarrier_29_io_y_pr),
    .io_y_ppp(pma_checker_OptimizationBarrier_29_io_y_ppp),
    .io_y_pal(pma_checker_OptimizationBarrier_29_io_y_pal),
    .io_y_paa(pma_checker_OptimizationBarrier_29_io_y_paa),
    .io_y_eff(pma_checker_OptimizationBarrier_29_io_y_eff),
    .io_y_c(pma_checker_OptimizationBarrier_29_io_y_c)
  );
  OptimizationBarrier pma_checker_OptimizationBarrier_30 ( // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179332.4]
    .io_x_ppn(pma_checker_OptimizationBarrier_30_io_x_ppn),
    .io_x_u(pma_checker_OptimizationBarrier_30_io_x_u),
    .io_x_ae(pma_checker_OptimizationBarrier_30_io_x_ae),
    .io_x_sw(pma_checker_OptimizationBarrier_30_io_x_sw),
    .io_x_sx(pma_checker_OptimizationBarrier_30_io_x_sx),
    .io_x_sr(pma_checker_OptimizationBarrier_30_io_x_sr),
    .io_x_pw(pma_checker_OptimizationBarrier_30_io_x_pw),
    .io_x_px(pma_checker_OptimizationBarrier_30_io_x_px),
    .io_x_pr(pma_checker_OptimizationBarrier_30_io_x_pr),
    .io_x_ppp(pma_checker_OptimizationBarrier_30_io_x_ppp),
    .io_x_pal(pma_checker_OptimizationBarrier_30_io_x_pal),
    .io_x_paa(pma_checker_OptimizationBarrier_30_io_x_paa),
    .io_x_eff(pma_checker_OptimizationBarrier_30_io_x_eff),
    .io_x_c(pma_checker_OptimizationBarrier_30_io_x_c),
    .io_y_ppn(pma_checker_OptimizationBarrier_30_io_y_ppn),
    .io_y_u(pma_checker_OptimizationBarrier_30_io_y_u),
    .io_y_ae(pma_checker_OptimizationBarrier_30_io_y_ae),
    .io_y_sw(pma_checker_OptimizationBarrier_30_io_y_sw),
    .io_y_sx(pma_checker_OptimizationBarrier_30_io_y_sx),
    .io_y_sr(pma_checker_OptimizationBarrier_30_io_y_sr),
    .io_y_pw(pma_checker_OptimizationBarrier_30_io_y_pw),
    .io_y_px(pma_checker_OptimizationBarrier_30_io_y_px),
    .io_y_pr(pma_checker_OptimizationBarrier_30_io_y_pr),
    .io_y_ppp(pma_checker_OptimizationBarrier_30_io_y_ppp),
    .io_y_pal(pma_checker_OptimizationBarrier_30_io_y_pal),
    .io_y_paa(pma_checker_OptimizationBarrier_30_io_y_paa),
    .io_y_eff(pma_checker_OptimizationBarrier_30_io_y_eff),
    .io_y_c(pma_checker_OptimizationBarrier_30_io_y_c)
  );
  OptimizationBarrier pma_checker_OptimizationBarrier_31 ( // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179375.4]
    .io_x_ppn(pma_checker_OptimizationBarrier_31_io_x_ppn),
    .io_x_u(pma_checker_OptimizationBarrier_31_io_x_u),
    .io_x_ae(pma_checker_OptimizationBarrier_31_io_x_ae),
    .io_x_sw(pma_checker_OptimizationBarrier_31_io_x_sw),
    .io_x_sx(pma_checker_OptimizationBarrier_31_io_x_sx),
    .io_x_sr(pma_checker_OptimizationBarrier_31_io_x_sr),
    .io_x_pw(pma_checker_OptimizationBarrier_31_io_x_pw),
    .io_x_px(pma_checker_OptimizationBarrier_31_io_x_px),
    .io_x_pr(pma_checker_OptimizationBarrier_31_io_x_pr),
    .io_x_ppp(pma_checker_OptimizationBarrier_31_io_x_ppp),
    .io_x_pal(pma_checker_OptimizationBarrier_31_io_x_pal),
    .io_x_paa(pma_checker_OptimizationBarrier_31_io_x_paa),
    .io_x_eff(pma_checker_OptimizationBarrier_31_io_x_eff),
    .io_x_c(pma_checker_OptimizationBarrier_31_io_x_c),
    .io_y_ppn(pma_checker_OptimizationBarrier_31_io_y_ppn),
    .io_y_u(pma_checker_OptimizationBarrier_31_io_y_u),
    .io_y_ae(pma_checker_OptimizationBarrier_31_io_y_ae),
    .io_y_sw(pma_checker_OptimizationBarrier_31_io_y_sw),
    .io_y_sx(pma_checker_OptimizationBarrier_31_io_y_sx),
    .io_y_sr(pma_checker_OptimizationBarrier_31_io_y_sr),
    .io_y_pw(pma_checker_OptimizationBarrier_31_io_y_pw),
    .io_y_px(pma_checker_OptimizationBarrier_31_io_y_px),
    .io_y_pr(pma_checker_OptimizationBarrier_31_io_y_pr),
    .io_y_ppp(pma_checker_OptimizationBarrier_31_io_y_ppp),
    .io_y_pal(pma_checker_OptimizationBarrier_31_io_y_pal),
    .io_y_paa(pma_checker_OptimizationBarrier_31_io_y_paa),
    .io_y_eff(pma_checker_OptimizationBarrier_31_io_y_eff),
    .io_y_c(pma_checker_OptimizationBarrier_31_io_y_c)
  );
  OptimizationBarrier pma_checker_OptimizationBarrier_32 ( // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179418.4]
    .io_x_ppn(pma_checker_OptimizationBarrier_32_io_x_ppn),
    .io_x_u(pma_checker_OptimizationBarrier_32_io_x_u),
    .io_x_ae(pma_checker_OptimizationBarrier_32_io_x_ae),
    .io_x_sw(pma_checker_OptimizationBarrier_32_io_x_sw),
    .io_x_sx(pma_checker_OptimizationBarrier_32_io_x_sx),
    .io_x_sr(pma_checker_OptimizationBarrier_32_io_x_sr),
    .io_x_pw(pma_checker_OptimizationBarrier_32_io_x_pw),
    .io_x_px(pma_checker_OptimizationBarrier_32_io_x_px),
    .io_x_pr(pma_checker_OptimizationBarrier_32_io_x_pr),
    .io_x_ppp(pma_checker_OptimizationBarrier_32_io_x_ppp),
    .io_x_pal(pma_checker_OptimizationBarrier_32_io_x_pal),
    .io_x_paa(pma_checker_OptimizationBarrier_32_io_x_paa),
    .io_x_eff(pma_checker_OptimizationBarrier_32_io_x_eff),
    .io_x_c(pma_checker_OptimizationBarrier_32_io_x_c),
    .io_y_ppn(pma_checker_OptimizationBarrier_32_io_y_ppn),
    .io_y_u(pma_checker_OptimizationBarrier_32_io_y_u),
    .io_y_ae(pma_checker_OptimizationBarrier_32_io_y_ae),
    .io_y_sw(pma_checker_OptimizationBarrier_32_io_y_sw),
    .io_y_sx(pma_checker_OptimizationBarrier_32_io_y_sx),
    .io_y_sr(pma_checker_OptimizationBarrier_32_io_y_sr),
    .io_y_pw(pma_checker_OptimizationBarrier_32_io_y_pw),
    .io_y_px(pma_checker_OptimizationBarrier_32_io_y_px),
    .io_y_pr(pma_checker_OptimizationBarrier_32_io_y_pr),
    .io_y_ppp(pma_checker_OptimizationBarrier_32_io_y_ppp),
    .io_y_pal(pma_checker_OptimizationBarrier_32_io_y_pal),
    .io_y_paa(pma_checker_OptimizationBarrier_32_io_y_paa),
    .io_y_eff(pma_checker_OptimizationBarrier_32_io_y_eff),
    .io_y_c(pma_checker_OptimizationBarrier_32_io_y_c)
  );
  OptimizationBarrier pma_checker_OptimizationBarrier_33 ( // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179461.4]
    .io_x_ppn(pma_checker_OptimizationBarrier_33_io_x_ppn),
    .io_x_u(pma_checker_OptimizationBarrier_33_io_x_u),
    .io_x_ae(pma_checker_OptimizationBarrier_33_io_x_ae),
    .io_x_sw(pma_checker_OptimizationBarrier_33_io_x_sw),
    .io_x_sx(pma_checker_OptimizationBarrier_33_io_x_sx),
    .io_x_sr(pma_checker_OptimizationBarrier_33_io_x_sr),
    .io_x_pw(pma_checker_OptimizationBarrier_33_io_x_pw),
    .io_x_px(pma_checker_OptimizationBarrier_33_io_x_px),
    .io_x_pr(pma_checker_OptimizationBarrier_33_io_x_pr),
    .io_x_ppp(pma_checker_OptimizationBarrier_33_io_x_ppp),
    .io_x_pal(pma_checker_OptimizationBarrier_33_io_x_pal),
    .io_x_paa(pma_checker_OptimizationBarrier_33_io_x_paa),
    .io_x_eff(pma_checker_OptimizationBarrier_33_io_x_eff),
    .io_x_c(pma_checker_OptimizationBarrier_33_io_x_c),
    .io_y_ppn(pma_checker_OptimizationBarrier_33_io_y_ppn),
    .io_y_u(pma_checker_OptimizationBarrier_33_io_y_u),
    .io_y_ae(pma_checker_OptimizationBarrier_33_io_y_ae),
    .io_y_sw(pma_checker_OptimizationBarrier_33_io_y_sw),
    .io_y_sx(pma_checker_OptimizationBarrier_33_io_y_sx),
    .io_y_sr(pma_checker_OptimizationBarrier_33_io_y_sr),
    .io_y_pw(pma_checker_OptimizationBarrier_33_io_y_pw),
    .io_y_px(pma_checker_OptimizationBarrier_33_io_y_px),
    .io_y_pr(pma_checker_OptimizationBarrier_33_io_y_pr),
    .io_y_ppp(pma_checker_OptimizationBarrier_33_io_y_ppp),
    .io_y_pal(pma_checker_OptimizationBarrier_33_io_y_pal),
    .io_y_paa(pma_checker_OptimizationBarrier_33_io_y_paa),
    .io_y_eff(pma_checker_OptimizationBarrier_33_io_y_eff),
    .io_y_c(pma_checker_OptimizationBarrier_33_io_y_c)
  );
  OptimizationBarrier pma_checker_OptimizationBarrier_34 ( // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179504.4]
    .io_x_ppn(pma_checker_OptimizationBarrier_34_io_x_ppn),
    .io_x_u(pma_checker_OptimizationBarrier_34_io_x_u),
    .io_x_ae(pma_checker_OptimizationBarrier_34_io_x_ae),
    .io_x_sw(pma_checker_OptimizationBarrier_34_io_x_sw),
    .io_x_sx(pma_checker_OptimizationBarrier_34_io_x_sx),
    .io_x_sr(pma_checker_OptimizationBarrier_34_io_x_sr),
    .io_x_pw(pma_checker_OptimizationBarrier_34_io_x_pw),
    .io_x_px(pma_checker_OptimizationBarrier_34_io_x_px),
    .io_x_pr(pma_checker_OptimizationBarrier_34_io_x_pr),
    .io_x_ppp(pma_checker_OptimizationBarrier_34_io_x_ppp),
    .io_x_pal(pma_checker_OptimizationBarrier_34_io_x_pal),
    .io_x_paa(pma_checker_OptimizationBarrier_34_io_x_paa),
    .io_x_eff(pma_checker_OptimizationBarrier_34_io_x_eff),
    .io_x_c(pma_checker_OptimizationBarrier_34_io_x_c),
    .io_y_ppn(pma_checker_OptimizationBarrier_34_io_y_ppn),
    .io_y_u(pma_checker_OptimizationBarrier_34_io_y_u),
    .io_y_ae(pma_checker_OptimizationBarrier_34_io_y_ae),
    .io_y_sw(pma_checker_OptimizationBarrier_34_io_y_sw),
    .io_y_sx(pma_checker_OptimizationBarrier_34_io_y_sx),
    .io_y_sr(pma_checker_OptimizationBarrier_34_io_y_sr),
    .io_y_pw(pma_checker_OptimizationBarrier_34_io_y_pw),
    .io_y_px(pma_checker_OptimizationBarrier_34_io_y_px),
    .io_y_pr(pma_checker_OptimizationBarrier_34_io_y_pr),
    .io_y_ppp(pma_checker_OptimizationBarrier_34_io_y_ppp),
    .io_y_pal(pma_checker_OptimizationBarrier_34_io_y_pal),
    .io_y_paa(pma_checker_OptimizationBarrier_34_io_y_paa),
    .io_y_eff(pma_checker_OptimizationBarrier_34_io_y_eff),
    .io_y_c(pma_checker_OptimizationBarrier_34_io_y_c)
  );
  OptimizationBarrier pma_checker_OptimizationBarrier_35 ( // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179546.4]
    .io_x_ppn(pma_checker_OptimizationBarrier_35_io_x_ppn),
    .io_x_u(pma_checker_OptimizationBarrier_35_io_x_u),
    .io_x_ae(pma_checker_OptimizationBarrier_35_io_x_ae),
    .io_x_sw(pma_checker_OptimizationBarrier_35_io_x_sw),
    .io_x_sx(pma_checker_OptimizationBarrier_35_io_x_sx),
    .io_x_sr(pma_checker_OptimizationBarrier_35_io_x_sr),
    .io_x_pw(pma_checker_OptimizationBarrier_35_io_x_pw),
    .io_x_px(pma_checker_OptimizationBarrier_35_io_x_px),
    .io_x_pr(pma_checker_OptimizationBarrier_35_io_x_pr),
    .io_x_ppp(pma_checker_OptimizationBarrier_35_io_x_ppp),
    .io_x_pal(pma_checker_OptimizationBarrier_35_io_x_pal),
    .io_x_paa(pma_checker_OptimizationBarrier_35_io_x_paa),
    .io_x_eff(pma_checker_OptimizationBarrier_35_io_x_eff),
    .io_x_c(pma_checker_OptimizationBarrier_35_io_x_c),
    .io_y_ppn(pma_checker_OptimizationBarrier_35_io_y_ppn),
    .io_y_u(pma_checker_OptimizationBarrier_35_io_y_u),
    .io_y_ae(pma_checker_OptimizationBarrier_35_io_y_ae),
    .io_y_sw(pma_checker_OptimizationBarrier_35_io_y_sw),
    .io_y_sx(pma_checker_OptimizationBarrier_35_io_y_sx),
    .io_y_sr(pma_checker_OptimizationBarrier_35_io_y_sr),
    .io_y_pw(pma_checker_OptimizationBarrier_35_io_y_pw),
    .io_y_px(pma_checker_OptimizationBarrier_35_io_y_px),
    .io_y_pr(pma_checker_OptimizationBarrier_35_io_y_pr),
    .io_y_ppp(pma_checker_OptimizationBarrier_35_io_y_ppp),
    .io_y_pal(pma_checker_OptimizationBarrier_35_io_y_pal),
    .io_y_paa(pma_checker_OptimizationBarrier_35_io_y_paa),
    .io_y_eff(pma_checker_OptimizationBarrier_35_io_y_eff),
    .io_y_c(pma_checker_OptimizationBarrier_35_io_y_c)
  );
  OptimizationBarrier pma_checker_OptimizationBarrier_36 ( // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179588.4]
    .io_x_ppn(pma_checker_OptimizationBarrier_36_io_x_ppn),
    .io_x_u(pma_checker_OptimizationBarrier_36_io_x_u),
    .io_x_ae(pma_checker_OptimizationBarrier_36_io_x_ae),
    .io_x_sw(pma_checker_OptimizationBarrier_36_io_x_sw),
    .io_x_sx(pma_checker_OptimizationBarrier_36_io_x_sx),
    .io_x_sr(pma_checker_OptimizationBarrier_36_io_x_sr),
    .io_x_pw(pma_checker_OptimizationBarrier_36_io_x_pw),
    .io_x_px(pma_checker_OptimizationBarrier_36_io_x_px),
    .io_x_pr(pma_checker_OptimizationBarrier_36_io_x_pr),
    .io_x_ppp(pma_checker_OptimizationBarrier_36_io_x_ppp),
    .io_x_pal(pma_checker_OptimizationBarrier_36_io_x_pal),
    .io_x_paa(pma_checker_OptimizationBarrier_36_io_x_paa),
    .io_x_eff(pma_checker_OptimizationBarrier_36_io_x_eff),
    .io_x_c(pma_checker_OptimizationBarrier_36_io_x_c),
    .io_y_ppn(pma_checker_OptimizationBarrier_36_io_y_ppn),
    .io_y_u(pma_checker_OptimizationBarrier_36_io_y_u),
    .io_y_ae(pma_checker_OptimizationBarrier_36_io_y_ae),
    .io_y_sw(pma_checker_OptimizationBarrier_36_io_y_sw),
    .io_y_sx(pma_checker_OptimizationBarrier_36_io_y_sx),
    .io_y_sr(pma_checker_OptimizationBarrier_36_io_y_sr),
    .io_y_pw(pma_checker_OptimizationBarrier_36_io_y_pw),
    .io_y_px(pma_checker_OptimizationBarrier_36_io_y_px),
    .io_y_pr(pma_checker_OptimizationBarrier_36_io_y_pr),
    .io_y_ppp(pma_checker_OptimizationBarrier_36_io_y_ppp),
    .io_y_pal(pma_checker_OptimizationBarrier_36_io_y_pal),
    .io_y_paa(pma_checker_OptimizationBarrier_36_io_y_paa),
    .io_y_eff(pma_checker_OptimizationBarrier_36_io_y_eff),
    .io_y_c(pma_checker_OptimizationBarrier_36_io_y_c)
  );
  OptimizationBarrier pma_checker_OptimizationBarrier_37 ( // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179630.4]
    .io_x_ppn(pma_checker_OptimizationBarrier_37_io_x_ppn),
    .io_x_u(pma_checker_OptimizationBarrier_37_io_x_u),
    .io_x_ae(pma_checker_OptimizationBarrier_37_io_x_ae),
    .io_x_sw(pma_checker_OptimizationBarrier_37_io_x_sw),
    .io_x_sx(pma_checker_OptimizationBarrier_37_io_x_sx),
    .io_x_sr(pma_checker_OptimizationBarrier_37_io_x_sr),
    .io_x_pw(pma_checker_OptimizationBarrier_37_io_x_pw),
    .io_x_px(pma_checker_OptimizationBarrier_37_io_x_px),
    .io_x_pr(pma_checker_OptimizationBarrier_37_io_x_pr),
    .io_x_ppp(pma_checker_OptimizationBarrier_37_io_x_ppp),
    .io_x_pal(pma_checker_OptimizationBarrier_37_io_x_pal),
    .io_x_paa(pma_checker_OptimizationBarrier_37_io_x_paa),
    .io_x_eff(pma_checker_OptimizationBarrier_37_io_x_eff),
    .io_x_c(pma_checker_OptimizationBarrier_37_io_x_c),
    .io_y_ppn(pma_checker_OptimizationBarrier_37_io_y_ppn),
    .io_y_u(pma_checker_OptimizationBarrier_37_io_y_u),
    .io_y_ae(pma_checker_OptimizationBarrier_37_io_y_ae),
    .io_y_sw(pma_checker_OptimizationBarrier_37_io_y_sw),
    .io_y_sx(pma_checker_OptimizationBarrier_37_io_y_sx),
    .io_y_sr(pma_checker_OptimizationBarrier_37_io_y_sr),
    .io_y_pw(pma_checker_OptimizationBarrier_37_io_y_pw),
    .io_y_px(pma_checker_OptimizationBarrier_37_io_y_px),
    .io_y_pr(pma_checker_OptimizationBarrier_37_io_y_pr),
    .io_y_ppp(pma_checker_OptimizationBarrier_37_io_y_ppp),
    .io_y_pal(pma_checker_OptimizationBarrier_37_io_y_pal),
    .io_y_paa(pma_checker_OptimizationBarrier_37_io_y_paa),
    .io_y_eff(pma_checker_OptimizationBarrier_37_io_y_eff),
    .io_y_c(pma_checker_OptimizationBarrier_37_io_y_c)
  );
  OptimizationBarrier pma_checker_OptimizationBarrier_38 ( // @[package.scala 231:25:freechips.rocketchip.system.DefaultRV32Config.fir@179672.4]
    .io_x_ppn(pma_checker_OptimizationBarrier_38_io_x_ppn),
    .io_x_u(pma_checker_OptimizationBarrier_38_io_x_u),
    .io_x_ae(pma_checker_OptimizationBarrier_38_io_x_ae),
    .io_x_sw(pma_checker_OptimizationBarrier_38_io_x_sw),
    .io_x_sx(pma_checker_OptimizationBarrier_38_io_x_sx),
    .io_x_sr(pma_checker_OptimizationBarrier_38_io_x_sr),
    .io_x_pw(pma_checker_OptimizationBarrier_38_io_x_pw),
    .io_x_px(pma_checker_OptimizationBarrier_38_io_x_px),
    .io_x_pr(pma_checker_OptimizationBarrier_38_io_x_pr),
    .io_x_ppp(pma_checker_OptimizationBarrier_38_io_x_ppp),
    .io_x_pal(pma_checker_OptimizationBarrier_38_io_x_pal),
    .io_x_paa(pma_checker_OptimizationBarrier_38_io_x_paa),
    .io_x_eff(pma_checker_OptimizationBarrier_38_io_x_eff),
    .io_x_c(pma_checker_OptimizationBarrier_38_io_x_c),
    .io_y_ppn(pma_checker_OptimizationBarrier_38_io_y_ppn),
    .io_y_u(pma_checker_OptimizationBarrier_38_io_y_u),
    .io_y_ae(pma_checker_OptimizationBarrier_38_io_y_ae),
    .io_y_sw(pma_checker_OptimizationBarrier_38_io_y_sw),
    .io_y_sx(pma_checker_OptimizationBarrier_38_io_y_sx),
    .io_y_sr(pma_checker_OptimizationBarrier_38_io_y_sr),
    .io_y_pw(pma_checker_OptimizationBarrier_38_io_y_pw),
    .io_y_px(pma_checker_OptimizationBarrier_38_io_y_px),
    .io_y_pr(pma_checker_OptimizationBarrier_38_io_y_pr),
    .io_y_ppp(pma_checker_OptimizationBarrier_38_io_y_ppp),
    .io_y_pal(pma_checker_OptimizationBarrier_38_io_y_pal),
    .io_y_paa(pma_checker_OptimizationBarrier_38_io_y_paa),
    .io_y_eff(pma_checker_OptimizationBarrier_38_io_y_eff),
    .io_y_c(pma_checker_OptimizationBarrier_38_io_y_c)
  );
  MaxPeriodFibonacciLFSR MaxPeriodFibonacciLFSR ( // @[PRNG.scala 82:22:freechips.rocketchip.system.DefaultRV32Config.fir@192119.4]
    .clock(MaxPeriodFibonacciLFSR_clock),
    .reset(MaxPeriodFibonacciLFSR_reset),
    .io_increment(MaxPeriodFibonacciLFSR_io_increment),
    .io_out_0(MaxPeriodFibonacciLFSR_io_out_0),
    .io_out_1(MaxPeriodFibonacciLFSR_io_out_1),
    .io_out_2(MaxPeriodFibonacciLFSR_io_out_2),
    .io_out_3(MaxPeriodFibonacciLFSR_io_out_3),
    .io_out_4(MaxPeriodFibonacciLFSR_io_out_4),
    .io_out_5(MaxPeriodFibonacciLFSR_io_out_5),
    .io_out_6(MaxPeriodFibonacciLFSR_io_out_6),
    .io_out_7(MaxPeriodFibonacciLFSR_io_out_7),
    .io_out_8(MaxPeriodFibonacciLFSR_io_out_8),
    .io_out_9(MaxPeriodFibonacciLFSR_io_out_9),
    .io_out_10(MaxPeriodFibonacciLFSR_io_out_10),
    .io_out_11(MaxPeriodFibonacciLFSR_io_out_11),
    .io_out_12(MaxPeriodFibonacciLFSR_io_out_12),
    .io_out_13(MaxPeriodFibonacciLFSR_io_out_13),
    .io_out_14(MaxPeriodFibonacciLFSR_io_out_14),
    .io_out_15(MaxPeriodFibonacciLFSR_io_out_15)
  );
  tag_array tag_array ( // @[DescribedSRAM.scala 23:26:freechips.rocketchip.system.DefaultRV32Config.fir@192159.4]
    .RW0_addr(tag_array_RW0_addr),
    .RW0_en(tag_array_RW0_en),
    .RW0_clk(tag_array_RW0_clk),
    .RW0_wmode(tag_array_RW0_wmode),
    .RW0_wdata_0(tag_array_RW0_wdata_0),
    .RW0_wdata_1(tag_array_RW0_wdata_1),
    .RW0_wdata_2(tag_array_RW0_wdata_2),
    .RW0_wdata_3(tag_array_RW0_wdata_3),
    .RW0_rdata_0(tag_array_RW0_rdata_0),
    .RW0_rdata_1(tag_array_RW0_rdata_1),
    .RW0_rdata_2(tag_array_RW0_rdata_2),
    .RW0_rdata_3(tag_array_RW0_rdata_3),
    .RW0_wmask_0(tag_array_RW0_wmask_0),
    .RW0_wmask_1(tag_array_RW0_wmask_1),
    .RW0_wmask_2(tag_array_RW0_wmask_2),
    .RW0_wmask_3(tag_array_RW0_wmask_3)
  );
  DCacheDataArray data ( // @[DCache.scala 130:20:freechips.rocketchip.system.DefaultRV32Config.fir@192160.4]
    .clock(data_clock),
    .io_req_valid(data_io_req_valid),
    .io_req_bits_addr(data_io_req_bits_addr),
    .io_req_bits_write(data_io_req_bits_write),
    .io_req_bits_wdata(data_io_req_bits_wdata),
    .io_req_bits_eccMask(data_io_req_bits_eccMask),
    .io_req_bits_way_en(data_io_req_bits_way_en),
    .io_resp_0(data_io_resp_0),
    .io_resp_1(data_io_resp_1),
    .io_resp_2(data_io_resp_2),
    .io_resp_3(data_io_resp_3)
  );
  AMOALU amoalu ( // @[DCache.scala 881:26:freechips.rocketchip.system.DefaultRV32Config.fir@195706.4]
    .io_mask(amoalu_io_mask),
    .io_cmd(amoalu_io_cmd),
    .io_lhs(amoalu_io_lhs),
    .io_rhs(amoalu_io_rhs),
    .io_out(amoalu_io_out)
  );
  assign tlb_priv_s = tlb_io_ptw_status_dprv[0]; // @[TLB.scala 177:20:freechips.rocketchip.system.DefaultRV32Config.fir@176856.4]
  assign tlb_priv_uses_vm = tlb_io_ptw_status_dprv <= 2'h1; // @[TLB.scala 178:27:freechips.rocketchip.system.DefaultRV32Config.fir@176857.4]
  assign tlb__T_2 = tlb_io_ptw_ptbr_mode & tlb_priv_uses_vm; // @[TLB.scala 179:83:freechips.rocketchip.system.DefaultRV32Config.fir@176860.4]
  assign tlb__T_3 = ~tlb_io_req_bits_passthrough; // @[TLB.scala 179:102:freechips.rocketchip.system.DefaultRV32Config.fir@176861.4]
  assign tlb_vm_enabled = tlb__T_2 & tlb__T_3; // @[TLB.scala 179:99:freechips.rocketchip.system.DefaultRV32Config.fir@176862.4]
  assign tlb_vpn = tlb_io_req_bits_vaddr[31:12]; // @[TLB.scala 182:30:freechips.rocketchip.system.DefaultRV32Config.fir@176863.4]
  assign tlb_refill_ppn = tlb_io_ptw_resp_bits_pte_ppn[19:0]; // @[TLB.scala 183:44:freechips.rocketchip.system.DefaultRV32Config.fir@176864.4]
  assign tlb__T_4 = tlb_state == 2'h1; // @[package.scala 15:47:freechips.rocketchip.system.DefaultRV32Config.fir@176866.4]
  assign tlb__T_5 = tlb_state == 2'h3; // @[package.scala 15:47:freechips.rocketchip.system.DefaultRV32Config.fir@176867.4]
  assign tlb_invalidate_refill = tlb__T_4 | tlb__T_5; // @[package.scala 64:59:freechips.rocketchip.system.DefaultRV32Config.fir@176868.4]
  assign tlb__T_22 = tlb_special_entry_data_0[13]; // @[TLB.scala 86:77:freechips.rocketchip.system.DefaultRV32Config.fir@176901.4]
  assign tlb__T_25 = tlb_OptimizationBarrier_io_y_ppn[19:10]; // @[TLB.scala 106:26:freechips.rocketchip.system.DefaultRV32Config.fir@176912.4]
  assign tlb__T_26 = tlb_special_entry_level < 1'h1; // @[TLB.scala 108:28:freechips.rocketchip.system.DefaultRV32Config.fir@176913.4]
  assign tlb__T_28 = tlb__T_26 ? tlb_vpn : 20'h0; // @[TLB.scala 109:28:freechips.rocketchip.system.DefaultRV32Config.fir@176915.4]
  assign tlb__T_29 = tlb__T_28 | tlb_OptimizationBarrier_io_y_ppn; // @[TLB.scala 109:47:freechips.rocketchip.system.DefaultRV32Config.fir@176916.4]
  assign tlb__T_30 = tlb__T_29[9:0]; // @[TLB.scala 109:58:freechips.rocketchip.system.DefaultRV32Config.fir@176917.4]
  assign tlb__T_31 = {tlb__T_25,tlb__T_30}; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@176918.4]
  assign tlb__T_32 = tlb_io_req_bits_vaddr[31:12]; // @[TLB.scala 187:123:freechips.rocketchip.system.DefaultRV32Config.fir@176919.4]
  assign tlb__T_33 = tlb_vm_enabled ? tlb__T_31 : tlb__T_32; // @[TLB.scala 187:20:freechips.rocketchip.system.DefaultRV32Config.fir@176920.4]
  assign tlb_mpu_ppn = tlb_io_ptw_resp_valid ? tlb_refill_ppn : tlb__T_33; // @[TLB.scala 186:20:freechips.rocketchip.system.DefaultRV32Config.fir@176921.4]
  assign tlb__T_34 = tlb_io_req_bits_vaddr[11:0]; // @[TLB.scala 188:52:freechips.rocketchip.system.DefaultRV32Config.fir@176922.4]
  assign tlb_mpu_physaddr = {tlb_mpu_ppn,tlb__T_34}; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@176923.4]
  assign tlb__T_35 = tlb_io_ptw_resp_valid | tlb_io_req_bits_passthrough; // @[TLB.scala 189:56:freechips.rocketchip.system.DefaultRV32Config.fir@176924.4]
  assign tlb__T_37 = {tlb_io_ptw_status_debug,tlb_io_ptw_status_dprv}; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@176926.4]
  assign tlb_mpu_priv = tlb__T_35 ? 3'h1 : tlb__T_37; // @[TLB.scala 189:27:freechips.rocketchip.system.DefaultRV32Config.fir@176927.4]
  assign tlb__T_38 = tlb_mpu_physaddr ^ 32'h3000; // @[Parameters.scala 137:31:freechips.rocketchip.system.DefaultRV32Config.fir@176943.4]
  assign tlb__T_39 = {1'b0,$signed(tlb__T_38)}; // @[Parameters.scala 137:49:freechips.rocketchip.system.DefaultRV32Config.fir@176944.4]
  assign tlb__T_41 = $signed(tlb__T_39) & -33'sh1000; // @[Parameters.scala 137:52:freechips.rocketchip.system.DefaultRV32Config.fir@176946.4]
  assign tlb__T_42 = $signed(tlb__T_41) == 33'sh0; // @[Parameters.scala 137:67:freechips.rocketchip.system.DefaultRV32Config.fir@176947.4]
  assign tlb__T_43 = tlb_mpu_physaddr ^ 32'hc000000; // @[Parameters.scala 137:31:freechips.rocketchip.system.DefaultRV32Config.fir@176948.4]
  assign tlb__T_44 = {1'b0,$signed(tlb__T_43)}; // @[Parameters.scala 137:49:freechips.rocketchip.system.DefaultRV32Config.fir@176949.4]
  assign tlb__T_46 = $signed(tlb__T_44) & -33'sh4000000; // @[Parameters.scala 137:52:freechips.rocketchip.system.DefaultRV32Config.fir@176951.4]
  assign tlb__T_47 = $signed(tlb__T_46) == 33'sh0; // @[Parameters.scala 137:67:freechips.rocketchip.system.DefaultRV32Config.fir@176952.4]
  assign tlb__T_48 = tlb_mpu_physaddr ^ 32'h2000000; // @[Parameters.scala 137:31:freechips.rocketchip.system.DefaultRV32Config.fir@176953.4]
  assign tlb__T_49 = {1'b0,$signed(tlb__T_48)}; // @[Parameters.scala 137:49:freechips.rocketchip.system.DefaultRV32Config.fir@176954.4]
  assign tlb__T_51 = $signed(tlb__T_49) & -33'sh10000; // @[Parameters.scala 137:52:freechips.rocketchip.system.DefaultRV32Config.fir@176956.4]
  assign tlb__T_52 = $signed(tlb__T_51) == 33'sh0; // @[Parameters.scala 137:67:freechips.rocketchip.system.DefaultRV32Config.fir@176957.4]
  assign tlb__T_54 = {1'b0,$signed(tlb_mpu_physaddr)}; // @[Parameters.scala 137:49:freechips.rocketchip.system.DefaultRV32Config.fir@176959.4]
  assign tlb__T_56 = $signed(tlb__T_54) & -33'sh1000; // @[Parameters.scala 137:52:freechips.rocketchip.system.DefaultRV32Config.fir@176961.4]
  assign tlb__T_57 = $signed(tlb__T_56) == 33'sh0; // @[Parameters.scala 137:67:freechips.rocketchip.system.DefaultRV32Config.fir@176962.4]
  assign tlb__T_58 = tlb_mpu_physaddr ^ 32'h10000; // @[Parameters.scala 137:31:freechips.rocketchip.system.DefaultRV32Config.fir@176963.4]
  assign tlb__T_59 = {1'b0,$signed(tlb__T_58)}; // @[Parameters.scala 137:49:freechips.rocketchip.system.DefaultRV32Config.fir@176964.4]
  assign tlb__T_61 = $signed(tlb__T_59) & -33'sh10000; // @[Parameters.scala 137:52:freechips.rocketchip.system.DefaultRV32Config.fir@176966.4]
  assign tlb__T_62 = $signed(tlb__T_61) == 33'sh0; // @[Parameters.scala 137:67:freechips.rocketchip.system.DefaultRV32Config.fir@176967.4]
  assign tlb__T_63 = tlb_mpu_physaddr ^ 32'h80000000; // @[Parameters.scala 137:31:freechips.rocketchip.system.DefaultRV32Config.fir@176968.4]
  assign tlb__T_64 = {1'b0,$signed(tlb__T_63)}; // @[Parameters.scala 137:49:freechips.rocketchip.system.DefaultRV32Config.fir@176969.4]
  assign tlb__T_66 = $signed(tlb__T_64) & -33'sh10000000; // @[Parameters.scala 137:52:freechips.rocketchip.system.DefaultRV32Config.fir@176971.4]
  assign tlb__T_67 = $signed(tlb__T_66) == 33'sh0; // @[Parameters.scala 137:67:freechips.rocketchip.system.DefaultRV32Config.fir@176972.4]
  assign tlb__T_68 = tlb_mpu_physaddr ^ 32'h60000000; // @[Parameters.scala 137:31:freechips.rocketchip.system.DefaultRV32Config.fir@176973.4]
  assign tlb__T_69 = {1'b0,$signed(tlb__T_68)}; // @[Parameters.scala 137:49:freechips.rocketchip.system.DefaultRV32Config.fir@176974.4]
  assign tlb__T_71 = $signed(tlb__T_69) & -33'sh20000000; // @[Parameters.scala 137:52:freechips.rocketchip.system.DefaultRV32Config.fir@176976.4]
  assign tlb__T_72 = $signed(tlb__T_71) == 33'sh0; // @[Parameters.scala 137:67:freechips.rocketchip.system.DefaultRV32Config.fir@176977.4]
  assign tlb__T_74 = tlb__T_42 | tlb__T_47; // @[TLB.scala 195:67:freechips.rocketchip.system.DefaultRV32Config.fir@176987.4]
  assign tlb__T_75 = tlb__T_74 | tlb__T_52; // @[TLB.scala 195:67:freechips.rocketchip.system.DefaultRV32Config.fir@176988.4]
  assign tlb__T_76 = tlb__T_75 | tlb__T_57; // @[TLB.scala 195:67:freechips.rocketchip.system.DefaultRV32Config.fir@176989.4]
  assign tlb__T_77 = tlb__T_76 | tlb__T_62; // @[TLB.scala 195:67:freechips.rocketchip.system.DefaultRV32Config.fir@176990.4]
  assign tlb__T_78 = tlb__T_77 | tlb__T_67; // @[TLB.scala 195:67:freechips.rocketchip.system.DefaultRV32Config.fir@176991.4]
  assign tlb_legal_address = tlb__T_78 | tlb__T_72; // @[TLB.scala 195:67:freechips.rocketchip.system.DefaultRV32Config.fir@176992.4]
  assign tlb__T_87 = $signed(tlb__T_64) & 33'sh80000000; // @[Parameters.scala 137:52:freechips.rocketchip.system.DefaultRV32Config.fir@177001.4]
  assign tlb__T_88 = $signed(tlb__T_87) == 33'sh0; // @[Parameters.scala 137:67:freechips.rocketchip.system.DefaultRV32Config.fir@177002.4]
  assign tlb__T_93 = tlb_legal_address & tlb__T_88; // @[TLB.scala 197:19:freechips.rocketchip.system.DefaultRV32Config.fir@177008.4]
  assign tlb__T_148 = tlb_mpu_physaddr ^ 32'h8000000; // @[Parameters.scala 137:31:freechips.rocketchip.system.DefaultRV32Config.fir@177065.4]
  assign tlb__T_149 = {1'b0,$signed(tlb__T_148)}; // @[Parameters.scala 137:49:freechips.rocketchip.system.DefaultRV32Config.fir@177066.4]
  assign tlb__T_151 = $signed(tlb__T_149) & 33'shc8000000; // @[Parameters.scala 137:52:freechips.rocketchip.system.DefaultRV32Config.fir@177068.4]
  assign tlb__T_152 = $signed(tlb__T_151) == 33'sh0; // @[Parameters.scala 137:67:freechips.rocketchip.system.DefaultRV32Config.fir@177069.4]
  assign tlb__T_165 = $signed(tlb__T_54) & 33'shc8010000; // @[Parameters.scala 137:52:freechips.rocketchip.system.DefaultRV32Config.fir@177082.4]
  assign tlb__T_166 = $signed(tlb__T_165) == 33'sh0; // @[Parameters.scala 137:67:freechips.rocketchip.system.DefaultRV32Config.fir@177083.4]
  assign tlb__T_173 = tlb__T_166 | tlb__T_152; // @[TLBPermissions.scala 82:66:freechips.rocketchip.system.DefaultRV32Config.fir@177090.4]
  assign tlb__T_186 = tlb_mpu_priv <= 3'h3; // @[TLB.scala 200:39:freechips.rocketchip.system.DefaultRV32Config.fir@177103.4]
  assign tlb_deny_access_to_debug = tlb__T_186 & tlb__T_57; // @[TLB.scala 200:48:freechips.rocketchip.system.DefaultRV32Config.fir@177109.4]
  assign tlb__T_198 = ~tlb_deny_access_to_debug; // @[TLB.scala 201:44:freechips.rocketchip.system.DefaultRV32Config.fir@177116.4]
  assign tlb__T_199 = tlb_legal_address & tlb__T_198; // @[TLB.scala 201:41:freechips.rocketchip.system.DefaultRV32Config.fir@177117.4]
  assign tlb_prot_r = tlb__T_199 & tlb_pmp_io_r; // @[TLB.scala 201:66:freechips.rocketchip.system.DefaultRV32Config.fir@177118.4]
  assign tlb__T_210 = tlb_mpu_physaddr ^ 32'h40000000; // @[Parameters.scala 137:31:freechips.rocketchip.system.DefaultRV32Config.fir@177129.4]
  assign tlb__T_211 = {1'b0,$signed(tlb__T_210)}; // @[Parameters.scala 137:49:freechips.rocketchip.system.DefaultRV32Config.fir@177130.4]
  assign tlb__T_213 = $signed(tlb__T_211) & 33'shc0000000; // @[Parameters.scala 137:52:freechips.rocketchip.system.DefaultRV32Config.fir@177132.4]
  assign tlb__T_214 = $signed(tlb__T_213) == 33'sh0; // @[Parameters.scala 137:67:freechips.rocketchip.system.DefaultRV32Config.fir@177133.4]
  assign tlb__T_218 = $signed(tlb__T_64) & 33'shc0000000; // @[Parameters.scala 137:52:freechips.rocketchip.system.DefaultRV32Config.fir@177137.4]
  assign tlb__T_219 = $signed(tlb__T_218) == 33'sh0; // @[Parameters.scala 137:67:freechips.rocketchip.system.DefaultRV32Config.fir@177138.4]
  assign tlb__T_221 = tlb__T_173 | tlb__T_214; // @[Parameters.scala 528:89:freechips.rocketchip.system.DefaultRV32Config.fir@177140.4]
  assign tlb__T_222 = tlb__T_221 | tlb__T_219; // @[Parameters.scala 528:89:freechips.rocketchip.system.DefaultRV32Config.fir@177141.4]
  assign tlb__T_232 = tlb_legal_address & tlb__T_222; // @[TLB.scala 197:19:freechips.rocketchip.system.DefaultRV32Config.fir@177152.4]
  assign tlb__T_234 = tlb__T_232 & tlb__T_198; // @[TLB.scala 202:45:freechips.rocketchip.system.DefaultRV32Config.fir@177154.4]
  assign tlb_prot_w = tlb__T_234 & tlb_pmp_io_w; // @[TLB.scala 202:70:freechips.rocketchip.system.DefaultRV32Config.fir@177155.4]
  assign tlb_prot_al = tlb_legal_address & tlb__T_173; // @[TLB.scala 197:19:freechips.rocketchip.system.DefaultRV32Config.fir@177223.4]
  assign tlb__T_334 = $signed(tlb__T_54) & 33'shca000000; // @[Parameters.scala 137:52:freechips.rocketchip.system.DefaultRV32Config.fir@177261.4]
  assign tlb__T_335 = $signed(tlb__T_334) == 33'sh0; // @[Parameters.scala 137:67:freechips.rocketchip.system.DefaultRV32Config.fir@177262.4]
  assign tlb__T_346 = tlb__T_335 | tlb__T_214; // @[Parameters.scala 528:89:freechips.rocketchip.system.DefaultRV32Config.fir@177273.4]
  assign tlb__T_347 = tlb__T_346 | tlb__T_219; // @[Parameters.scala 528:89:freechips.rocketchip.system.DefaultRV32Config.fir@177274.4]
  assign tlb__T_363 = tlb_legal_address & tlb__T_347; // @[TLB.scala 197:19:freechips.rocketchip.system.DefaultRV32Config.fir@177291.4]
  assign tlb__T_365 = tlb__T_363 & tlb__T_198; // @[TLB.scala 206:40:freechips.rocketchip.system.DefaultRV32Config.fir@177293.4]
  assign tlb_prot_x = tlb__T_365 & tlb_pmp_io_x; // @[TLB.scala 206:65:freechips.rocketchip.system.DefaultRV32Config.fir@177294.4]
  assign tlb__T_386 = $signed(tlb__T_54) & 33'shca012000; // @[Parameters.scala 137:52:freechips.rocketchip.system.DefaultRV32Config.fir@177315.4]
  assign tlb__T_387 = $signed(tlb__T_386) == 33'sh0; // @[Parameters.scala 137:67:freechips.rocketchip.system.DefaultRV32Config.fir@177316.4]
  assign tlb__T_391 = $signed(tlb__T_49) & 33'shca010000; // @[Parameters.scala 137:52:freechips.rocketchip.system.DefaultRV32Config.fir@177320.4]
  assign tlb__T_392 = $signed(tlb__T_391) == 33'sh0; // @[Parameters.scala 137:67:freechips.rocketchip.system.DefaultRV32Config.fir@177321.4]
  assign tlb__T_403 = tlb__T_387 | tlb__T_392; // @[Parameters.scala 528:89:freechips.rocketchip.system.DefaultRV32Config.fir@177332.4]
  assign tlb__T_404 = tlb__T_403 | tlb__T_152; // @[Parameters.scala 528:89:freechips.rocketchip.system.DefaultRV32Config.fir@177333.4]
  assign tlb__T_405 = tlb__T_404 | tlb__T_214; // @[Parameters.scala 528:89:freechips.rocketchip.system.DefaultRV32Config.fir@177334.4]
  assign tlb_prot_eff = tlb_legal_address & tlb__T_405; // @[TLB.scala 197:19:freechips.rocketchip.system.DefaultRV32Config.fir@177340.4]
  assign tlb__T_410 = tlb_sectored_entries_0_valid_0 | tlb_sectored_entries_0_valid_1; // @[package.scala 64:59:freechips.rocketchip.system.DefaultRV32Config.fir@177341.4]
  assign tlb__T_411 = tlb__T_410 | tlb_sectored_entries_0_valid_2; // @[package.scala 64:59:freechips.rocketchip.system.DefaultRV32Config.fir@177342.4]
  assign tlb__T_412 = tlb__T_411 | tlb_sectored_entries_0_valid_3; // @[package.scala 64:59:freechips.rocketchip.system.DefaultRV32Config.fir@177343.4]
  assign tlb__T_413 = tlb_sectored_entries_0_tag ^ tlb_vpn; // @[TLB.scala 88:41:freechips.rocketchip.system.DefaultRV32Config.fir@177344.4]
  assign tlb__T_414 = tlb__T_413[19:2]; // @[TLB.scala 88:48:freechips.rocketchip.system.DefaultRV32Config.fir@177345.4]
  assign tlb__T_415 = tlb__T_414 == 18'h0; // @[TLB.scala 88:66:freechips.rocketchip.system.DefaultRV32Config.fir@177346.4]
  assign tlb_sector_hits_0 = tlb__T_412 & tlb__T_415; // @[TLB.scala 87:40:freechips.rocketchip.system.DefaultRV32Config.fir@177347.4]
  assign tlb__T_416 = tlb_sectored_entries_1_valid_0 | tlb_sectored_entries_1_valid_1; // @[package.scala 64:59:freechips.rocketchip.system.DefaultRV32Config.fir@177348.4]
  assign tlb__T_417 = tlb__T_416 | tlb_sectored_entries_1_valid_2; // @[package.scala 64:59:freechips.rocketchip.system.DefaultRV32Config.fir@177349.4]
  assign tlb__T_418 = tlb__T_417 | tlb_sectored_entries_1_valid_3; // @[package.scala 64:59:freechips.rocketchip.system.DefaultRV32Config.fir@177350.4]
  assign tlb__T_419 = tlb_sectored_entries_1_tag ^ tlb_vpn; // @[TLB.scala 88:41:freechips.rocketchip.system.DefaultRV32Config.fir@177351.4]
  assign tlb__T_420 = tlb__T_419[19:2]; // @[TLB.scala 88:48:freechips.rocketchip.system.DefaultRV32Config.fir@177352.4]
  assign tlb__T_421 = tlb__T_420 == 18'h0; // @[TLB.scala 88:66:freechips.rocketchip.system.DefaultRV32Config.fir@177353.4]
  assign tlb_sector_hits_1 = tlb__T_418 & tlb__T_421; // @[TLB.scala 87:40:freechips.rocketchip.system.DefaultRV32Config.fir@177354.4]
  assign tlb__T_422 = tlb_sectored_entries_2_valid_0 | tlb_sectored_entries_2_valid_1; // @[package.scala 64:59:freechips.rocketchip.system.DefaultRV32Config.fir@177355.4]
  assign tlb__T_423 = tlb__T_422 | tlb_sectored_entries_2_valid_2; // @[package.scala 64:59:freechips.rocketchip.system.DefaultRV32Config.fir@177356.4]
  assign tlb__T_424 = tlb__T_423 | tlb_sectored_entries_2_valid_3; // @[package.scala 64:59:freechips.rocketchip.system.DefaultRV32Config.fir@177357.4]
  assign tlb__T_425 = tlb_sectored_entries_2_tag ^ tlb_vpn; // @[TLB.scala 88:41:freechips.rocketchip.system.DefaultRV32Config.fir@177358.4]
  assign tlb__T_426 = tlb__T_425[19:2]; // @[TLB.scala 88:48:freechips.rocketchip.system.DefaultRV32Config.fir@177359.4]
  assign tlb__T_427 = tlb__T_426 == 18'h0; // @[TLB.scala 88:66:freechips.rocketchip.system.DefaultRV32Config.fir@177360.4]
  assign tlb_sector_hits_2 = tlb__T_424 & tlb__T_427; // @[TLB.scala 87:40:freechips.rocketchip.system.DefaultRV32Config.fir@177361.4]
  assign tlb__T_428 = tlb_sectored_entries_3_valid_0 | tlb_sectored_entries_3_valid_1; // @[package.scala 64:59:freechips.rocketchip.system.DefaultRV32Config.fir@177362.4]
  assign tlb__T_429 = tlb__T_428 | tlb_sectored_entries_3_valid_2; // @[package.scala 64:59:freechips.rocketchip.system.DefaultRV32Config.fir@177363.4]
  assign tlb__T_430 = tlb__T_429 | tlb_sectored_entries_3_valid_3; // @[package.scala 64:59:freechips.rocketchip.system.DefaultRV32Config.fir@177364.4]
  assign tlb__T_431 = tlb_sectored_entries_3_tag ^ tlb_vpn; // @[TLB.scala 88:41:freechips.rocketchip.system.DefaultRV32Config.fir@177365.4]
  assign tlb__T_432 = tlb__T_431[19:2]; // @[TLB.scala 88:48:freechips.rocketchip.system.DefaultRV32Config.fir@177366.4]
  assign tlb__T_433 = tlb__T_432 == 18'h0; // @[TLB.scala 88:66:freechips.rocketchip.system.DefaultRV32Config.fir@177367.4]
  assign tlb_sector_hits_3 = tlb__T_430 & tlb__T_433; // @[TLB.scala 87:40:freechips.rocketchip.system.DefaultRV32Config.fir@177368.4]
  assign tlb__T_434 = tlb_sectored_entries_4_valid_0 | tlb_sectored_entries_4_valid_1; // @[package.scala 64:59:freechips.rocketchip.system.DefaultRV32Config.fir@177369.4]
  assign tlb__T_435 = tlb__T_434 | tlb_sectored_entries_4_valid_2; // @[package.scala 64:59:freechips.rocketchip.system.DefaultRV32Config.fir@177370.4]
  assign tlb__T_436 = tlb__T_435 | tlb_sectored_entries_4_valid_3; // @[package.scala 64:59:freechips.rocketchip.system.DefaultRV32Config.fir@177371.4]
  assign tlb__T_437 = tlb_sectored_entries_4_tag ^ tlb_vpn; // @[TLB.scala 88:41:freechips.rocketchip.system.DefaultRV32Config.fir@177372.4]
  assign tlb__T_438 = tlb__T_437[19:2]; // @[TLB.scala 88:48:freechips.rocketchip.system.DefaultRV32Config.fir@177373.4]
  assign tlb__T_439 = tlb__T_438 == 18'h0; // @[TLB.scala 88:66:freechips.rocketchip.system.DefaultRV32Config.fir@177374.4]
  assign tlb_sector_hits_4 = tlb__T_436 & tlb__T_439; // @[TLB.scala 87:40:freechips.rocketchip.system.DefaultRV32Config.fir@177375.4]
  assign tlb__T_440 = tlb_sectored_entries_5_valid_0 | tlb_sectored_entries_5_valid_1; // @[package.scala 64:59:freechips.rocketchip.system.DefaultRV32Config.fir@177376.4]
  assign tlb__T_441 = tlb__T_440 | tlb_sectored_entries_5_valid_2; // @[package.scala 64:59:freechips.rocketchip.system.DefaultRV32Config.fir@177377.4]
  assign tlb__T_442 = tlb__T_441 | tlb_sectored_entries_5_valid_3; // @[package.scala 64:59:freechips.rocketchip.system.DefaultRV32Config.fir@177378.4]
  assign tlb__T_443 = tlb_sectored_entries_5_tag ^ tlb_vpn; // @[TLB.scala 88:41:freechips.rocketchip.system.DefaultRV32Config.fir@177379.4]
  assign tlb__T_444 = tlb__T_443[19:2]; // @[TLB.scala 88:48:freechips.rocketchip.system.DefaultRV32Config.fir@177380.4]
  assign tlb__T_445 = tlb__T_444 == 18'h0; // @[TLB.scala 88:66:freechips.rocketchip.system.DefaultRV32Config.fir@177381.4]
  assign tlb_sector_hits_5 = tlb__T_442 & tlb__T_445; // @[TLB.scala 87:40:freechips.rocketchip.system.DefaultRV32Config.fir@177382.4]
  assign tlb__T_446 = tlb_sectored_entries_6_valid_0 | tlb_sectored_entries_6_valid_1; // @[package.scala 64:59:freechips.rocketchip.system.DefaultRV32Config.fir@177383.4]
  assign tlb__T_447 = tlb__T_446 | tlb_sectored_entries_6_valid_2; // @[package.scala 64:59:freechips.rocketchip.system.DefaultRV32Config.fir@177384.4]
  assign tlb__T_448 = tlb__T_447 | tlb_sectored_entries_6_valid_3; // @[package.scala 64:59:freechips.rocketchip.system.DefaultRV32Config.fir@177385.4]
  assign tlb__T_449 = tlb_sectored_entries_6_tag ^ tlb_vpn; // @[TLB.scala 88:41:freechips.rocketchip.system.DefaultRV32Config.fir@177386.4]
  assign tlb__T_450 = tlb__T_449[19:2]; // @[TLB.scala 88:48:freechips.rocketchip.system.DefaultRV32Config.fir@177387.4]
  assign tlb__T_451 = tlb__T_450 == 18'h0; // @[TLB.scala 88:66:freechips.rocketchip.system.DefaultRV32Config.fir@177388.4]
  assign tlb_sector_hits_6 = tlb__T_448 & tlb__T_451; // @[TLB.scala 87:40:freechips.rocketchip.system.DefaultRV32Config.fir@177389.4]
  assign tlb__T_452 = tlb_sectored_entries_7_valid_0 | tlb_sectored_entries_7_valid_1; // @[package.scala 64:59:freechips.rocketchip.system.DefaultRV32Config.fir@177390.4]
  assign tlb__T_453 = tlb__T_452 | tlb_sectored_entries_7_valid_2; // @[package.scala 64:59:freechips.rocketchip.system.DefaultRV32Config.fir@177391.4]
  assign tlb__T_454 = tlb__T_453 | tlb_sectored_entries_7_valid_3; // @[package.scala 64:59:freechips.rocketchip.system.DefaultRV32Config.fir@177392.4]
  assign tlb__T_455 = tlb_sectored_entries_7_tag ^ tlb_vpn; // @[TLB.scala 88:41:freechips.rocketchip.system.DefaultRV32Config.fir@177393.4]
  assign tlb__T_456 = tlb__T_455[19:2]; // @[TLB.scala 88:48:freechips.rocketchip.system.DefaultRV32Config.fir@177394.4]
  assign tlb__T_457 = tlb__T_456 == 18'h0; // @[TLB.scala 88:66:freechips.rocketchip.system.DefaultRV32Config.fir@177395.4]
  assign tlb_sector_hits_7 = tlb__T_454 & tlb__T_457; // @[TLB.scala 87:40:freechips.rocketchip.system.DefaultRV32Config.fir@177396.4]
  assign tlb__T_460 = tlb_superpage_entries_0_tag[19:10]; // @[TLB.scala 95:46:freechips.rocketchip.system.DefaultRV32Config.fir@177399.4]
  assign tlb__T_461 = tlb_vpn[19:10]; // @[TLB.scala 95:84:freechips.rocketchip.system.DefaultRV32Config.fir@177400.4]
  assign tlb__T_462 = tlb__T_460 == tlb__T_461; // @[TLB.scala 95:77:freechips.rocketchip.system.DefaultRV32Config.fir@177401.4]
  assign tlb__T_464 = tlb_superpage_entries_0_valid_0 & tlb__T_462; // @[TLB.scala 95:29:freechips.rocketchip.system.DefaultRV32Config.fir@177403.4]
  assign tlb__T_468 = tlb_vpn[9:0]; // @[TLB.scala 95:84:freechips.rocketchip.system.DefaultRV32Config.fir@177407.4]
  assign tlb__T_473 = tlb_superpage_entries_1_tag[19:10]; // @[TLB.scala 95:46:freechips.rocketchip.system.DefaultRV32Config.fir@177413.4]
  assign tlb__T_475 = tlb__T_473 == tlb__T_461; // @[TLB.scala 95:77:freechips.rocketchip.system.DefaultRV32Config.fir@177415.4]
  assign tlb__T_477 = tlb_superpage_entries_1_valid_0 & tlb__T_475; // @[TLB.scala 95:29:freechips.rocketchip.system.DefaultRV32Config.fir@177417.4]
  assign tlb__T_486 = tlb_superpage_entries_2_tag[19:10]; // @[TLB.scala 95:46:freechips.rocketchip.system.DefaultRV32Config.fir@177427.4]
  assign tlb__T_488 = tlb__T_486 == tlb__T_461; // @[TLB.scala 95:77:freechips.rocketchip.system.DefaultRV32Config.fir@177429.4]
  assign tlb__T_490 = tlb_superpage_entries_2_valid_0 & tlb__T_488; // @[TLB.scala 95:29:freechips.rocketchip.system.DefaultRV32Config.fir@177431.4]
  assign tlb__T_499 = tlb_superpage_entries_3_tag[19:10]; // @[TLB.scala 95:46:freechips.rocketchip.system.DefaultRV32Config.fir@177441.4]
  assign tlb__T_501 = tlb__T_499 == tlb__T_461; // @[TLB.scala 95:77:freechips.rocketchip.system.DefaultRV32Config.fir@177443.4]
  assign tlb__T_503 = tlb_superpage_entries_3_valid_0 & tlb__T_501; // @[TLB.scala 95:29:freechips.rocketchip.system.DefaultRV32Config.fir@177445.4]
  assign tlb__T_510 = tlb_vpn[1:0]; // @[package.scala 138:13:freechips.rocketchip.system.DefaultRV32Config.fir@177453.4]
  assign tlb__GEN_1 = 2'h1 == tlb__T_510 ? tlb_sectored_entries_0_valid_1 : tlb_sectored_entries_0_valid_0; // @[TLB.scala 100:18:freechips.rocketchip.system.DefaultRV32Config.fir@177457.4]
  assign tlb__GEN_2 = 2'h2 == tlb__T_510 ? tlb_sectored_entries_0_valid_2 : tlb__GEN_1; // @[TLB.scala 100:18:freechips.rocketchip.system.DefaultRV32Config.fir@177457.4]
  assign tlb__GEN_3 = 2'h3 == tlb__T_510 ? tlb_sectored_entries_0_valid_3 : tlb__GEN_2; // @[TLB.scala 100:18:freechips.rocketchip.system.DefaultRV32Config.fir@177457.4]
  assign tlb__T_514 = tlb__GEN_3 & tlb__T_415; // @[TLB.scala 100:18:freechips.rocketchip.system.DefaultRV32Config.fir@177457.4]
  assign tlb_hitsVec_0 = tlb_vm_enabled & tlb__T_514; // @[TLB.scala 211:44:freechips.rocketchip.system.DefaultRV32Config.fir@177458.4]
  assign tlb__GEN_5 = 2'h1 == tlb__T_510 ? tlb_sectored_entries_1_valid_1 : tlb_sectored_entries_1_valid_0; // @[TLB.scala 100:18:freechips.rocketchip.system.DefaultRV32Config.fir@177463.4]
  assign tlb__GEN_6 = 2'h2 == tlb__T_510 ? tlb_sectored_entries_1_valid_2 : tlb__GEN_5; // @[TLB.scala 100:18:freechips.rocketchip.system.DefaultRV32Config.fir@177463.4]
  assign tlb__GEN_7 = 2'h3 == tlb__T_510 ? tlb_sectored_entries_1_valid_3 : tlb__GEN_6; // @[TLB.scala 100:18:freechips.rocketchip.system.DefaultRV32Config.fir@177463.4]
  assign tlb__T_519 = tlb__GEN_7 & tlb__T_421; // @[TLB.scala 100:18:freechips.rocketchip.system.DefaultRV32Config.fir@177463.4]
  assign tlb_hitsVec_1 = tlb_vm_enabled & tlb__T_519; // @[TLB.scala 211:44:freechips.rocketchip.system.DefaultRV32Config.fir@177464.4]
  assign tlb__GEN_9 = 2'h1 == tlb__T_510 ? tlb_sectored_entries_2_valid_1 : tlb_sectored_entries_2_valid_0; // @[TLB.scala 100:18:freechips.rocketchip.system.DefaultRV32Config.fir@177469.4]
  assign tlb__GEN_10 = 2'h2 == tlb__T_510 ? tlb_sectored_entries_2_valid_2 : tlb__GEN_9; // @[TLB.scala 100:18:freechips.rocketchip.system.DefaultRV32Config.fir@177469.4]
  assign tlb__GEN_11 = 2'h3 == tlb__T_510 ? tlb_sectored_entries_2_valid_3 : tlb__GEN_10; // @[TLB.scala 100:18:freechips.rocketchip.system.DefaultRV32Config.fir@177469.4]
  assign tlb__T_524 = tlb__GEN_11 & tlb__T_427; // @[TLB.scala 100:18:freechips.rocketchip.system.DefaultRV32Config.fir@177469.4]
  assign tlb_hitsVec_2 = tlb_vm_enabled & tlb__T_524; // @[TLB.scala 211:44:freechips.rocketchip.system.DefaultRV32Config.fir@177470.4]
  assign tlb__GEN_13 = 2'h1 == tlb__T_510 ? tlb_sectored_entries_3_valid_1 : tlb_sectored_entries_3_valid_0; // @[TLB.scala 100:18:freechips.rocketchip.system.DefaultRV32Config.fir@177475.4]
  assign tlb__GEN_14 = 2'h2 == tlb__T_510 ? tlb_sectored_entries_3_valid_2 : tlb__GEN_13; // @[TLB.scala 100:18:freechips.rocketchip.system.DefaultRV32Config.fir@177475.4]
  assign tlb__GEN_15 = 2'h3 == tlb__T_510 ? tlb_sectored_entries_3_valid_3 : tlb__GEN_14; // @[TLB.scala 100:18:freechips.rocketchip.system.DefaultRV32Config.fir@177475.4]
  assign tlb__T_529 = tlb__GEN_15 & tlb__T_433; // @[TLB.scala 100:18:freechips.rocketchip.system.DefaultRV32Config.fir@177475.4]
  assign tlb_hitsVec_3 = tlb_vm_enabled & tlb__T_529; // @[TLB.scala 211:44:freechips.rocketchip.system.DefaultRV32Config.fir@177476.4]
  assign tlb__GEN_17 = 2'h1 == tlb__T_510 ? tlb_sectored_entries_4_valid_1 : tlb_sectored_entries_4_valid_0; // @[TLB.scala 100:18:freechips.rocketchip.system.DefaultRV32Config.fir@177481.4]
  assign tlb__GEN_18 = 2'h2 == tlb__T_510 ? tlb_sectored_entries_4_valid_2 : tlb__GEN_17; // @[TLB.scala 100:18:freechips.rocketchip.system.DefaultRV32Config.fir@177481.4]
  assign tlb__GEN_19 = 2'h3 == tlb__T_510 ? tlb_sectored_entries_4_valid_3 : tlb__GEN_18; // @[TLB.scala 100:18:freechips.rocketchip.system.DefaultRV32Config.fir@177481.4]
  assign tlb__T_534 = tlb__GEN_19 & tlb__T_439; // @[TLB.scala 100:18:freechips.rocketchip.system.DefaultRV32Config.fir@177481.4]
  assign tlb_hitsVec_4 = tlb_vm_enabled & tlb__T_534; // @[TLB.scala 211:44:freechips.rocketchip.system.DefaultRV32Config.fir@177482.4]
  assign tlb__GEN_21 = 2'h1 == tlb__T_510 ? tlb_sectored_entries_5_valid_1 : tlb_sectored_entries_5_valid_0; // @[TLB.scala 100:18:freechips.rocketchip.system.DefaultRV32Config.fir@177487.4]
  assign tlb__GEN_22 = 2'h2 == tlb__T_510 ? tlb_sectored_entries_5_valid_2 : tlb__GEN_21; // @[TLB.scala 100:18:freechips.rocketchip.system.DefaultRV32Config.fir@177487.4]
  assign tlb__GEN_23 = 2'h3 == tlb__T_510 ? tlb_sectored_entries_5_valid_3 : tlb__GEN_22; // @[TLB.scala 100:18:freechips.rocketchip.system.DefaultRV32Config.fir@177487.4]
  assign tlb__T_539 = tlb__GEN_23 & tlb__T_445; // @[TLB.scala 100:18:freechips.rocketchip.system.DefaultRV32Config.fir@177487.4]
  assign tlb_hitsVec_5 = tlb_vm_enabled & tlb__T_539; // @[TLB.scala 211:44:freechips.rocketchip.system.DefaultRV32Config.fir@177488.4]
  assign tlb__GEN_25 = 2'h1 == tlb__T_510 ? tlb_sectored_entries_6_valid_1 : tlb_sectored_entries_6_valid_0; // @[TLB.scala 100:18:freechips.rocketchip.system.DefaultRV32Config.fir@177493.4]
  assign tlb__GEN_26 = 2'h2 == tlb__T_510 ? tlb_sectored_entries_6_valid_2 : tlb__GEN_25; // @[TLB.scala 100:18:freechips.rocketchip.system.DefaultRV32Config.fir@177493.4]
  assign tlb__GEN_27 = 2'h3 == tlb__T_510 ? tlb_sectored_entries_6_valid_3 : tlb__GEN_26; // @[TLB.scala 100:18:freechips.rocketchip.system.DefaultRV32Config.fir@177493.4]
  assign tlb__T_544 = tlb__GEN_27 & tlb__T_451; // @[TLB.scala 100:18:freechips.rocketchip.system.DefaultRV32Config.fir@177493.4]
  assign tlb_hitsVec_6 = tlb_vm_enabled & tlb__T_544; // @[TLB.scala 211:44:freechips.rocketchip.system.DefaultRV32Config.fir@177494.4]
  assign tlb__GEN_29 = 2'h1 == tlb__T_510 ? tlb_sectored_entries_7_valid_1 : tlb_sectored_entries_7_valid_0; // @[TLB.scala 100:18:freechips.rocketchip.system.DefaultRV32Config.fir@177499.4]
  assign tlb__GEN_30 = 2'h2 == tlb__T_510 ? tlb_sectored_entries_7_valid_2 : tlb__GEN_29; // @[TLB.scala 100:18:freechips.rocketchip.system.DefaultRV32Config.fir@177499.4]
  assign tlb__GEN_31 = 2'h3 == tlb__T_510 ? tlb_sectored_entries_7_valid_3 : tlb__GEN_30; // @[TLB.scala 100:18:freechips.rocketchip.system.DefaultRV32Config.fir@177499.4]
  assign tlb__T_549 = tlb__GEN_31 & tlb__T_457; // @[TLB.scala 100:18:freechips.rocketchip.system.DefaultRV32Config.fir@177499.4]
  assign tlb_hitsVec_7 = tlb_vm_enabled & tlb__T_549; // @[TLB.scala 211:44:freechips.rocketchip.system.DefaultRV32Config.fir@177500.4]
  assign tlb_hitsVec_8 = tlb_vm_enabled & tlb__T_464; // @[TLB.scala 211:44:freechips.rocketchip.system.DefaultRV32Config.fir@177515.4]
  assign tlb_hitsVec_9 = tlb_vm_enabled & tlb__T_477; // @[TLB.scala 211:44:freechips.rocketchip.system.DefaultRV32Config.fir@177530.4]
  assign tlb_hitsVec_10 = tlb_vm_enabled & tlb__T_490; // @[TLB.scala 211:44:freechips.rocketchip.system.DefaultRV32Config.fir@177545.4]
  assign tlb_hitsVec_11 = tlb_vm_enabled & tlb__T_503; // @[TLB.scala 211:44:freechips.rocketchip.system.DefaultRV32Config.fir@177560.4]
  assign tlb__T_608 = tlb_special_entry_tag[19:10]; // @[TLB.scala 95:46:freechips.rocketchip.system.DefaultRV32Config.fir@177563.4]
  assign tlb__T_610 = tlb__T_608 == tlb__T_461; // @[TLB.scala 95:77:freechips.rocketchip.system.DefaultRV32Config.fir@177565.4]
  assign tlb__T_612 = tlb_special_entry_valid_0 & tlb__T_610; // @[TLB.scala 95:29:freechips.rocketchip.system.DefaultRV32Config.fir@177567.4]
  assign tlb__T_615 = tlb_special_entry_tag[9:0]; // @[TLB.scala 95:46:freechips.rocketchip.system.DefaultRV32Config.fir@177570.4]
  assign tlb__T_617 = tlb__T_615 == tlb__T_468; // @[TLB.scala 95:77:freechips.rocketchip.system.DefaultRV32Config.fir@177572.4]
  assign tlb__T_618 = tlb__T_26 | tlb__T_617; // @[TLB.scala 95:40:freechips.rocketchip.system.DefaultRV32Config.fir@177573.4]
  assign tlb__T_619 = tlb__T_612 & tlb__T_618; // @[TLB.scala 95:29:freechips.rocketchip.system.DefaultRV32Config.fir@177574.4]
  assign tlb_hitsVec_12 = tlb_vm_enabled & tlb__T_619; // @[TLB.scala 211:44:freechips.rocketchip.system.DefaultRV32Config.fir@177575.4]
  assign tlb__T_624 = {tlb_hitsVec_5,tlb_hitsVec_4,tlb_hitsVec_3,tlb_hitsVec_2,tlb_hitsVec_1,tlb_hitsVec_0}; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@177580.4]
  assign tlb_real_hits = {tlb_hitsVec_12,tlb_hitsVec_11,tlb_hitsVec_10,tlb_hitsVec_9,tlb_hitsVec_8,tlb_hitsVec_7,tlb_hitsVec_6,tlb__T_624}; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@177587.4]
  assign tlb__T_631 = ~tlb_vm_enabled; // @[TLB.scala 213:18:freechips.rocketchip.system.DefaultRV32Config.fir@177588.4]
  assign tlb_hits = {tlb__T_631,tlb_hitsVec_12,tlb_hitsVec_11,tlb_hitsVec_10,tlb_hitsVec_9,tlb_hitsVec_8,tlb_hitsVec_7,tlb_hitsVec_6,tlb__T_624}; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@177589.4]
  assign tlb__GEN_33 = 2'h1 == tlb__T_510 ? tlb_sectored_entries_0_data_1 : tlb_sectored_entries_0_data_0; // @[:freechips.rocketchip.system.DefaultRV32Config.fir@177596.4]
  assign tlb__GEN_34 = 2'h2 == tlb__T_510 ? tlb_sectored_entries_0_data_2 : tlb__GEN_33; // @[:freechips.rocketchip.system.DefaultRV32Config.fir@177596.4]
  assign tlb__GEN_35 = 2'h3 == tlb__T_510 ? tlb_sectored_entries_0_data_3 : tlb__GEN_34; // @[:freechips.rocketchip.system.DefaultRV32Config.fir@177596.4]
  assign tlb__GEN_37 = 2'h1 == tlb__T_510 ? tlb_sectored_entries_1_data_1 : tlb_sectored_entries_1_data_0; // @[:freechips.rocketchip.system.DefaultRV32Config.fir@177639.4]
  assign tlb__GEN_38 = 2'h2 == tlb__T_510 ? tlb_sectored_entries_1_data_2 : tlb__GEN_37; // @[:freechips.rocketchip.system.DefaultRV32Config.fir@177639.4]
  assign tlb__GEN_39 = 2'h3 == tlb__T_510 ? tlb_sectored_entries_1_data_3 : tlb__GEN_38; // @[:freechips.rocketchip.system.DefaultRV32Config.fir@177639.4]
  assign tlb__GEN_41 = 2'h1 == tlb__T_510 ? tlb_sectored_entries_2_data_1 : tlb_sectored_entries_2_data_0; // @[:freechips.rocketchip.system.DefaultRV32Config.fir@177682.4]
  assign tlb__GEN_42 = 2'h2 == tlb__T_510 ? tlb_sectored_entries_2_data_2 : tlb__GEN_41; // @[:freechips.rocketchip.system.DefaultRV32Config.fir@177682.4]
  assign tlb__GEN_43 = 2'h3 == tlb__T_510 ? tlb_sectored_entries_2_data_3 : tlb__GEN_42; // @[:freechips.rocketchip.system.DefaultRV32Config.fir@177682.4]
  assign tlb__GEN_45 = 2'h1 == tlb__T_510 ? tlb_sectored_entries_3_data_1 : tlb_sectored_entries_3_data_0; // @[:freechips.rocketchip.system.DefaultRV32Config.fir@177725.4]
  assign tlb__GEN_46 = 2'h2 == tlb__T_510 ? tlb_sectored_entries_3_data_2 : tlb__GEN_45; // @[:freechips.rocketchip.system.DefaultRV32Config.fir@177725.4]
  assign tlb__GEN_47 = 2'h3 == tlb__T_510 ? tlb_sectored_entries_3_data_3 : tlb__GEN_46; // @[:freechips.rocketchip.system.DefaultRV32Config.fir@177725.4]
  assign tlb__GEN_49 = 2'h1 == tlb__T_510 ? tlb_sectored_entries_4_data_1 : tlb_sectored_entries_4_data_0; // @[:freechips.rocketchip.system.DefaultRV32Config.fir@177768.4]
  assign tlb__GEN_50 = 2'h2 == tlb__T_510 ? tlb_sectored_entries_4_data_2 : tlb__GEN_49; // @[:freechips.rocketchip.system.DefaultRV32Config.fir@177768.4]
  assign tlb__GEN_51 = 2'h3 == tlb__T_510 ? tlb_sectored_entries_4_data_3 : tlb__GEN_50; // @[:freechips.rocketchip.system.DefaultRV32Config.fir@177768.4]
  assign tlb__GEN_53 = 2'h1 == tlb__T_510 ? tlb_sectored_entries_5_data_1 : tlb_sectored_entries_5_data_0; // @[:freechips.rocketchip.system.DefaultRV32Config.fir@177811.4]
  assign tlb__GEN_54 = 2'h2 == tlb__T_510 ? tlb_sectored_entries_5_data_2 : tlb__GEN_53; // @[:freechips.rocketchip.system.DefaultRV32Config.fir@177811.4]
  assign tlb__GEN_55 = 2'h3 == tlb__T_510 ? tlb_sectored_entries_5_data_3 : tlb__GEN_54; // @[:freechips.rocketchip.system.DefaultRV32Config.fir@177811.4]
  assign tlb__GEN_57 = 2'h1 == tlb__T_510 ? tlb_sectored_entries_6_data_1 : tlb_sectored_entries_6_data_0; // @[:freechips.rocketchip.system.DefaultRV32Config.fir@177854.4]
  assign tlb__GEN_58 = 2'h2 == tlb__T_510 ? tlb_sectored_entries_6_data_2 : tlb__GEN_57; // @[:freechips.rocketchip.system.DefaultRV32Config.fir@177854.4]
  assign tlb__GEN_59 = 2'h3 == tlb__T_510 ? tlb_sectored_entries_6_data_3 : tlb__GEN_58; // @[:freechips.rocketchip.system.DefaultRV32Config.fir@177854.4]
  assign tlb__GEN_61 = 2'h1 == tlb__T_510 ? tlb_sectored_entries_7_data_1 : tlb_sectored_entries_7_data_0; // @[:freechips.rocketchip.system.DefaultRV32Config.fir@177897.4]
  assign tlb__GEN_62 = 2'h2 == tlb__T_510 ? tlb_sectored_entries_7_data_2 : tlb__GEN_61; // @[:freechips.rocketchip.system.DefaultRV32Config.fir@177897.4]
  assign tlb__GEN_63 = 2'h3 == tlb__T_510 ? tlb_sectored_entries_7_data_3 : tlb__GEN_62; // @[:freechips.rocketchip.system.DefaultRV32Config.fir@177897.4]
  assign tlb__T_800 = tlb_superpage_entries_0_data_0[13]; // @[TLB.scala 86:77:freechips.rocketchip.system.DefaultRV32Config.fir@177966.4]
  assign tlb__T_803 = tlb_OptimizationBarrier_9_io_y_ppn[19:10]; // @[TLB.scala 106:26:freechips.rocketchip.system.DefaultRV32Config.fir@177977.4]
  assign tlb__T_807 = tlb_vpn | tlb_OptimizationBarrier_9_io_y_ppn; // @[TLB.scala 109:47:freechips.rocketchip.system.DefaultRV32Config.fir@177981.4]
  assign tlb__T_808 = tlb__T_807[9:0]; // @[TLB.scala 109:58:freechips.rocketchip.system.DefaultRV32Config.fir@177982.4]
  assign tlb__T_809 = {tlb__T_803,tlb__T_808}; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@177983.4]
  assign tlb__T_825 = tlb_superpage_entries_1_data_0[13]; // @[TLB.scala 86:77:freechips.rocketchip.system.DefaultRV32Config.fir@178015.4]
  assign tlb__T_828 = tlb_OptimizationBarrier_10_io_y_ppn[19:10]; // @[TLB.scala 106:26:freechips.rocketchip.system.DefaultRV32Config.fir@178026.4]
  assign tlb__T_832 = tlb_vpn | tlb_OptimizationBarrier_10_io_y_ppn; // @[TLB.scala 109:47:freechips.rocketchip.system.DefaultRV32Config.fir@178030.4]
  assign tlb__T_833 = tlb__T_832[9:0]; // @[TLB.scala 109:58:freechips.rocketchip.system.DefaultRV32Config.fir@178031.4]
  assign tlb__T_834 = {tlb__T_828,tlb__T_833}; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@178032.4]
  assign tlb__T_850 = tlb_superpage_entries_2_data_0[13]; // @[TLB.scala 86:77:freechips.rocketchip.system.DefaultRV32Config.fir@178064.4]
  assign tlb__T_853 = tlb_OptimizationBarrier_11_io_y_ppn[19:10]; // @[TLB.scala 106:26:freechips.rocketchip.system.DefaultRV32Config.fir@178075.4]
  assign tlb__T_857 = tlb_vpn | tlb_OptimizationBarrier_11_io_y_ppn; // @[TLB.scala 109:47:freechips.rocketchip.system.DefaultRV32Config.fir@178079.4]
  assign tlb__T_858 = tlb__T_857[9:0]; // @[TLB.scala 109:58:freechips.rocketchip.system.DefaultRV32Config.fir@178080.4]
  assign tlb__T_859 = {tlb__T_853,tlb__T_858}; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@178081.4]
  assign tlb__T_875 = tlb_superpage_entries_3_data_0[13]; // @[TLB.scala 86:77:freechips.rocketchip.system.DefaultRV32Config.fir@178113.4]
  assign tlb__T_878 = tlb_OptimizationBarrier_12_io_y_ppn[19:10]; // @[TLB.scala 106:26:freechips.rocketchip.system.DefaultRV32Config.fir@178124.4]
  assign tlb__T_882 = tlb_vpn | tlb_OptimizationBarrier_12_io_y_ppn; // @[TLB.scala 109:47:freechips.rocketchip.system.DefaultRV32Config.fir@178128.4]
  assign tlb__T_883 = tlb__T_882[9:0]; // @[TLB.scala 109:58:freechips.rocketchip.system.DefaultRV32Config.fir@178129.4]
  assign tlb__T_884 = {tlb__T_878,tlb__T_883}; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@178130.4]
  assign tlb__T_903 = tlb_OptimizationBarrier_13_io_y_ppn[19:10]; // @[TLB.scala 106:26:freechips.rocketchip.system.DefaultRV32Config.fir@178173.4]
  assign tlb__T_907 = tlb__T_28 | tlb_OptimizationBarrier_13_io_y_ppn; // @[TLB.scala 109:47:freechips.rocketchip.system.DefaultRV32Config.fir@178177.4]
  assign tlb__T_908 = tlb__T_907[9:0]; // @[TLB.scala 109:58:freechips.rocketchip.system.DefaultRV32Config.fir@178178.4]
  assign tlb__T_909 = {tlb__T_903,tlb__T_908}; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@178179.4]
  assign tlb__T_911 = tlb_hitsVec_0 ? tlb_OptimizationBarrier_1_io_y_ppn : 20'h0; // @[Mux.scala 27:72:freechips.rocketchip.system.DefaultRV32Config.fir@178181.4]
  assign tlb__T_912 = tlb_hitsVec_1 ? tlb_OptimizationBarrier_2_io_y_ppn : 20'h0; // @[Mux.scala 27:72:freechips.rocketchip.system.DefaultRV32Config.fir@178182.4]
  assign tlb__T_913 = tlb_hitsVec_2 ? tlb_OptimizationBarrier_3_io_y_ppn : 20'h0; // @[Mux.scala 27:72:freechips.rocketchip.system.DefaultRV32Config.fir@178183.4]
  assign tlb__T_914 = tlb_hitsVec_3 ? tlb_OptimizationBarrier_4_io_y_ppn : 20'h0; // @[Mux.scala 27:72:freechips.rocketchip.system.DefaultRV32Config.fir@178184.4]
  assign tlb__T_915 = tlb_hitsVec_4 ? tlb_OptimizationBarrier_5_io_y_ppn : 20'h0; // @[Mux.scala 27:72:freechips.rocketchip.system.DefaultRV32Config.fir@178185.4]
  assign tlb__T_916 = tlb_hitsVec_5 ? tlb_OptimizationBarrier_6_io_y_ppn : 20'h0; // @[Mux.scala 27:72:freechips.rocketchip.system.DefaultRV32Config.fir@178186.4]
  assign tlb__T_917 = tlb_hitsVec_6 ? tlb_OptimizationBarrier_7_io_y_ppn : 20'h0; // @[Mux.scala 27:72:freechips.rocketchip.system.DefaultRV32Config.fir@178187.4]
  assign tlb__T_918 = tlb_hitsVec_7 ? tlb_OptimizationBarrier_8_io_y_ppn : 20'h0; // @[Mux.scala 27:72:freechips.rocketchip.system.DefaultRV32Config.fir@178188.4]
  assign tlb__T_919 = tlb_hitsVec_8 ? tlb__T_809 : 20'h0; // @[Mux.scala 27:72:freechips.rocketchip.system.DefaultRV32Config.fir@178189.4]
  assign tlb__T_920 = tlb_hitsVec_9 ? tlb__T_834 : 20'h0; // @[Mux.scala 27:72:freechips.rocketchip.system.DefaultRV32Config.fir@178190.4]
  assign tlb__T_921 = tlb_hitsVec_10 ? tlb__T_859 : 20'h0; // @[Mux.scala 27:72:freechips.rocketchip.system.DefaultRV32Config.fir@178191.4]
  assign tlb__T_922 = tlb_hitsVec_11 ? tlb__T_884 : 20'h0; // @[Mux.scala 27:72:freechips.rocketchip.system.DefaultRV32Config.fir@178192.4]
  assign tlb__T_923 = tlb_hitsVec_12 ? tlb__T_909 : 20'h0; // @[Mux.scala 27:72:freechips.rocketchip.system.DefaultRV32Config.fir@178193.4]
  assign tlb__T_924 = tlb__T_631 ? tlb_vpn : 20'h0; // @[Mux.scala 27:72:freechips.rocketchip.system.DefaultRV32Config.fir@178194.4]
  assign tlb__T_925 = tlb__T_911 | tlb__T_912; // @[Mux.scala 27:72:freechips.rocketchip.system.DefaultRV32Config.fir@178195.4]
  assign tlb__T_926 = tlb__T_925 | tlb__T_913; // @[Mux.scala 27:72:freechips.rocketchip.system.DefaultRV32Config.fir@178196.4]
  assign tlb__T_927 = tlb__T_926 | tlb__T_914; // @[Mux.scala 27:72:freechips.rocketchip.system.DefaultRV32Config.fir@178197.4]
  assign tlb__T_928 = tlb__T_927 | tlb__T_915; // @[Mux.scala 27:72:freechips.rocketchip.system.DefaultRV32Config.fir@178198.4]
  assign tlb__T_929 = tlb__T_928 | tlb__T_916; // @[Mux.scala 27:72:freechips.rocketchip.system.DefaultRV32Config.fir@178199.4]
  assign tlb__T_930 = tlb__T_929 | tlb__T_917; // @[Mux.scala 27:72:freechips.rocketchip.system.DefaultRV32Config.fir@178200.4]
  assign tlb__T_931 = tlb__T_930 | tlb__T_918; // @[Mux.scala 27:72:freechips.rocketchip.system.DefaultRV32Config.fir@178201.4]
  assign tlb__T_932 = tlb__T_931 | tlb__T_919; // @[Mux.scala 27:72:freechips.rocketchip.system.DefaultRV32Config.fir@178202.4]
  assign tlb__T_933 = tlb__T_932 | tlb__T_920; // @[Mux.scala 27:72:freechips.rocketchip.system.DefaultRV32Config.fir@178203.4]
  assign tlb__T_934 = tlb__T_933 | tlb__T_921; // @[Mux.scala 27:72:freechips.rocketchip.system.DefaultRV32Config.fir@178204.4]
  assign tlb__T_935 = tlb__T_934 | tlb__T_922; // @[Mux.scala 27:72:freechips.rocketchip.system.DefaultRV32Config.fir@178205.4]
  assign tlb__T_936 = tlb__T_935 | tlb__T_923; // @[Mux.scala 27:72:freechips.rocketchip.system.DefaultRV32Config.fir@178206.4]
  assign tlb__T_937 = tlb__T_936 | tlb__T_924; // @[Mux.scala 27:72:freechips.rocketchip.system.DefaultRV32Config.fir@178207.4]
  assign tlb__T_938 = ~tlb_invalidate_refill; // @[TLB.scala 217:22:freechips.rocketchip.system.DefaultRV32Config.fir@178210.4]
  assign tlb__T_939 = tlb_io_ptw_resp_valid & tlb__T_938; // @[TLB.scala 217:19:freechips.rocketchip.system.DefaultRV32Config.fir@178211.4]
  assign tlb__T_941 = tlb_io_ptw_resp_bits_pte_g & tlb_io_ptw_resp_bits_pte_v; // @[TLB.scala 223:25:freechips.rocketchip.system.DefaultRV32Config.fir@178218.6]
  assign tlb__T_942 = ~tlb_io_ptw_resp_bits_pte_w; // @[PTW.scala 69:47:freechips.rocketchip.system.DefaultRV32Config.fir@178221.6]
  assign tlb__T_943 = tlb_io_ptw_resp_bits_pte_x & tlb__T_942; // @[PTW.scala 69:44:freechips.rocketchip.system.DefaultRV32Config.fir@178222.6]
  assign tlb__T_944 = tlb_io_ptw_resp_bits_pte_r | tlb__T_943; // @[PTW.scala 69:38:freechips.rocketchip.system.DefaultRV32Config.fir@178223.6]
  assign tlb__T_945 = tlb_io_ptw_resp_bits_pte_v & tlb__T_944; // @[PTW.scala 69:32:freechips.rocketchip.system.DefaultRV32Config.fir@178224.6]
  assign tlb__T_946 = tlb__T_945 & tlb_io_ptw_resp_bits_pte_a; // @[PTW.scala 69:52:freechips.rocketchip.system.DefaultRV32Config.fir@178225.6]
  assign tlb__T_947 = tlb__T_946 & tlb_io_ptw_resp_bits_pte_r; // @[PTW.scala 73:35:freechips.rocketchip.system.DefaultRV32Config.fir@178226.6]
  assign tlb__T_953 = tlb__T_946 & tlb_io_ptw_resp_bits_pte_w; // @[PTW.scala 74:35:freechips.rocketchip.system.DefaultRV32Config.fir@178233.6]
  assign tlb__T_954 = tlb__T_953 & tlb_io_ptw_resp_bits_pte_d; // @[PTW.scala 74:40:freechips.rocketchip.system.DefaultRV32Config.fir@178234.6]
  assign tlb__T_960 = tlb__T_946 & tlb_io_ptw_resp_bits_pte_x; // @[PTW.scala 75:35:freechips.rocketchip.system.DefaultRV32Config.fir@178241.6]
  assign tlb__T_961 = ~tlb_io_ptw_resp_bits_homogeneous; // @[TLB.scala 237:37:freechips.rocketchip.system.DefaultRV32Config.fir@178251.6]
  assign tlb__T_970 = {tlb_prot_x,tlb_prot_r,tlb__T_232,tlb_prot_al,tlb_prot_al,tlb_prot_eff,tlb__T_93,1'h0}; // @[TLB.scala 123:24:freechips.rocketchip.system.DefaultRV32Config.fir@178264.8]
  assign tlb__T_978 = {tlb_refill_ppn,tlb_io_ptw_resp_bits_pte_u,tlb__T_941,tlb_io_ptw_resp_bits_ae,tlb__T_954,tlb__T_960,tlb__T_947,tlb_prot_w,tlb__T_970}; // @[TLB.scala 123:24:freechips.rocketchip.system.DefaultRV32Config.fir@178272.8]
  assign tlb__T_979 = tlb_io_ptw_resp_bits_level < 1'h1; // @[TLB.scala 239:40:freechips.rocketchip.system.DefaultRV32Config.fir@178276.8]
  assign tlb__T_980 = tlb_r_superpage_repl_addr == 2'h0; // @[TLB.scala 240:82:freechips.rocketchip.system.DefaultRV32Config.fir@178278.10]
  assign tlb__GEN_66 = tlb__T_980 | tlb_superpage_entries_0_valid_0; // @[TLB.scala 240:89:freechips.rocketchip.system.DefaultRV32Config.fir@178279.10]
  assign tlb__T_996 = tlb_r_superpage_repl_addr == 2'h1; // @[TLB.scala 240:82:freechips.rocketchip.system.DefaultRV32Config.fir@178300.10]
  assign tlb__GEN_70 = tlb__T_996 | tlb_superpage_entries_1_valid_0; // @[TLB.scala 240:89:freechips.rocketchip.system.DefaultRV32Config.fir@178301.10]
  assign tlb__T_1012 = tlb_r_superpage_repl_addr == 2'h2; // @[TLB.scala 240:82:freechips.rocketchip.system.DefaultRV32Config.fir@178322.10]
  assign tlb__GEN_74 = tlb__T_1012 | tlb_superpage_entries_2_valid_0; // @[TLB.scala 240:89:freechips.rocketchip.system.DefaultRV32Config.fir@178323.10]
  assign tlb__T_1028 = tlb_r_superpage_repl_addr == 2'h3; // @[TLB.scala 240:82:freechips.rocketchip.system.DefaultRV32Config.fir@178344.10]
  assign tlb__GEN_78 = tlb__T_1028 | tlb_superpage_entries_3_valid_0; // @[TLB.scala 240:89:freechips.rocketchip.system.DefaultRV32Config.fir@178345.10]
  assign tlb__T_1044 = tlb_r_sectored_hit ? tlb_r_sectored_hit_addr : tlb_r_sectored_repl_addr; // @[TLB.scala 244:22:freechips.rocketchip.system.DefaultRV32Config.fir@178368.10]
  assign tlb__T_1045 = tlb__T_1044 == 3'h0; // @[TLB.scala 245:65:freechips.rocketchip.system.DefaultRV32Config.fir@178369.10]
  assign tlb__T_1046 = ~tlb_r_sectored_hit; // @[TLB.scala 246:15:freechips.rocketchip.system.DefaultRV32Config.fir@178371.12]
  assign tlb__GEN_80 = tlb__T_1046 ? 1'h0 : tlb_sectored_entries_0_valid_0; // @[TLB.scala 246:32:freechips.rocketchip.system.DefaultRV32Config.fir@178372.12]
  assign tlb__GEN_81 = tlb__T_1046 ? 1'h0 : tlb_sectored_entries_0_valid_1; // @[TLB.scala 246:32:freechips.rocketchip.system.DefaultRV32Config.fir@178372.12]
  assign tlb__GEN_82 = tlb__T_1046 ? 1'h0 : tlb_sectored_entries_0_valid_2; // @[TLB.scala 246:32:freechips.rocketchip.system.DefaultRV32Config.fir@178372.12]
  assign tlb__GEN_83 = tlb__T_1046 ? 1'h0 : tlb_sectored_entries_0_valid_3; // @[TLB.scala 246:32:freechips.rocketchip.system.DefaultRV32Config.fir@178372.12]
  assign tlb__T_1047 = tlb_r_refill_tag[1:0]; // @[package.scala 138:13:freechips.rocketchip.system.DefaultRV32Config.fir@178380.12]
  assign _GEN_343 = 2'h0 == tlb__T_1047; // @[TLB.scala 122:16:freechips.rocketchip.system.DefaultRV32Config.fir@178381.12]
  assign tlb__GEN_84 = _GEN_343 | tlb__GEN_80; // @[TLB.scala 122:16:freechips.rocketchip.system.DefaultRV32Config.fir@178381.12]
  assign _GEN_344 = 2'h1 == tlb__T_1047; // @[TLB.scala 122:16:freechips.rocketchip.system.DefaultRV32Config.fir@178381.12]
  assign tlb__GEN_85 = _GEN_344 | tlb__GEN_81; // @[TLB.scala 122:16:freechips.rocketchip.system.DefaultRV32Config.fir@178381.12]
  assign _GEN_345 = 2'h2 == tlb__T_1047; // @[TLB.scala 122:16:freechips.rocketchip.system.DefaultRV32Config.fir@178381.12]
  assign tlb__GEN_86 = _GEN_345 | tlb__GEN_82; // @[TLB.scala 122:16:freechips.rocketchip.system.DefaultRV32Config.fir@178381.12]
  assign _GEN_346 = 2'h3 == tlb__T_1047; // @[TLB.scala 122:16:freechips.rocketchip.system.DefaultRV32Config.fir@178381.12]
  assign tlb__GEN_87 = _GEN_346 | tlb__GEN_83; // @[TLB.scala 122:16:freechips.rocketchip.system.DefaultRV32Config.fir@178381.12]
  assign tlb__GEN_92 = tlb__T_1045 ? tlb__GEN_84 : tlb_sectored_entries_0_valid_0; // @[TLB.scala 245:72:freechips.rocketchip.system.DefaultRV32Config.fir@178370.10]
  assign tlb__GEN_93 = tlb__T_1045 ? tlb__GEN_85 : tlb_sectored_entries_0_valid_1; // @[TLB.scala 245:72:freechips.rocketchip.system.DefaultRV32Config.fir@178370.10]
  assign tlb__GEN_94 = tlb__T_1045 ? tlb__GEN_86 : tlb_sectored_entries_0_valid_2; // @[TLB.scala 245:72:freechips.rocketchip.system.DefaultRV32Config.fir@178370.10]
  assign tlb__GEN_95 = tlb__T_1045 ? tlb__GEN_87 : tlb_sectored_entries_0_valid_3; // @[TLB.scala 245:72:freechips.rocketchip.system.DefaultRV32Config.fir@178370.10]
  assign tlb__T_1063 = tlb__T_1044 == 3'h1; // @[TLB.scala 245:65:freechips.rocketchip.system.DefaultRV32Config.fir@178399.10]
  assign tlb__GEN_102 = tlb__T_1046 ? 1'h0 : tlb_sectored_entries_1_valid_0; // @[TLB.scala 246:32:freechips.rocketchip.system.DefaultRV32Config.fir@178402.12]
  assign tlb__GEN_103 = tlb__T_1046 ? 1'h0 : tlb_sectored_entries_1_valid_1; // @[TLB.scala 246:32:freechips.rocketchip.system.DefaultRV32Config.fir@178402.12]
  assign tlb__GEN_104 = tlb__T_1046 ? 1'h0 : tlb_sectored_entries_1_valid_2; // @[TLB.scala 246:32:freechips.rocketchip.system.DefaultRV32Config.fir@178402.12]
  assign tlb__GEN_105 = tlb__T_1046 ? 1'h0 : tlb_sectored_entries_1_valid_3; // @[TLB.scala 246:32:freechips.rocketchip.system.DefaultRV32Config.fir@178402.12]
  assign tlb__GEN_106 = _GEN_343 | tlb__GEN_102; // @[TLB.scala 122:16:freechips.rocketchip.system.DefaultRV32Config.fir@178411.12]
  assign tlb__GEN_107 = _GEN_344 | tlb__GEN_103; // @[TLB.scala 122:16:freechips.rocketchip.system.DefaultRV32Config.fir@178411.12]
  assign tlb__GEN_108 = _GEN_345 | tlb__GEN_104; // @[TLB.scala 122:16:freechips.rocketchip.system.DefaultRV32Config.fir@178411.12]
  assign tlb__GEN_109 = _GEN_346 | tlb__GEN_105; // @[TLB.scala 122:16:freechips.rocketchip.system.DefaultRV32Config.fir@178411.12]
  assign tlb__GEN_114 = tlb__T_1063 ? tlb__GEN_106 : tlb_sectored_entries_1_valid_0; // @[TLB.scala 245:72:freechips.rocketchip.system.DefaultRV32Config.fir@178400.10]
  assign tlb__GEN_115 = tlb__T_1063 ? tlb__GEN_107 : tlb_sectored_entries_1_valid_1; // @[TLB.scala 245:72:freechips.rocketchip.system.DefaultRV32Config.fir@178400.10]
  assign tlb__GEN_116 = tlb__T_1063 ? tlb__GEN_108 : tlb_sectored_entries_1_valid_2; // @[TLB.scala 245:72:freechips.rocketchip.system.DefaultRV32Config.fir@178400.10]
  assign tlb__GEN_117 = tlb__T_1063 ? tlb__GEN_109 : tlb_sectored_entries_1_valid_3; // @[TLB.scala 245:72:freechips.rocketchip.system.DefaultRV32Config.fir@178400.10]
  assign tlb__T_1081 = tlb__T_1044 == 3'h2; // @[TLB.scala 245:65:freechips.rocketchip.system.DefaultRV32Config.fir@178429.10]
  assign tlb__GEN_124 = tlb__T_1046 ? 1'h0 : tlb_sectored_entries_2_valid_0; // @[TLB.scala 246:32:freechips.rocketchip.system.DefaultRV32Config.fir@178432.12]
  assign tlb__GEN_125 = tlb__T_1046 ? 1'h0 : tlb_sectored_entries_2_valid_1; // @[TLB.scala 246:32:freechips.rocketchip.system.DefaultRV32Config.fir@178432.12]
  assign tlb__GEN_126 = tlb__T_1046 ? 1'h0 : tlb_sectored_entries_2_valid_2; // @[TLB.scala 246:32:freechips.rocketchip.system.DefaultRV32Config.fir@178432.12]
  assign tlb__GEN_127 = tlb__T_1046 ? 1'h0 : tlb_sectored_entries_2_valid_3; // @[TLB.scala 246:32:freechips.rocketchip.system.DefaultRV32Config.fir@178432.12]
  assign tlb__GEN_128 = _GEN_343 | tlb__GEN_124; // @[TLB.scala 122:16:freechips.rocketchip.system.DefaultRV32Config.fir@178441.12]
  assign tlb__GEN_129 = _GEN_344 | tlb__GEN_125; // @[TLB.scala 122:16:freechips.rocketchip.system.DefaultRV32Config.fir@178441.12]
  assign tlb__GEN_130 = _GEN_345 | tlb__GEN_126; // @[TLB.scala 122:16:freechips.rocketchip.system.DefaultRV32Config.fir@178441.12]
  assign tlb__GEN_131 = _GEN_346 | tlb__GEN_127; // @[TLB.scala 122:16:freechips.rocketchip.system.DefaultRV32Config.fir@178441.12]
  assign tlb__GEN_136 = tlb__T_1081 ? tlb__GEN_128 : tlb_sectored_entries_2_valid_0; // @[TLB.scala 245:72:freechips.rocketchip.system.DefaultRV32Config.fir@178430.10]
  assign tlb__GEN_137 = tlb__T_1081 ? tlb__GEN_129 : tlb_sectored_entries_2_valid_1; // @[TLB.scala 245:72:freechips.rocketchip.system.DefaultRV32Config.fir@178430.10]
  assign tlb__GEN_138 = tlb__T_1081 ? tlb__GEN_130 : tlb_sectored_entries_2_valid_2; // @[TLB.scala 245:72:freechips.rocketchip.system.DefaultRV32Config.fir@178430.10]
  assign tlb__GEN_139 = tlb__T_1081 ? tlb__GEN_131 : tlb_sectored_entries_2_valid_3; // @[TLB.scala 245:72:freechips.rocketchip.system.DefaultRV32Config.fir@178430.10]
  assign tlb__T_1099 = tlb__T_1044 == 3'h3; // @[TLB.scala 245:65:freechips.rocketchip.system.DefaultRV32Config.fir@178459.10]
  assign tlb__GEN_146 = tlb__T_1046 ? 1'h0 : tlb_sectored_entries_3_valid_0; // @[TLB.scala 246:32:freechips.rocketchip.system.DefaultRV32Config.fir@178462.12]
  assign tlb__GEN_147 = tlb__T_1046 ? 1'h0 : tlb_sectored_entries_3_valid_1; // @[TLB.scala 246:32:freechips.rocketchip.system.DefaultRV32Config.fir@178462.12]
  assign tlb__GEN_148 = tlb__T_1046 ? 1'h0 : tlb_sectored_entries_3_valid_2; // @[TLB.scala 246:32:freechips.rocketchip.system.DefaultRV32Config.fir@178462.12]
  assign tlb__GEN_149 = tlb__T_1046 ? 1'h0 : tlb_sectored_entries_3_valid_3; // @[TLB.scala 246:32:freechips.rocketchip.system.DefaultRV32Config.fir@178462.12]
  assign tlb__GEN_150 = _GEN_343 | tlb__GEN_146; // @[TLB.scala 122:16:freechips.rocketchip.system.DefaultRV32Config.fir@178471.12]
  assign tlb__GEN_151 = _GEN_344 | tlb__GEN_147; // @[TLB.scala 122:16:freechips.rocketchip.system.DefaultRV32Config.fir@178471.12]
  assign tlb__GEN_152 = _GEN_345 | tlb__GEN_148; // @[TLB.scala 122:16:freechips.rocketchip.system.DefaultRV32Config.fir@178471.12]
  assign tlb__GEN_153 = _GEN_346 | tlb__GEN_149; // @[TLB.scala 122:16:freechips.rocketchip.system.DefaultRV32Config.fir@178471.12]
  assign tlb__GEN_158 = tlb__T_1099 ? tlb__GEN_150 : tlb_sectored_entries_3_valid_0; // @[TLB.scala 245:72:freechips.rocketchip.system.DefaultRV32Config.fir@178460.10]
  assign tlb__GEN_159 = tlb__T_1099 ? tlb__GEN_151 : tlb_sectored_entries_3_valid_1; // @[TLB.scala 245:72:freechips.rocketchip.system.DefaultRV32Config.fir@178460.10]
  assign tlb__GEN_160 = tlb__T_1099 ? tlb__GEN_152 : tlb_sectored_entries_3_valid_2; // @[TLB.scala 245:72:freechips.rocketchip.system.DefaultRV32Config.fir@178460.10]
  assign tlb__GEN_161 = tlb__T_1099 ? tlb__GEN_153 : tlb_sectored_entries_3_valid_3; // @[TLB.scala 245:72:freechips.rocketchip.system.DefaultRV32Config.fir@178460.10]
  assign tlb__T_1117 = tlb__T_1044 == 3'h4; // @[TLB.scala 245:65:freechips.rocketchip.system.DefaultRV32Config.fir@178489.10]
  assign tlb__GEN_168 = tlb__T_1046 ? 1'h0 : tlb_sectored_entries_4_valid_0; // @[TLB.scala 246:32:freechips.rocketchip.system.DefaultRV32Config.fir@178492.12]
  assign tlb__GEN_169 = tlb__T_1046 ? 1'h0 : tlb_sectored_entries_4_valid_1; // @[TLB.scala 246:32:freechips.rocketchip.system.DefaultRV32Config.fir@178492.12]
  assign tlb__GEN_170 = tlb__T_1046 ? 1'h0 : tlb_sectored_entries_4_valid_2; // @[TLB.scala 246:32:freechips.rocketchip.system.DefaultRV32Config.fir@178492.12]
  assign tlb__GEN_171 = tlb__T_1046 ? 1'h0 : tlb_sectored_entries_4_valid_3; // @[TLB.scala 246:32:freechips.rocketchip.system.DefaultRV32Config.fir@178492.12]
  assign tlb__GEN_172 = _GEN_343 | tlb__GEN_168; // @[TLB.scala 122:16:freechips.rocketchip.system.DefaultRV32Config.fir@178501.12]
  assign tlb__GEN_173 = _GEN_344 | tlb__GEN_169; // @[TLB.scala 122:16:freechips.rocketchip.system.DefaultRV32Config.fir@178501.12]
  assign tlb__GEN_174 = _GEN_345 | tlb__GEN_170; // @[TLB.scala 122:16:freechips.rocketchip.system.DefaultRV32Config.fir@178501.12]
  assign tlb__GEN_175 = _GEN_346 | tlb__GEN_171; // @[TLB.scala 122:16:freechips.rocketchip.system.DefaultRV32Config.fir@178501.12]
  assign tlb__GEN_180 = tlb__T_1117 ? tlb__GEN_172 : tlb_sectored_entries_4_valid_0; // @[TLB.scala 245:72:freechips.rocketchip.system.DefaultRV32Config.fir@178490.10]
  assign tlb__GEN_181 = tlb__T_1117 ? tlb__GEN_173 : tlb_sectored_entries_4_valid_1; // @[TLB.scala 245:72:freechips.rocketchip.system.DefaultRV32Config.fir@178490.10]
  assign tlb__GEN_182 = tlb__T_1117 ? tlb__GEN_174 : tlb_sectored_entries_4_valid_2; // @[TLB.scala 245:72:freechips.rocketchip.system.DefaultRV32Config.fir@178490.10]
  assign tlb__GEN_183 = tlb__T_1117 ? tlb__GEN_175 : tlb_sectored_entries_4_valid_3; // @[TLB.scala 245:72:freechips.rocketchip.system.DefaultRV32Config.fir@178490.10]
  assign tlb__T_1135 = tlb__T_1044 == 3'h5; // @[TLB.scala 245:65:freechips.rocketchip.system.DefaultRV32Config.fir@178519.10]
  assign tlb__GEN_190 = tlb__T_1046 ? 1'h0 : tlb_sectored_entries_5_valid_0; // @[TLB.scala 246:32:freechips.rocketchip.system.DefaultRV32Config.fir@178522.12]
  assign tlb__GEN_191 = tlb__T_1046 ? 1'h0 : tlb_sectored_entries_5_valid_1; // @[TLB.scala 246:32:freechips.rocketchip.system.DefaultRV32Config.fir@178522.12]
  assign tlb__GEN_192 = tlb__T_1046 ? 1'h0 : tlb_sectored_entries_5_valid_2; // @[TLB.scala 246:32:freechips.rocketchip.system.DefaultRV32Config.fir@178522.12]
  assign tlb__GEN_193 = tlb__T_1046 ? 1'h0 : tlb_sectored_entries_5_valid_3; // @[TLB.scala 246:32:freechips.rocketchip.system.DefaultRV32Config.fir@178522.12]
  assign tlb__GEN_194 = _GEN_343 | tlb__GEN_190; // @[TLB.scala 122:16:freechips.rocketchip.system.DefaultRV32Config.fir@178531.12]
  assign tlb__GEN_195 = _GEN_344 | tlb__GEN_191; // @[TLB.scala 122:16:freechips.rocketchip.system.DefaultRV32Config.fir@178531.12]
  assign tlb__GEN_196 = _GEN_345 | tlb__GEN_192; // @[TLB.scala 122:16:freechips.rocketchip.system.DefaultRV32Config.fir@178531.12]
  assign tlb__GEN_197 = _GEN_346 | tlb__GEN_193; // @[TLB.scala 122:16:freechips.rocketchip.system.DefaultRV32Config.fir@178531.12]
  assign tlb__GEN_202 = tlb__T_1135 ? tlb__GEN_194 : tlb_sectored_entries_5_valid_0; // @[TLB.scala 245:72:freechips.rocketchip.system.DefaultRV32Config.fir@178520.10]
  assign tlb__GEN_203 = tlb__T_1135 ? tlb__GEN_195 : tlb_sectored_entries_5_valid_1; // @[TLB.scala 245:72:freechips.rocketchip.system.DefaultRV32Config.fir@178520.10]
  assign tlb__GEN_204 = tlb__T_1135 ? tlb__GEN_196 : tlb_sectored_entries_5_valid_2; // @[TLB.scala 245:72:freechips.rocketchip.system.DefaultRV32Config.fir@178520.10]
  assign tlb__GEN_205 = tlb__T_1135 ? tlb__GEN_197 : tlb_sectored_entries_5_valid_3; // @[TLB.scala 245:72:freechips.rocketchip.system.DefaultRV32Config.fir@178520.10]
  assign tlb__T_1153 = tlb__T_1044 == 3'h6; // @[TLB.scala 245:65:freechips.rocketchip.system.DefaultRV32Config.fir@178549.10]
  assign tlb__GEN_212 = tlb__T_1046 ? 1'h0 : tlb_sectored_entries_6_valid_0; // @[TLB.scala 246:32:freechips.rocketchip.system.DefaultRV32Config.fir@178552.12]
  assign tlb__GEN_213 = tlb__T_1046 ? 1'h0 : tlb_sectored_entries_6_valid_1; // @[TLB.scala 246:32:freechips.rocketchip.system.DefaultRV32Config.fir@178552.12]
  assign tlb__GEN_214 = tlb__T_1046 ? 1'h0 : tlb_sectored_entries_6_valid_2; // @[TLB.scala 246:32:freechips.rocketchip.system.DefaultRV32Config.fir@178552.12]
  assign tlb__GEN_215 = tlb__T_1046 ? 1'h0 : tlb_sectored_entries_6_valid_3; // @[TLB.scala 246:32:freechips.rocketchip.system.DefaultRV32Config.fir@178552.12]
  assign tlb__GEN_216 = _GEN_343 | tlb__GEN_212; // @[TLB.scala 122:16:freechips.rocketchip.system.DefaultRV32Config.fir@178561.12]
  assign tlb__GEN_217 = _GEN_344 | tlb__GEN_213; // @[TLB.scala 122:16:freechips.rocketchip.system.DefaultRV32Config.fir@178561.12]
  assign tlb__GEN_218 = _GEN_345 | tlb__GEN_214; // @[TLB.scala 122:16:freechips.rocketchip.system.DefaultRV32Config.fir@178561.12]
  assign tlb__GEN_219 = _GEN_346 | tlb__GEN_215; // @[TLB.scala 122:16:freechips.rocketchip.system.DefaultRV32Config.fir@178561.12]
  assign tlb__GEN_224 = tlb__T_1153 ? tlb__GEN_216 : tlb_sectored_entries_6_valid_0; // @[TLB.scala 245:72:freechips.rocketchip.system.DefaultRV32Config.fir@178550.10]
  assign tlb__GEN_225 = tlb__T_1153 ? tlb__GEN_217 : tlb_sectored_entries_6_valid_1; // @[TLB.scala 245:72:freechips.rocketchip.system.DefaultRV32Config.fir@178550.10]
  assign tlb__GEN_226 = tlb__T_1153 ? tlb__GEN_218 : tlb_sectored_entries_6_valid_2; // @[TLB.scala 245:72:freechips.rocketchip.system.DefaultRV32Config.fir@178550.10]
  assign tlb__GEN_227 = tlb__T_1153 ? tlb__GEN_219 : tlb_sectored_entries_6_valid_3; // @[TLB.scala 245:72:freechips.rocketchip.system.DefaultRV32Config.fir@178550.10]
  assign tlb__T_1171 = tlb__T_1044 == 3'h7; // @[TLB.scala 245:65:freechips.rocketchip.system.DefaultRV32Config.fir@178579.10]
  assign tlb__GEN_234 = tlb__T_1046 ? 1'h0 : tlb_sectored_entries_7_valid_0; // @[TLB.scala 246:32:freechips.rocketchip.system.DefaultRV32Config.fir@178582.12]
  assign tlb__GEN_235 = tlb__T_1046 ? 1'h0 : tlb_sectored_entries_7_valid_1; // @[TLB.scala 246:32:freechips.rocketchip.system.DefaultRV32Config.fir@178582.12]
  assign tlb__GEN_236 = tlb__T_1046 ? 1'h0 : tlb_sectored_entries_7_valid_2; // @[TLB.scala 246:32:freechips.rocketchip.system.DefaultRV32Config.fir@178582.12]
  assign tlb__GEN_237 = tlb__T_1046 ? 1'h0 : tlb_sectored_entries_7_valid_3; // @[TLB.scala 246:32:freechips.rocketchip.system.DefaultRV32Config.fir@178582.12]
  assign tlb__GEN_238 = _GEN_343 | tlb__GEN_234; // @[TLB.scala 122:16:freechips.rocketchip.system.DefaultRV32Config.fir@178591.12]
  assign tlb__GEN_239 = _GEN_344 | tlb__GEN_235; // @[TLB.scala 122:16:freechips.rocketchip.system.DefaultRV32Config.fir@178591.12]
  assign tlb__GEN_240 = _GEN_345 | tlb__GEN_236; // @[TLB.scala 122:16:freechips.rocketchip.system.DefaultRV32Config.fir@178591.12]
  assign tlb__GEN_241 = _GEN_346 | tlb__GEN_237; // @[TLB.scala 122:16:freechips.rocketchip.system.DefaultRV32Config.fir@178591.12]
  assign tlb__GEN_246 = tlb__T_1171 ? tlb__GEN_238 : tlb_sectored_entries_7_valid_0; // @[TLB.scala 245:72:freechips.rocketchip.system.DefaultRV32Config.fir@178580.10]
  assign tlb__GEN_247 = tlb__T_1171 ? tlb__GEN_239 : tlb_sectored_entries_7_valid_1; // @[TLB.scala 245:72:freechips.rocketchip.system.DefaultRV32Config.fir@178580.10]
  assign tlb__GEN_248 = tlb__T_1171 ? tlb__GEN_240 : tlb_sectored_entries_7_valid_2; // @[TLB.scala 245:72:freechips.rocketchip.system.DefaultRV32Config.fir@178580.10]
  assign tlb__GEN_249 = tlb__T_1171 ? tlb__GEN_241 : tlb_sectored_entries_7_valid_3; // @[TLB.scala 245:72:freechips.rocketchip.system.DefaultRV32Config.fir@178580.10]
  assign tlb__GEN_258 = tlb__T_979 ? tlb__GEN_66 : tlb_superpage_entries_0_valid_0; // @[TLB.scala 239:54:freechips.rocketchip.system.DefaultRV32Config.fir@178277.8]
  assign tlb__GEN_262 = tlb__T_979 ? tlb__GEN_70 : tlb_superpage_entries_1_valid_0; // @[TLB.scala 239:54:freechips.rocketchip.system.DefaultRV32Config.fir@178277.8]
  assign tlb__GEN_266 = tlb__T_979 ? tlb__GEN_74 : tlb_superpage_entries_2_valid_0; // @[TLB.scala 239:54:freechips.rocketchip.system.DefaultRV32Config.fir@178277.8]
  assign tlb__GEN_270 = tlb__T_979 ? tlb__GEN_78 : tlb_superpage_entries_3_valid_0; // @[TLB.scala 239:54:freechips.rocketchip.system.DefaultRV32Config.fir@178277.8]
  assign tlb__GEN_272 = tlb__T_979 ? tlb_sectored_entries_0_valid_0 : tlb__GEN_92; // @[TLB.scala 239:54:freechips.rocketchip.system.DefaultRV32Config.fir@178277.8]
  assign tlb__GEN_273 = tlb__T_979 ? tlb_sectored_entries_0_valid_1 : tlb__GEN_93; // @[TLB.scala 239:54:freechips.rocketchip.system.DefaultRV32Config.fir@178277.8]
  assign tlb__GEN_274 = tlb__T_979 ? tlb_sectored_entries_0_valid_2 : tlb__GEN_94; // @[TLB.scala 239:54:freechips.rocketchip.system.DefaultRV32Config.fir@178277.8]
  assign tlb__GEN_275 = tlb__T_979 ? tlb_sectored_entries_0_valid_3 : tlb__GEN_95; // @[TLB.scala 239:54:freechips.rocketchip.system.DefaultRV32Config.fir@178277.8]
  assign tlb__GEN_282 = tlb__T_979 ? tlb_sectored_entries_1_valid_0 : tlb__GEN_114; // @[TLB.scala 239:54:freechips.rocketchip.system.DefaultRV32Config.fir@178277.8]
  assign tlb__GEN_283 = tlb__T_979 ? tlb_sectored_entries_1_valid_1 : tlb__GEN_115; // @[TLB.scala 239:54:freechips.rocketchip.system.DefaultRV32Config.fir@178277.8]
  assign tlb__GEN_284 = tlb__T_979 ? tlb_sectored_entries_1_valid_2 : tlb__GEN_116; // @[TLB.scala 239:54:freechips.rocketchip.system.DefaultRV32Config.fir@178277.8]
  assign tlb__GEN_285 = tlb__T_979 ? tlb_sectored_entries_1_valid_3 : tlb__GEN_117; // @[TLB.scala 239:54:freechips.rocketchip.system.DefaultRV32Config.fir@178277.8]
  assign tlb__GEN_292 = tlb__T_979 ? tlb_sectored_entries_2_valid_0 : tlb__GEN_136; // @[TLB.scala 239:54:freechips.rocketchip.system.DefaultRV32Config.fir@178277.8]
  assign tlb__GEN_293 = tlb__T_979 ? tlb_sectored_entries_2_valid_1 : tlb__GEN_137; // @[TLB.scala 239:54:freechips.rocketchip.system.DefaultRV32Config.fir@178277.8]
  assign tlb__GEN_294 = tlb__T_979 ? tlb_sectored_entries_2_valid_2 : tlb__GEN_138; // @[TLB.scala 239:54:freechips.rocketchip.system.DefaultRV32Config.fir@178277.8]
  assign tlb__GEN_295 = tlb__T_979 ? tlb_sectored_entries_2_valid_3 : tlb__GEN_139; // @[TLB.scala 239:54:freechips.rocketchip.system.DefaultRV32Config.fir@178277.8]
  assign tlb__GEN_302 = tlb__T_979 ? tlb_sectored_entries_3_valid_0 : tlb__GEN_158; // @[TLB.scala 239:54:freechips.rocketchip.system.DefaultRV32Config.fir@178277.8]
  assign tlb__GEN_303 = tlb__T_979 ? tlb_sectored_entries_3_valid_1 : tlb__GEN_159; // @[TLB.scala 239:54:freechips.rocketchip.system.DefaultRV32Config.fir@178277.8]
  assign tlb__GEN_304 = tlb__T_979 ? tlb_sectored_entries_3_valid_2 : tlb__GEN_160; // @[TLB.scala 239:54:freechips.rocketchip.system.DefaultRV32Config.fir@178277.8]
  assign tlb__GEN_305 = tlb__T_979 ? tlb_sectored_entries_3_valid_3 : tlb__GEN_161; // @[TLB.scala 239:54:freechips.rocketchip.system.DefaultRV32Config.fir@178277.8]
  assign tlb__GEN_312 = tlb__T_979 ? tlb_sectored_entries_4_valid_0 : tlb__GEN_180; // @[TLB.scala 239:54:freechips.rocketchip.system.DefaultRV32Config.fir@178277.8]
  assign tlb__GEN_313 = tlb__T_979 ? tlb_sectored_entries_4_valid_1 : tlb__GEN_181; // @[TLB.scala 239:54:freechips.rocketchip.system.DefaultRV32Config.fir@178277.8]
  assign tlb__GEN_314 = tlb__T_979 ? tlb_sectored_entries_4_valid_2 : tlb__GEN_182; // @[TLB.scala 239:54:freechips.rocketchip.system.DefaultRV32Config.fir@178277.8]
  assign tlb__GEN_315 = tlb__T_979 ? tlb_sectored_entries_4_valid_3 : tlb__GEN_183; // @[TLB.scala 239:54:freechips.rocketchip.system.DefaultRV32Config.fir@178277.8]
  assign tlb__GEN_322 = tlb__T_979 ? tlb_sectored_entries_5_valid_0 : tlb__GEN_202; // @[TLB.scala 239:54:freechips.rocketchip.system.DefaultRV32Config.fir@178277.8]
  assign tlb__GEN_323 = tlb__T_979 ? tlb_sectored_entries_5_valid_1 : tlb__GEN_203; // @[TLB.scala 239:54:freechips.rocketchip.system.DefaultRV32Config.fir@178277.8]
  assign tlb__GEN_324 = tlb__T_979 ? tlb_sectored_entries_5_valid_2 : tlb__GEN_204; // @[TLB.scala 239:54:freechips.rocketchip.system.DefaultRV32Config.fir@178277.8]
  assign tlb__GEN_325 = tlb__T_979 ? tlb_sectored_entries_5_valid_3 : tlb__GEN_205; // @[TLB.scala 239:54:freechips.rocketchip.system.DefaultRV32Config.fir@178277.8]
  assign tlb__GEN_332 = tlb__T_979 ? tlb_sectored_entries_6_valid_0 : tlb__GEN_224; // @[TLB.scala 239:54:freechips.rocketchip.system.DefaultRV32Config.fir@178277.8]
  assign tlb__GEN_333 = tlb__T_979 ? tlb_sectored_entries_6_valid_1 : tlb__GEN_225; // @[TLB.scala 239:54:freechips.rocketchip.system.DefaultRV32Config.fir@178277.8]
  assign tlb__GEN_334 = tlb__T_979 ? tlb_sectored_entries_6_valid_2 : tlb__GEN_226; // @[TLB.scala 239:54:freechips.rocketchip.system.DefaultRV32Config.fir@178277.8]
  assign tlb__GEN_335 = tlb__T_979 ? tlb_sectored_entries_6_valid_3 : tlb__GEN_227; // @[TLB.scala 239:54:freechips.rocketchip.system.DefaultRV32Config.fir@178277.8]
  assign tlb__GEN_342 = tlb__T_979 ? tlb_sectored_entries_7_valid_0 : tlb__GEN_246; // @[TLB.scala 239:54:freechips.rocketchip.system.DefaultRV32Config.fir@178277.8]
  assign tlb__GEN_343 = tlb__T_979 ? tlb_sectored_entries_7_valid_1 : tlb__GEN_247; // @[TLB.scala 239:54:freechips.rocketchip.system.DefaultRV32Config.fir@178277.8]
  assign tlb__GEN_344 = tlb__T_979 ? tlb_sectored_entries_7_valid_2 : tlb__GEN_248; // @[TLB.scala 239:54:freechips.rocketchip.system.DefaultRV32Config.fir@178277.8]
  assign tlb__GEN_345 = tlb__T_979 ? tlb_sectored_entries_7_valid_3 : tlb__GEN_249; // @[TLB.scala 239:54:freechips.rocketchip.system.DefaultRV32Config.fir@178277.8]
  assign tlb__GEN_354 = tlb__T_961 | tlb_special_entry_valid_0; // @[TLB.scala 237:68:freechips.rocketchip.system.DefaultRV32Config.fir@178253.6]
  assign tlb__GEN_358 = tlb__T_961 ? tlb_superpage_entries_0_valid_0 : tlb__GEN_258; // @[TLB.scala 237:68:freechips.rocketchip.system.DefaultRV32Config.fir@178253.6]
  assign tlb__GEN_362 = tlb__T_961 ? tlb_superpage_entries_1_valid_0 : tlb__GEN_262; // @[TLB.scala 237:68:freechips.rocketchip.system.DefaultRV32Config.fir@178253.6]
  assign tlb__GEN_366 = tlb__T_961 ? tlb_superpage_entries_2_valid_0 : tlb__GEN_266; // @[TLB.scala 237:68:freechips.rocketchip.system.DefaultRV32Config.fir@178253.6]
  assign tlb__GEN_370 = tlb__T_961 ? tlb_superpage_entries_3_valid_0 : tlb__GEN_270; // @[TLB.scala 237:68:freechips.rocketchip.system.DefaultRV32Config.fir@178253.6]
  assign tlb__GEN_372 = tlb__T_961 ? tlb_sectored_entries_0_valid_0 : tlb__GEN_272; // @[TLB.scala 237:68:freechips.rocketchip.system.DefaultRV32Config.fir@178253.6]
  assign tlb__GEN_373 = tlb__T_961 ? tlb_sectored_entries_0_valid_1 : tlb__GEN_273; // @[TLB.scala 237:68:freechips.rocketchip.system.DefaultRV32Config.fir@178253.6]
  assign tlb__GEN_374 = tlb__T_961 ? tlb_sectored_entries_0_valid_2 : tlb__GEN_274; // @[TLB.scala 237:68:freechips.rocketchip.system.DefaultRV32Config.fir@178253.6]
  assign tlb__GEN_375 = tlb__T_961 ? tlb_sectored_entries_0_valid_3 : tlb__GEN_275; // @[TLB.scala 237:68:freechips.rocketchip.system.DefaultRV32Config.fir@178253.6]
  assign tlb__GEN_382 = tlb__T_961 ? tlb_sectored_entries_1_valid_0 : tlb__GEN_282; // @[TLB.scala 237:68:freechips.rocketchip.system.DefaultRV32Config.fir@178253.6]
  assign tlb__GEN_383 = tlb__T_961 ? tlb_sectored_entries_1_valid_1 : tlb__GEN_283; // @[TLB.scala 237:68:freechips.rocketchip.system.DefaultRV32Config.fir@178253.6]
  assign tlb__GEN_384 = tlb__T_961 ? tlb_sectored_entries_1_valid_2 : tlb__GEN_284; // @[TLB.scala 237:68:freechips.rocketchip.system.DefaultRV32Config.fir@178253.6]
  assign tlb__GEN_385 = tlb__T_961 ? tlb_sectored_entries_1_valid_3 : tlb__GEN_285; // @[TLB.scala 237:68:freechips.rocketchip.system.DefaultRV32Config.fir@178253.6]
  assign tlb__GEN_392 = tlb__T_961 ? tlb_sectored_entries_2_valid_0 : tlb__GEN_292; // @[TLB.scala 237:68:freechips.rocketchip.system.DefaultRV32Config.fir@178253.6]
  assign tlb__GEN_393 = tlb__T_961 ? tlb_sectored_entries_2_valid_1 : tlb__GEN_293; // @[TLB.scala 237:68:freechips.rocketchip.system.DefaultRV32Config.fir@178253.6]
  assign tlb__GEN_394 = tlb__T_961 ? tlb_sectored_entries_2_valid_2 : tlb__GEN_294; // @[TLB.scala 237:68:freechips.rocketchip.system.DefaultRV32Config.fir@178253.6]
  assign tlb__GEN_395 = tlb__T_961 ? tlb_sectored_entries_2_valid_3 : tlb__GEN_295; // @[TLB.scala 237:68:freechips.rocketchip.system.DefaultRV32Config.fir@178253.6]
  assign tlb__GEN_402 = tlb__T_961 ? tlb_sectored_entries_3_valid_0 : tlb__GEN_302; // @[TLB.scala 237:68:freechips.rocketchip.system.DefaultRV32Config.fir@178253.6]
  assign tlb__GEN_403 = tlb__T_961 ? tlb_sectored_entries_3_valid_1 : tlb__GEN_303; // @[TLB.scala 237:68:freechips.rocketchip.system.DefaultRV32Config.fir@178253.6]
  assign tlb__GEN_404 = tlb__T_961 ? tlb_sectored_entries_3_valid_2 : tlb__GEN_304; // @[TLB.scala 237:68:freechips.rocketchip.system.DefaultRV32Config.fir@178253.6]
  assign tlb__GEN_405 = tlb__T_961 ? tlb_sectored_entries_3_valid_3 : tlb__GEN_305; // @[TLB.scala 237:68:freechips.rocketchip.system.DefaultRV32Config.fir@178253.6]
  assign tlb__GEN_412 = tlb__T_961 ? tlb_sectored_entries_4_valid_0 : tlb__GEN_312; // @[TLB.scala 237:68:freechips.rocketchip.system.DefaultRV32Config.fir@178253.6]
  assign tlb__GEN_413 = tlb__T_961 ? tlb_sectored_entries_4_valid_1 : tlb__GEN_313; // @[TLB.scala 237:68:freechips.rocketchip.system.DefaultRV32Config.fir@178253.6]
  assign tlb__GEN_414 = tlb__T_961 ? tlb_sectored_entries_4_valid_2 : tlb__GEN_314; // @[TLB.scala 237:68:freechips.rocketchip.system.DefaultRV32Config.fir@178253.6]
  assign tlb__GEN_415 = tlb__T_961 ? tlb_sectored_entries_4_valid_3 : tlb__GEN_315; // @[TLB.scala 237:68:freechips.rocketchip.system.DefaultRV32Config.fir@178253.6]
  assign tlb__GEN_422 = tlb__T_961 ? tlb_sectored_entries_5_valid_0 : tlb__GEN_322; // @[TLB.scala 237:68:freechips.rocketchip.system.DefaultRV32Config.fir@178253.6]
  assign tlb__GEN_423 = tlb__T_961 ? tlb_sectored_entries_5_valid_1 : tlb__GEN_323; // @[TLB.scala 237:68:freechips.rocketchip.system.DefaultRV32Config.fir@178253.6]
  assign tlb__GEN_424 = tlb__T_961 ? tlb_sectored_entries_5_valid_2 : tlb__GEN_324; // @[TLB.scala 237:68:freechips.rocketchip.system.DefaultRV32Config.fir@178253.6]
  assign tlb__GEN_425 = tlb__T_961 ? tlb_sectored_entries_5_valid_3 : tlb__GEN_325; // @[TLB.scala 237:68:freechips.rocketchip.system.DefaultRV32Config.fir@178253.6]
  assign tlb__GEN_432 = tlb__T_961 ? tlb_sectored_entries_6_valid_0 : tlb__GEN_332; // @[TLB.scala 237:68:freechips.rocketchip.system.DefaultRV32Config.fir@178253.6]
  assign tlb__GEN_433 = tlb__T_961 ? tlb_sectored_entries_6_valid_1 : tlb__GEN_333; // @[TLB.scala 237:68:freechips.rocketchip.system.DefaultRV32Config.fir@178253.6]
  assign tlb__GEN_434 = tlb__T_961 ? tlb_sectored_entries_6_valid_2 : tlb__GEN_334; // @[TLB.scala 237:68:freechips.rocketchip.system.DefaultRV32Config.fir@178253.6]
  assign tlb__GEN_435 = tlb__T_961 ? tlb_sectored_entries_6_valid_3 : tlb__GEN_335; // @[TLB.scala 237:68:freechips.rocketchip.system.DefaultRV32Config.fir@178253.6]
  assign tlb__GEN_442 = tlb__T_961 ? tlb_sectored_entries_7_valid_0 : tlb__GEN_342; // @[TLB.scala 237:68:freechips.rocketchip.system.DefaultRV32Config.fir@178253.6]
  assign tlb__GEN_443 = tlb__T_961 ? tlb_sectored_entries_7_valid_1 : tlb__GEN_343; // @[TLB.scala 237:68:freechips.rocketchip.system.DefaultRV32Config.fir@178253.6]
  assign tlb__GEN_444 = tlb__T_961 ? tlb_sectored_entries_7_valid_2 : tlb__GEN_344; // @[TLB.scala 237:68:freechips.rocketchip.system.DefaultRV32Config.fir@178253.6]
  assign tlb__GEN_445 = tlb__T_961 ? tlb_sectored_entries_7_valid_3 : tlb__GEN_345; // @[TLB.scala 237:68:freechips.rocketchip.system.DefaultRV32Config.fir@178253.6]
  assign tlb__GEN_454 = tlb__T_939 ? tlb__GEN_354 : tlb_special_entry_valid_0; // @[TLB.scala 217:42:freechips.rocketchip.system.DefaultRV32Config.fir@178212.4]
  assign tlb__GEN_458 = tlb__T_939 ? tlb__GEN_358 : tlb_superpage_entries_0_valid_0; // @[TLB.scala 217:42:freechips.rocketchip.system.DefaultRV32Config.fir@178212.4]
  assign tlb__GEN_462 = tlb__T_939 ? tlb__GEN_362 : tlb_superpage_entries_1_valid_0; // @[TLB.scala 217:42:freechips.rocketchip.system.DefaultRV32Config.fir@178212.4]
  assign tlb__GEN_466 = tlb__T_939 ? tlb__GEN_366 : tlb_superpage_entries_2_valid_0; // @[TLB.scala 217:42:freechips.rocketchip.system.DefaultRV32Config.fir@178212.4]
  assign tlb__GEN_470 = tlb__T_939 ? tlb__GEN_370 : tlb_superpage_entries_3_valid_0; // @[TLB.scala 217:42:freechips.rocketchip.system.DefaultRV32Config.fir@178212.4]
  assign tlb__GEN_472 = tlb__T_939 ? tlb__GEN_372 : tlb_sectored_entries_0_valid_0; // @[TLB.scala 217:42:freechips.rocketchip.system.DefaultRV32Config.fir@178212.4]
  assign tlb__GEN_473 = tlb__T_939 ? tlb__GEN_373 : tlb_sectored_entries_0_valid_1; // @[TLB.scala 217:42:freechips.rocketchip.system.DefaultRV32Config.fir@178212.4]
  assign tlb__GEN_474 = tlb__T_939 ? tlb__GEN_374 : tlb_sectored_entries_0_valid_2; // @[TLB.scala 217:42:freechips.rocketchip.system.DefaultRV32Config.fir@178212.4]
  assign tlb__GEN_475 = tlb__T_939 ? tlb__GEN_375 : tlb_sectored_entries_0_valid_3; // @[TLB.scala 217:42:freechips.rocketchip.system.DefaultRV32Config.fir@178212.4]
  assign tlb__GEN_482 = tlb__T_939 ? tlb__GEN_382 : tlb_sectored_entries_1_valid_0; // @[TLB.scala 217:42:freechips.rocketchip.system.DefaultRV32Config.fir@178212.4]
  assign tlb__GEN_483 = tlb__T_939 ? tlb__GEN_383 : tlb_sectored_entries_1_valid_1; // @[TLB.scala 217:42:freechips.rocketchip.system.DefaultRV32Config.fir@178212.4]
  assign tlb__GEN_484 = tlb__T_939 ? tlb__GEN_384 : tlb_sectored_entries_1_valid_2; // @[TLB.scala 217:42:freechips.rocketchip.system.DefaultRV32Config.fir@178212.4]
  assign tlb__GEN_485 = tlb__T_939 ? tlb__GEN_385 : tlb_sectored_entries_1_valid_3; // @[TLB.scala 217:42:freechips.rocketchip.system.DefaultRV32Config.fir@178212.4]
  assign tlb__GEN_492 = tlb__T_939 ? tlb__GEN_392 : tlb_sectored_entries_2_valid_0; // @[TLB.scala 217:42:freechips.rocketchip.system.DefaultRV32Config.fir@178212.4]
  assign tlb__GEN_493 = tlb__T_939 ? tlb__GEN_393 : tlb_sectored_entries_2_valid_1; // @[TLB.scala 217:42:freechips.rocketchip.system.DefaultRV32Config.fir@178212.4]
  assign tlb__GEN_494 = tlb__T_939 ? tlb__GEN_394 : tlb_sectored_entries_2_valid_2; // @[TLB.scala 217:42:freechips.rocketchip.system.DefaultRV32Config.fir@178212.4]
  assign tlb__GEN_495 = tlb__T_939 ? tlb__GEN_395 : tlb_sectored_entries_2_valid_3; // @[TLB.scala 217:42:freechips.rocketchip.system.DefaultRV32Config.fir@178212.4]
  assign tlb__GEN_502 = tlb__T_939 ? tlb__GEN_402 : tlb_sectored_entries_3_valid_0; // @[TLB.scala 217:42:freechips.rocketchip.system.DefaultRV32Config.fir@178212.4]
  assign tlb__GEN_503 = tlb__T_939 ? tlb__GEN_403 : tlb_sectored_entries_3_valid_1; // @[TLB.scala 217:42:freechips.rocketchip.system.DefaultRV32Config.fir@178212.4]
  assign tlb__GEN_504 = tlb__T_939 ? tlb__GEN_404 : tlb_sectored_entries_3_valid_2; // @[TLB.scala 217:42:freechips.rocketchip.system.DefaultRV32Config.fir@178212.4]
  assign tlb__GEN_505 = tlb__T_939 ? tlb__GEN_405 : tlb_sectored_entries_3_valid_3; // @[TLB.scala 217:42:freechips.rocketchip.system.DefaultRV32Config.fir@178212.4]
  assign tlb__GEN_512 = tlb__T_939 ? tlb__GEN_412 : tlb_sectored_entries_4_valid_0; // @[TLB.scala 217:42:freechips.rocketchip.system.DefaultRV32Config.fir@178212.4]
  assign tlb__GEN_513 = tlb__T_939 ? tlb__GEN_413 : tlb_sectored_entries_4_valid_1; // @[TLB.scala 217:42:freechips.rocketchip.system.DefaultRV32Config.fir@178212.4]
  assign tlb__GEN_514 = tlb__T_939 ? tlb__GEN_414 : tlb_sectored_entries_4_valid_2; // @[TLB.scala 217:42:freechips.rocketchip.system.DefaultRV32Config.fir@178212.4]
  assign tlb__GEN_515 = tlb__T_939 ? tlb__GEN_415 : tlb_sectored_entries_4_valid_3; // @[TLB.scala 217:42:freechips.rocketchip.system.DefaultRV32Config.fir@178212.4]
  assign tlb__GEN_522 = tlb__T_939 ? tlb__GEN_422 : tlb_sectored_entries_5_valid_0; // @[TLB.scala 217:42:freechips.rocketchip.system.DefaultRV32Config.fir@178212.4]
  assign tlb__GEN_523 = tlb__T_939 ? tlb__GEN_423 : tlb_sectored_entries_5_valid_1; // @[TLB.scala 217:42:freechips.rocketchip.system.DefaultRV32Config.fir@178212.4]
  assign tlb__GEN_524 = tlb__T_939 ? tlb__GEN_424 : tlb_sectored_entries_5_valid_2; // @[TLB.scala 217:42:freechips.rocketchip.system.DefaultRV32Config.fir@178212.4]
  assign tlb__GEN_525 = tlb__T_939 ? tlb__GEN_425 : tlb_sectored_entries_5_valid_3; // @[TLB.scala 217:42:freechips.rocketchip.system.DefaultRV32Config.fir@178212.4]
  assign tlb__GEN_532 = tlb__T_939 ? tlb__GEN_432 : tlb_sectored_entries_6_valid_0; // @[TLB.scala 217:42:freechips.rocketchip.system.DefaultRV32Config.fir@178212.4]
  assign tlb__GEN_533 = tlb__T_939 ? tlb__GEN_433 : tlb_sectored_entries_6_valid_1; // @[TLB.scala 217:42:freechips.rocketchip.system.DefaultRV32Config.fir@178212.4]
  assign tlb__GEN_534 = tlb__T_939 ? tlb__GEN_434 : tlb_sectored_entries_6_valid_2; // @[TLB.scala 217:42:freechips.rocketchip.system.DefaultRV32Config.fir@178212.4]
  assign tlb__GEN_535 = tlb__T_939 ? tlb__GEN_435 : tlb_sectored_entries_6_valid_3; // @[TLB.scala 217:42:freechips.rocketchip.system.DefaultRV32Config.fir@178212.4]
  assign tlb__GEN_542 = tlb__T_939 ? tlb__GEN_442 : tlb_sectored_entries_7_valid_0; // @[TLB.scala 217:42:freechips.rocketchip.system.DefaultRV32Config.fir@178212.4]
  assign tlb__GEN_543 = tlb__T_939 ? tlb__GEN_443 : tlb_sectored_entries_7_valid_1; // @[TLB.scala 217:42:freechips.rocketchip.system.DefaultRV32Config.fir@178212.4]
  assign tlb__GEN_544 = tlb__T_939 ? tlb__GEN_444 : tlb_sectored_entries_7_valid_2; // @[TLB.scala 217:42:freechips.rocketchip.system.DefaultRV32Config.fir@178212.4]
  assign tlb__GEN_545 = tlb__T_939 ? tlb__GEN_445 : tlb_sectored_entries_7_valid_3; // @[TLB.scala 217:42:freechips.rocketchip.system.DefaultRV32Config.fir@178212.4]
  assign tlb__T_1659 = {tlb_OptimizationBarrier_19_io_y_ae,tlb_OptimizationBarrier_18_io_y_ae,tlb_OptimizationBarrier_17_io_y_ae,tlb_OptimizationBarrier_16_io_y_ae,tlb_OptimizationBarrier_15_io_y_ae,tlb_OptimizationBarrier_14_io_y_ae}; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@179681.4]
  assign tlb_ptw_ae_array = {1'h0,tlb_OptimizationBarrier_26_io_y_ae,tlb_OptimizationBarrier_25_io_y_ae,tlb_OptimizationBarrier_24_io_y_ae,tlb_OptimizationBarrier_23_io_y_ae,tlb_OptimizationBarrier_22_io_y_ae,tlb_OptimizationBarrier_21_io_y_ae,tlb_OptimizationBarrier_20_io_y_ae,tlb__T_1659}; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@179689.4]
  assign tlb__T_1667 = ~tlb_priv_s; // @[TLB.scala 256:24:freechips.rocketchip.system.DefaultRV32Config.fir@179690.4]
  assign tlb__T_1668 = tlb__T_1667 | tlb_io_ptw_status_sum; // @[TLB.scala 256:32:freechips.rocketchip.system.DefaultRV32Config.fir@179691.4]
  assign tlb__T_1673 = {tlb_OptimizationBarrier_19_io_y_u,tlb_OptimizationBarrier_18_io_y_u,tlb_OptimizationBarrier_17_io_y_u,tlb_OptimizationBarrier_16_io_y_u,tlb_OptimizationBarrier_15_io_y_u,tlb_OptimizationBarrier_14_io_y_u}; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@179696.4]
  assign tlb__T_1680 = {tlb_OptimizationBarrier_26_io_y_u,tlb_OptimizationBarrier_25_io_y_u,tlb_OptimizationBarrier_24_io_y_u,tlb_OptimizationBarrier_23_io_y_u,tlb_OptimizationBarrier_22_io_y_u,tlb_OptimizationBarrier_21_io_y_u,tlb_OptimizationBarrier_20_io_y_u,tlb__T_1673}; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@179703.4]
  assign tlb__T_1681 = tlb__T_1668 ? tlb__T_1680 : 13'h0; // @[TLB.scala 256:23:freechips.rocketchip.system.DefaultRV32Config.fir@179704.4]
  assign tlb__T_1694 = ~tlb__T_1680; // @[TLB.scala 256:98:freechips.rocketchip.system.DefaultRV32Config.fir@179717.4]
  assign tlb__T_1695 = tlb_priv_s ? tlb__T_1694 : 13'h0; // @[TLB.scala 256:89:freechips.rocketchip.system.DefaultRV32Config.fir@179718.4]
  assign tlb_priv_rw_ok = tlb__T_1681 | tlb__T_1695; // @[TLB.scala 256:84:freechips.rocketchip.system.DefaultRV32Config.fir@179719.4]
  assign tlb__T_1725 = {tlb_OptimizationBarrier_19_io_y_sr,tlb_OptimizationBarrier_18_io_y_sr,tlb_OptimizationBarrier_17_io_y_sr,tlb_OptimizationBarrier_16_io_y_sr,tlb_OptimizationBarrier_15_io_y_sr,tlb_OptimizationBarrier_14_io_y_sr}; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@179750.4]
  assign tlb__T_1732 = {tlb_OptimizationBarrier_26_io_y_sr,tlb_OptimizationBarrier_25_io_y_sr,tlb_OptimizationBarrier_24_io_y_sr,tlb_OptimizationBarrier_23_io_y_sr,tlb_OptimizationBarrier_22_io_y_sr,tlb_OptimizationBarrier_21_io_y_sr,tlb_OptimizationBarrier_20_io_y_sr,tlb__T_1725}; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@179757.4]
  assign tlb__T_1737 = {tlb_OptimizationBarrier_19_io_y_sx,tlb_OptimizationBarrier_18_io_y_sx,tlb_OptimizationBarrier_17_io_y_sx,tlb_OptimizationBarrier_16_io_y_sx,tlb_OptimizationBarrier_15_io_y_sx,tlb_OptimizationBarrier_14_io_y_sx}; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@179762.4]
  assign tlb__T_1744 = {tlb_OptimizationBarrier_26_io_y_sx,tlb_OptimizationBarrier_25_io_y_sx,tlb_OptimizationBarrier_24_io_y_sx,tlb_OptimizationBarrier_23_io_y_sx,tlb_OptimizationBarrier_22_io_y_sx,tlb_OptimizationBarrier_21_io_y_sx,tlb_OptimizationBarrier_20_io_y_sx,tlb__T_1737}; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@179769.4]
  assign tlb__T_1745 = tlb_io_ptw_status_mxr ? tlb__T_1744 : 13'h0; // @[TLB.scala 258:73:freechips.rocketchip.system.DefaultRV32Config.fir@179770.4]
  assign tlb__T_1746 = tlb__T_1732 | tlb__T_1745; // @[TLB.scala 258:68:freechips.rocketchip.system.DefaultRV32Config.fir@179771.4]
  assign tlb__T_1747 = tlb_priv_rw_ok & tlb__T_1746; // @[TLB.scala 258:40:freechips.rocketchip.system.DefaultRV32Config.fir@179772.4]
  assign tlb_r_array = {1'h1,tlb__T_1747}; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@179773.4]
  assign tlb__T_1752 = {tlb_OptimizationBarrier_19_io_y_sw,tlb_OptimizationBarrier_18_io_y_sw,tlb_OptimizationBarrier_17_io_y_sw,tlb_OptimizationBarrier_16_io_y_sw,tlb_OptimizationBarrier_15_io_y_sw,tlb_OptimizationBarrier_14_io_y_sw}; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@179778.4]
  assign tlb__T_1759 = {tlb_OptimizationBarrier_26_io_y_sw,tlb_OptimizationBarrier_25_io_y_sw,tlb_OptimizationBarrier_24_io_y_sw,tlb_OptimizationBarrier_23_io_y_sw,tlb_OptimizationBarrier_22_io_y_sw,tlb_OptimizationBarrier_21_io_y_sw,tlb_OptimizationBarrier_20_io_y_sw,tlb__T_1752}; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@179785.4]
  assign tlb__T_1760 = tlb_priv_rw_ok & tlb__T_1759; // @[TLB.scala 259:40:freechips.rocketchip.system.DefaultRV32Config.fir@179786.4]
  assign tlb_w_array = {1'h1,tlb__T_1760}; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@179787.4]
  assign tlb__T_1775 = tlb_prot_r ? 2'h3 : 2'h0; // @[Bitwise.scala 72:12:freechips.rocketchip.system.DefaultRV32Config.fir@179803.4]
  assign tlb__T_1780 = {tlb_OptimizationBarrier_32_io_y_pr,tlb_OptimizationBarrier_31_io_y_pr,tlb_OptimizationBarrier_30_io_y_pr,tlb_OptimizationBarrier_29_io_y_pr,tlb_OptimizationBarrier_28_io_y_pr,tlb_OptimizationBarrier_27_io_y_pr}; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@179808.4]
  assign tlb__T_1787 = {tlb__T_1775,tlb_OptimizationBarrier_38_io_y_pr,tlb_OptimizationBarrier_37_io_y_pr,tlb_OptimizationBarrier_36_io_y_pr,tlb_OptimizationBarrier_35_io_y_pr,tlb_OptimizationBarrier_34_io_y_pr,tlb_OptimizationBarrier_33_io_y_pr,tlb__T_1780}; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@179815.4]
  assign tlb__T_1788 = ~tlb_ptw_ae_array; // @[TLB.scala 261:89:freechips.rocketchip.system.DefaultRV32Config.fir@179816.4]
  assign tlb_pr_array = tlb__T_1787 & tlb__T_1788; // @[TLB.scala 261:87:freechips.rocketchip.system.DefaultRV32Config.fir@179817.4]
  assign tlb__T_1790 = tlb_prot_w ? 2'h3 : 2'h0; // @[Bitwise.scala 72:12:freechips.rocketchip.system.DefaultRV32Config.fir@179819.4]
  assign tlb__T_1795 = {tlb_OptimizationBarrier_32_io_y_pw,tlb_OptimizationBarrier_31_io_y_pw,tlb_OptimizationBarrier_30_io_y_pw,tlb_OptimizationBarrier_29_io_y_pw,tlb_OptimizationBarrier_28_io_y_pw,tlb_OptimizationBarrier_27_io_y_pw}; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@179824.4]
  assign tlb__T_1802 = {tlb__T_1790,tlb_OptimizationBarrier_38_io_y_pw,tlb_OptimizationBarrier_37_io_y_pw,tlb_OptimizationBarrier_36_io_y_pw,tlb_OptimizationBarrier_35_io_y_pw,tlb_OptimizationBarrier_34_io_y_pw,tlb_OptimizationBarrier_33_io_y_pw,tlb__T_1795}; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@179831.4]
  assign tlb_pw_array = tlb__T_1802 & tlb__T_1788; // @[TLB.scala 262:87:freechips.rocketchip.system.DefaultRV32Config.fir@179833.4]
  assign tlb__T_1820 = tlb_prot_eff ? 2'h3 : 2'h0; // @[Bitwise.scala 72:12:freechips.rocketchip.system.DefaultRV32Config.fir@179851.4]
  assign tlb__T_1825 = {tlb_OptimizationBarrier_32_io_y_eff,tlb_OptimizationBarrier_31_io_y_eff,tlb_OptimizationBarrier_30_io_y_eff,tlb_OptimizationBarrier_29_io_y_eff,tlb_OptimizationBarrier_28_io_y_eff,tlb_OptimizationBarrier_27_io_y_eff}; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@179856.4]
  assign tlb_eff_array = {tlb__T_1820,tlb_OptimizationBarrier_38_io_y_eff,tlb_OptimizationBarrier_37_io_y_eff,tlb_OptimizationBarrier_36_io_y_eff,tlb_OptimizationBarrier_35_io_y_eff,tlb_OptimizationBarrier_34_io_y_eff,tlb_OptimizationBarrier_33_io_y_eff,tlb__T_1825}; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@179863.4]
  assign tlb__T_1833 = tlb__T_93 ? 2'h3 : 2'h0; // @[Bitwise.scala 72:12:freechips.rocketchip.system.DefaultRV32Config.fir@179865.4]
  assign tlb__T_1838 = {tlb_OptimizationBarrier_32_io_y_c,tlb_OptimizationBarrier_31_io_y_c,tlb_OptimizationBarrier_30_io_y_c,tlb_OptimizationBarrier_29_io_y_c,tlb_OptimizationBarrier_28_io_y_c,tlb_OptimizationBarrier_27_io_y_c}; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@179870.4]
  assign tlb_c_array = {tlb__T_1833,tlb_OptimizationBarrier_38_io_y_c,tlb_OptimizationBarrier_37_io_y_c,tlb_OptimizationBarrier_36_io_y_c,tlb_OptimizationBarrier_35_io_y_c,tlb_OptimizationBarrier_34_io_y_c,tlb_OptimizationBarrier_33_io_y_c,tlb__T_1838}; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@179877.4]
  assign tlb__T_1846 = tlb__T_232 ? 2'h3 : 2'h0; // @[Bitwise.scala 72:12:freechips.rocketchip.system.DefaultRV32Config.fir@179879.4]
  assign tlb__T_1851 = {tlb_OptimizationBarrier_32_io_y_ppp,tlb_OptimizationBarrier_31_io_y_ppp,tlb_OptimizationBarrier_30_io_y_ppp,tlb_OptimizationBarrier_29_io_y_ppp,tlb_OptimizationBarrier_28_io_y_ppp,tlb_OptimizationBarrier_27_io_y_ppp}; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@179884.4]
  assign tlb_ppp_array = {tlb__T_1846,tlb_OptimizationBarrier_38_io_y_ppp,tlb_OptimizationBarrier_37_io_y_ppp,tlb_OptimizationBarrier_36_io_y_ppp,tlb_OptimizationBarrier_35_io_y_ppp,tlb_OptimizationBarrier_34_io_y_ppp,tlb_OptimizationBarrier_33_io_y_ppp,tlb__T_1851}; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@179891.4]
  assign tlb__T_1859 = tlb_prot_al ? 2'h3 : 2'h0; // @[Bitwise.scala 72:12:freechips.rocketchip.system.DefaultRV32Config.fir@179893.4]
  assign tlb__T_1864 = {tlb_OptimizationBarrier_32_io_y_paa,tlb_OptimizationBarrier_31_io_y_paa,tlb_OptimizationBarrier_30_io_y_paa,tlb_OptimizationBarrier_29_io_y_paa,tlb_OptimizationBarrier_28_io_y_paa,tlb_OptimizationBarrier_27_io_y_paa}; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@179898.4]
  assign tlb_paa_array = {tlb__T_1859,tlb_OptimizationBarrier_38_io_y_paa,tlb_OptimizationBarrier_37_io_y_paa,tlb_OptimizationBarrier_36_io_y_paa,tlb_OptimizationBarrier_35_io_y_paa,tlb_OptimizationBarrier_34_io_y_paa,tlb_OptimizationBarrier_33_io_y_paa,tlb__T_1864}; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@179905.4]
  assign tlb__T_1877 = {tlb_OptimizationBarrier_32_io_y_pal,tlb_OptimizationBarrier_31_io_y_pal,tlb_OptimizationBarrier_30_io_y_pal,tlb_OptimizationBarrier_29_io_y_pal,tlb_OptimizationBarrier_28_io_y_pal,tlb_OptimizationBarrier_27_io_y_pal}; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@179912.4]
  assign tlb_pal_array = {tlb__T_1859,tlb_OptimizationBarrier_38_io_y_pal,tlb_OptimizationBarrier_37_io_y_pal,tlb_OptimizationBarrier_36_io_y_pal,tlb_OptimizationBarrier_35_io_y_pal,tlb_OptimizationBarrier_34_io_y_pal,tlb_OptimizationBarrier_33_io_y_pal,tlb__T_1877}; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@179919.4]
  assign tlb_ppp_array_if_cached = tlb_ppp_array | tlb_c_array; // @[TLB.scala 269:39:freechips.rocketchip.system.DefaultRV32Config.fir@179920.4]
  assign tlb_paa_array_if_cached = tlb_paa_array | tlb_c_array; // @[TLB.scala 270:39:freechips.rocketchip.system.DefaultRV32Config.fir@179922.4]
  assign tlb_pal_array_if_cached = tlb_pal_array | tlb_c_array; // @[TLB.scala 271:39:freechips.rocketchip.system.DefaultRV32Config.fir@179924.4]
  assign tlb__T_1899 = 4'h1 << tlb_io_req_bits_size; // @[OneHot.scala 58:35:freechips.rocketchip.system.DefaultRV32Config.fir@179939.4]
  assign tlb__T_1901 = tlb__T_1899 - 4'h1; // @[TLB.scala 274:69:freechips.rocketchip.system.DefaultRV32Config.fir@179941.4]
  assign _GEN_375 = {{28'd0}, tlb__T_1901}; // @[TLB.scala 274:39:freechips.rocketchip.system.DefaultRV32Config.fir@179942.4]
  assign tlb__T_1902 = tlb_io_req_bits_vaddr & _GEN_375; // @[TLB.scala 274:39:freechips.rocketchip.system.DefaultRV32Config.fir@179942.4]
  assign tlb_misaligned = |tlb__T_1902; // @[TLB.scala 274:75:freechips.rocketchip.system.DefaultRV32Config.fir@179943.4]
  assign tlb__T_1903 = tlb_io_req_bits_cmd == 5'h6; // @[package.scala 15:47:freechips.rocketchip.system.DefaultRV32Config.fir@179944.4]
  assign tlb__T_1904 = tlb_io_req_bits_cmd == 5'h7; // @[package.scala 15:47:freechips.rocketchip.system.DefaultRV32Config.fir@179945.4]
  assign tlb__T_1905 = tlb__T_1903 | tlb__T_1904; // @[package.scala 64:59:freechips.rocketchip.system.DefaultRV32Config.fir@179946.4]
  assign tlb__T_1906 = tlb_io_req_bits_cmd == 5'h4; // @[package.scala 15:47:freechips.rocketchip.system.DefaultRV32Config.fir@179948.4]
  assign tlb__T_1907 = tlb_io_req_bits_cmd == 5'h9; // @[package.scala 15:47:freechips.rocketchip.system.DefaultRV32Config.fir@179949.4]
  assign tlb__T_1908 = tlb_io_req_bits_cmd == 5'ha; // @[package.scala 15:47:freechips.rocketchip.system.DefaultRV32Config.fir@179950.4]
  assign tlb__T_1909 = tlb_io_req_bits_cmd == 5'hb; // @[package.scala 15:47:freechips.rocketchip.system.DefaultRV32Config.fir@179951.4]
  assign tlb__T_1910 = tlb__T_1906 | tlb__T_1907; // @[package.scala 64:59:freechips.rocketchip.system.DefaultRV32Config.fir@179952.4]
  assign tlb__T_1911 = tlb__T_1910 | tlb__T_1908; // @[package.scala 64:59:freechips.rocketchip.system.DefaultRV32Config.fir@179953.4]
  assign tlb__T_1912 = tlb__T_1911 | tlb__T_1909; // @[package.scala 64:59:freechips.rocketchip.system.DefaultRV32Config.fir@179954.4]
  assign tlb__T_1913 = tlb_io_req_bits_cmd == 5'h8; // @[package.scala 15:47:freechips.rocketchip.system.DefaultRV32Config.fir@179956.4]
  assign tlb__T_1914 = tlb_io_req_bits_cmd == 5'hc; // @[package.scala 15:47:freechips.rocketchip.system.DefaultRV32Config.fir@179957.4]
  assign tlb__T_1915 = tlb_io_req_bits_cmd == 5'hd; // @[package.scala 15:47:freechips.rocketchip.system.DefaultRV32Config.fir@179958.4]
  assign tlb__T_1916 = tlb_io_req_bits_cmd == 5'he; // @[package.scala 15:47:freechips.rocketchip.system.DefaultRV32Config.fir@179959.4]
  assign tlb__T_1917 = tlb_io_req_bits_cmd == 5'hf; // @[package.scala 15:47:freechips.rocketchip.system.DefaultRV32Config.fir@179960.4]
  assign tlb__T_1918 = tlb__T_1913 | tlb__T_1914; // @[package.scala 64:59:freechips.rocketchip.system.DefaultRV32Config.fir@179961.4]
  assign tlb__T_1919 = tlb__T_1918 | tlb__T_1915; // @[package.scala 64:59:freechips.rocketchip.system.DefaultRV32Config.fir@179962.4]
  assign tlb__T_1920 = tlb__T_1919 | tlb__T_1916; // @[package.scala 64:59:freechips.rocketchip.system.DefaultRV32Config.fir@179963.4]
  assign tlb__T_1921 = tlb__T_1920 | tlb__T_1917; // @[package.scala 64:59:freechips.rocketchip.system.DefaultRV32Config.fir@179964.4]
  assign tlb_cmd_put_partial = tlb_io_req_bits_cmd == 5'h11; // @[TLB.scala 288:41:freechips.rocketchip.system.DefaultRV32Config.fir@179966.4]
  assign tlb__T_1922 = tlb_io_req_bits_cmd == 5'h0; // @[Consts.scala 82:31:freechips.rocketchip.system.DefaultRV32Config.fir@179967.4]
  assign tlb__T_1924 = tlb__T_1922 | tlb__T_1903; // @[Consts.scala 82:41:freechips.rocketchip.system.DefaultRV32Config.fir@179969.4]
  assign tlb__T_1926 = tlb__T_1924 | tlb__T_1904; // @[Consts.scala 82:58:freechips.rocketchip.system.DefaultRV32Config.fir@179971.4]
  assign tlb__T_1943 = tlb__T_1912 | tlb__T_1921; // @[Consts.scala 80:44:freechips.rocketchip.system.DefaultRV32Config.fir@179988.4]
  assign tlb_cmd_read = tlb__T_1926 | tlb__T_1943; // @[Consts.scala 82:75:freechips.rocketchip.system.DefaultRV32Config.fir@179989.4]
  assign tlb__T_1944 = tlb_io_req_bits_cmd == 5'h1; // @[Consts.scala 83:32:freechips.rocketchip.system.DefaultRV32Config.fir@179990.4]
  assign tlb__T_1946 = tlb__T_1944 | tlb_cmd_put_partial; // @[Consts.scala 83:42:freechips.rocketchip.system.DefaultRV32Config.fir@179992.4]
  assign tlb__T_1948 = tlb__T_1946 | tlb__T_1904; // @[Consts.scala 83:59:freechips.rocketchip.system.DefaultRV32Config.fir@179994.4]
  assign tlb_cmd_write = tlb__T_1948 | tlb__T_1943; // @[Consts.scala 83:76:freechips.rocketchip.system.DefaultRV32Config.fir@180012.4]
  assign tlb__T_1966 = tlb_io_req_bits_cmd == 5'h5; // @[package.scala 15:47:freechips.rocketchip.system.DefaultRV32Config.fir@180013.4]
  assign tlb__T_1967 = tlb_io_req_bits_cmd == 5'h17; // @[package.scala 15:47:freechips.rocketchip.system.DefaultRV32Config.fir@180014.4]
  assign tlb__T_1968 = tlb__T_1966 | tlb__T_1967; // @[package.scala 64:59:freechips.rocketchip.system.DefaultRV32Config.fir@180015.4]
  assign tlb_cmd_write_perms = tlb_cmd_write | tlb__T_1968; // @[TLB.scala 291:35:freechips.rocketchip.system.DefaultRV32Config.fir@180016.4]
  assign tlb__T_1969 = tlb_misaligned ? tlb_eff_array : 14'h0; // @[TLB.scala 296:8:freechips.rocketchip.system.DefaultRV32Config.fir@180018.4]
  assign tlb__T_1970 = ~tlb_c_array; // @[TLB.scala 297:19:freechips.rocketchip.system.DefaultRV32Config.fir@180019.4]
  assign tlb__T_1971 = tlb__T_1905 ? tlb__T_1970 : 14'h0; // @[TLB.scala 297:8:freechips.rocketchip.system.DefaultRV32Config.fir@180020.4]
  assign tlb_ae_array = tlb__T_1969 | tlb__T_1971; // @[TLB.scala 296:37:freechips.rocketchip.system.DefaultRV32Config.fir@180021.4]
  assign tlb__T_1972 = ~tlb_pr_array; // @[TLB.scala 298:46:freechips.rocketchip.system.DefaultRV32Config.fir@180022.4]
  assign tlb__T_1973 = tlb_ae_array | tlb__T_1972; // @[TLB.scala 298:44:freechips.rocketchip.system.DefaultRV32Config.fir@180023.4]
  assign tlb_ae_ld_array = tlb_cmd_read ? tlb__T_1973 : 14'h0; // @[TLB.scala 298:24:freechips.rocketchip.system.DefaultRV32Config.fir@180024.4]
  assign tlb__T_1974 = ~tlb_pw_array; // @[TLB.scala 300:37:freechips.rocketchip.system.DefaultRV32Config.fir@180025.4]
  assign tlb__T_1975 = tlb_ae_array | tlb__T_1974; // @[TLB.scala 300:35:freechips.rocketchip.system.DefaultRV32Config.fir@180026.4]
  assign tlb__T_1976 = tlb_cmd_write_perms ? tlb__T_1975 : 14'h0; // @[TLB.scala 300:8:freechips.rocketchip.system.DefaultRV32Config.fir@180027.4]
  assign tlb__T_1977 = ~tlb_ppp_array_if_cached; // @[TLB.scala 301:26:freechips.rocketchip.system.DefaultRV32Config.fir@180028.4]
  assign tlb__T_1978 = tlb_cmd_put_partial ? tlb__T_1977 : 14'h0; // @[TLB.scala 301:8:freechips.rocketchip.system.DefaultRV32Config.fir@180029.4]
  assign tlb__T_1979 = tlb__T_1976 | tlb__T_1978; // @[TLB.scala 300:53:freechips.rocketchip.system.DefaultRV32Config.fir@180030.4]
  assign tlb__T_1980 = ~tlb_pal_array_if_cached; // @[TLB.scala 302:26:freechips.rocketchip.system.DefaultRV32Config.fir@180031.4]
  assign tlb__T_1981 = tlb__T_1912 ? tlb__T_1980 : 14'h0; // @[TLB.scala 302:8:freechips.rocketchip.system.DefaultRV32Config.fir@180032.4]
  assign tlb__T_1982 = tlb__T_1979 | tlb__T_1981; // @[TLB.scala 301:53:freechips.rocketchip.system.DefaultRV32Config.fir@180033.4]
  assign tlb__T_1983 = ~tlb_paa_array_if_cached; // @[TLB.scala 303:29:freechips.rocketchip.system.DefaultRV32Config.fir@180034.4]
  assign tlb__T_1984 = tlb__T_1921 ? tlb__T_1983 : 14'h0; // @[TLB.scala 303:8:freechips.rocketchip.system.DefaultRV32Config.fir@180035.4]
  assign tlb_ae_st_array = tlb__T_1982 | tlb__T_1984; // @[TLB.scala 302:53:freechips.rocketchip.system.DefaultRV32Config.fir@180036.4]
  assign tlb__T_1995 = tlb_misaligned & tlb_cmd_read; // @[TLB.scala 309:36:freechips.rocketchip.system.DefaultRV32Config.fir@180048.4]
  assign tlb__T_1996 = ~tlb_eff_array; // @[TLB.scala 309:49:freechips.rocketchip.system.DefaultRV32Config.fir@180049.4]
  assign tlb_ma_ld_array = tlb__T_1995 ? tlb__T_1996 : 14'h0; // @[TLB.scala 309:24:freechips.rocketchip.system.DefaultRV32Config.fir@180050.4]
  assign tlb__T_1997 = tlb_misaligned & tlb_cmd_write; // @[TLB.scala 310:36:freechips.rocketchip.system.DefaultRV32Config.fir@180051.4]
  assign tlb_ma_st_array = tlb__T_1997 ? tlb__T_1996 : 14'h0; // @[TLB.scala 310:24:freechips.rocketchip.system.DefaultRV32Config.fir@180053.4]
  assign tlb__T_1999 = tlb_r_array | tlb_ptw_ae_array; // @[TLB.scala 311:45:freechips.rocketchip.system.DefaultRV32Config.fir@180054.4]
  assign tlb__T_2000 = ~tlb__T_1999; // @[TLB.scala 311:35:freechips.rocketchip.system.DefaultRV32Config.fir@180055.4]
  assign tlb_pf_ld_array = tlb_cmd_read ? tlb__T_2000 : 14'h0; // @[TLB.scala 311:24:freechips.rocketchip.system.DefaultRV32Config.fir@180056.4]
  assign tlb__T_2001 = tlb_w_array | tlb_ptw_ae_array; // @[TLB.scala 312:52:freechips.rocketchip.system.DefaultRV32Config.fir@180057.4]
  assign tlb__T_2002 = ~tlb__T_2001; // @[TLB.scala 312:42:freechips.rocketchip.system.DefaultRV32Config.fir@180058.4]
  assign tlb_pf_st_array = tlb_cmd_write_perms ? tlb__T_2002 : 14'h0; // @[TLB.scala 312:24:freechips.rocketchip.system.DefaultRV32Config.fir@180059.4]
  assign tlb_tlb_hit = |tlb_real_hits; // @[TLB.scala 315:27:freechips.rocketchip.system.DefaultRV32Config.fir@180062.4]
  assign tlb__T_2006 = ~tlb_tlb_hit; // @[TLB.scala 316:43:freechips.rocketchip.system.DefaultRV32Config.fir@180065.4]
  assign tlb_tlb_miss = tlb_vm_enabled & tlb__T_2006; // @[TLB.scala 316:40:freechips.rocketchip.system.DefaultRV32Config.fir@180066.4]
  assign tlb__T_2009 = tlb_io_req_valid & tlb_vm_enabled; // @[TLB.scala 320:22:freechips.rocketchip.system.DefaultRV32Config.fir@180069.4]
  assign tlb__T_2010 = tlb_sector_hits_0 | tlb_sector_hits_1; // @[package.scala 64:59:freechips.rocketchip.system.DefaultRV32Config.fir@180071.6]
  assign tlb__T_2011 = tlb__T_2010 | tlb_sector_hits_2; // @[package.scala 64:59:freechips.rocketchip.system.DefaultRV32Config.fir@180072.6]
  assign tlb__T_2012 = tlb__T_2011 | tlb_sector_hits_3; // @[package.scala 64:59:freechips.rocketchip.system.DefaultRV32Config.fir@180073.6]
  assign tlb__T_2013 = tlb__T_2012 | tlb_sector_hits_4; // @[package.scala 64:59:freechips.rocketchip.system.DefaultRV32Config.fir@180074.6]
  assign tlb__T_2014 = tlb__T_2013 | tlb_sector_hits_5; // @[package.scala 64:59:freechips.rocketchip.system.DefaultRV32Config.fir@180075.6]
  assign tlb__T_2015 = tlb__T_2014 | tlb_sector_hits_6; // @[package.scala 64:59:freechips.rocketchip.system.DefaultRV32Config.fir@180076.6]
  assign tlb__T_2016 = tlb__T_2015 | tlb_sector_hits_7; // @[package.scala 64:59:freechips.rocketchip.system.DefaultRV32Config.fir@180077.6]
  assign tlb__T_2023 = {tlb_sector_hits_7,tlb_sector_hits_6,tlb_sector_hits_5,tlb_sector_hits_4,tlb_sector_hits_3,tlb_sector_hits_2,tlb_sector_hits_1,tlb_sector_hits_0}; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@180085.8]
  assign tlb__T_2024 = tlb__T_2023[7:4]; // @[OneHot.scala 30:18:freechips.rocketchip.system.DefaultRV32Config.fir@180086.8]
  assign tlb__T_2025 = tlb__T_2023[3:0]; // @[OneHot.scala 31:18:freechips.rocketchip.system.DefaultRV32Config.fir@180087.8]
  assign tlb__T_2026 = |tlb__T_2024; // @[OneHot.scala 32:14:freechips.rocketchip.system.DefaultRV32Config.fir@180088.8]
  assign tlb__T_2027 = tlb__T_2024 | tlb__T_2025; // @[OneHot.scala 32:28:freechips.rocketchip.system.DefaultRV32Config.fir@180089.8]
  assign tlb__T_2028 = tlb__T_2027[3:2]; // @[OneHot.scala 30:18:freechips.rocketchip.system.DefaultRV32Config.fir@180090.8]
  assign tlb__T_2029 = tlb__T_2027[1:0]; // @[OneHot.scala 31:18:freechips.rocketchip.system.DefaultRV32Config.fir@180091.8]
  assign tlb__T_2030 = |tlb__T_2028; // @[OneHot.scala 32:14:freechips.rocketchip.system.DefaultRV32Config.fir@180092.8]
  assign tlb__T_2031 = tlb__T_2028 | tlb__T_2029; // @[OneHot.scala 32:28:freechips.rocketchip.system.DefaultRV32Config.fir@180093.8]
  assign tlb__T_2032 = tlb__T_2031[1]; // @[CircuitMath.scala 30:8:freechips.rocketchip.system.DefaultRV32Config.fir@180094.8]
  assign tlb__T_2034 = {tlb__T_2026,tlb__T_2030,tlb__T_2032}; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@180096.8]
  assign tlb__T_2036 = tlb__T_2034[2]; // @[Replacement.scala 186:43:freechips.rocketchip.system.DefaultRV32Config.fir@180098.8]
  assign tlb__T_2037 = ~tlb__T_2036; // @[Replacement.scala 186:33:freechips.rocketchip.system.DefaultRV32Config.fir@180099.8]
  assign tlb__T_2038 = tlb__T_2007[5:3]; // @[package.scala 138:13:freechips.rocketchip.system.DefaultRV32Config.fir@180100.8]
  assign tlb__T_2039 = tlb__T_2007[2:0]; // @[Replacement.scala 188:38:freechips.rocketchip.system.DefaultRV32Config.fir@180101.8]
  assign tlb__T_2040 = tlb__T_2034[1:0]; // @[package.scala 138:13:freechips.rocketchip.system.DefaultRV32Config.fir@180102.8]
  assign tlb__T_2041 = tlb__T_2040[1]; // @[Replacement.scala 186:43:freechips.rocketchip.system.DefaultRV32Config.fir@180103.8]
  assign tlb__T_2042 = ~tlb__T_2041; // @[Replacement.scala 186:33:freechips.rocketchip.system.DefaultRV32Config.fir@180104.8]
  assign tlb__T_2043 = tlb__T_2038[1]; // @[package.scala 138:13:freechips.rocketchip.system.DefaultRV32Config.fir@180105.8]
  assign tlb__T_2044 = tlb__T_2038[0]; // @[Replacement.scala 188:38:freechips.rocketchip.system.DefaultRV32Config.fir@180106.8]
  assign tlb__T_2045 = tlb__T_2040[0]; // @[package.scala 138:13:freechips.rocketchip.system.DefaultRV32Config.fir@180107.8]
  assign tlb__T_2047 = ~tlb__T_2045; // @[Replacement.scala 208:7:freechips.rocketchip.system.DefaultRV32Config.fir@180109.8]
  assign tlb__T_2048 = tlb__T_2042 ? tlb__T_2043 : tlb__T_2047; // @[Replacement.scala 193:16:freechips.rocketchip.system.DefaultRV32Config.fir@180110.8]
  assign tlb__T_2052 = tlb__T_2042 ? tlb__T_2047 : tlb__T_2044; // @[Replacement.scala 196:16:freechips.rocketchip.system.DefaultRV32Config.fir@180114.8]
  assign tlb__T_2054 = {tlb__T_2042,tlb__T_2048,tlb__T_2052}; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@180116.8]
  assign tlb__T_2055 = tlb__T_2037 ? tlb__T_2038 : tlb__T_2054; // @[Replacement.scala 193:16:freechips.rocketchip.system.DefaultRV32Config.fir@180117.8]
  assign tlb__T_2059 = tlb__T_2039[1]; // @[package.scala 138:13:freechips.rocketchip.system.DefaultRV32Config.fir@180121.8]
  assign tlb__T_2060 = tlb__T_2039[0]; // @[Replacement.scala 188:38:freechips.rocketchip.system.DefaultRV32Config.fir@180122.8]
  assign tlb__T_2064 = tlb__T_2042 ? tlb__T_2059 : tlb__T_2047; // @[Replacement.scala 193:16:freechips.rocketchip.system.DefaultRV32Config.fir@180126.8]
  assign tlb__T_2068 = tlb__T_2042 ? tlb__T_2047 : tlb__T_2060; // @[Replacement.scala 196:16:freechips.rocketchip.system.DefaultRV32Config.fir@180130.8]
  assign tlb__T_2070 = {tlb__T_2042,tlb__T_2064,tlb__T_2068}; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@180132.8]
  assign tlb__T_2071 = tlb__T_2037 ? tlb__T_2070 : tlb__T_2039; // @[Replacement.scala 196:16:freechips.rocketchip.system.DefaultRV32Config.fir@180133.8]
  assign tlb__T_2073 = {tlb__T_2037,tlb__T_2055,tlb__T_2071}; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@180135.8]
  assign tlb__T_2074 = tlb__T_464 | tlb__T_477; // @[package.scala 64:59:freechips.rocketchip.system.DefaultRV32Config.fir@180138.6]
  assign tlb__T_2075 = tlb__T_2074 | tlb__T_490; // @[package.scala 64:59:freechips.rocketchip.system.DefaultRV32Config.fir@180139.6]
  assign tlb__T_2076 = tlb__T_2075 | tlb__T_503; // @[package.scala 64:59:freechips.rocketchip.system.DefaultRV32Config.fir@180140.6]
  assign tlb__T_2079 = {tlb__T_503,tlb__T_490,tlb__T_477,tlb__T_464}; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@180144.8]
  assign tlb__T_2080 = tlb__T_2079[3:2]; // @[OneHot.scala 30:18:freechips.rocketchip.system.DefaultRV32Config.fir@180145.8]
  assign tlb__T_2081 = tlb__T_2079[1:0]; // @[OneHot.scala 31:18:freechips.rocketchip.system.DefaultRV32Config.fir@180146.8]
  assign tlb__T_2082 = |tlb__T_2080; // @[OneHot.scala 32:14:freechips.rocketchip.system.DefaultRV32Config.fir@180147.8]
  assign tlb__T_2083 = tlb__T_2080 | tlb__T_2081; // @[OneHot.scala 32:28:freechips.rocketchip.system.DefaultRV32Config.fir@180148.8]
  assign tlb__T_2084 = tlb__T_2083[1]; // @[CircuitMath.scala 30:8:freechips.rocketchip.system.DefaultRV32Config.fir@180149.8]
  assign tlb__T_2085 = {tlb__T_2082,tlb__T_2084}; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@180150.8]
  assign tlb__T_2087 = tlb__T_2085[1]; // @[Replacement.scala 186:43:freechips.rocketchip.system.DefaultRV32Config.fir@180152.8]
  assign tlb__T_2088 = ~tlb__T_2087; // @[Replacement.scala 186:33:freechips.rocketchip.system.DefaultRV32Config.fir@180153.8]
  assign tlb__T_2089 = tlb__T_2008[1]; // @[package.scala 138:13:freechips.rocketchip.system.DefaultRV32Config.fir@180154.8]
  assign tlb__T_2090 = tlb__T_2008[0]; // @[Replacement.scala 188:38:freechips.rocketchip.system.DefaultRV32Config.fir@180155.8]
  assign tlb__T_2091 = tlb__T_2085[0]; // @[package.scala 138:13:freechips.rocketchip.system.DefaultRV32Config.fir@180156.8]
  assign tlb__T_2093 = ~tlb__T_2091; // @[Replacement.scala 208:7:freechips.rocketchip.system.DefaultRV32Config.fir@180158.8]
  assign tlb__T_2094 = tlb__T_2088 ? tlb__T_2089 : tlb__T_2093; // @[Replacement.scala 193:16:freechips.rocketchip.system.DefaultRV32Config.fir@180159.8]
  assign tlb__T_2098 = tlb__T_2088 ? tlb__T_2093 : tlb__T_2090; // @[Replacement.scala 196:16:freechips.rocketchip.system.DefaultRV32Config.fir@180163.8]
  assign tlb__T_2100 = {tlb__T_2088,tlb__T_2094,tlb__T_2098}; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@180165.8]
  assign tlb__T_2101 = tlb_real_hits[5:0]; // @[Misc.scala 180:37:freechips.rocketchip.system.DefaultRV32Config.fir@180169.4]
  assign tlb__T_2102 = tlb__T_2101[2:0]; // @[Misc.scala 180:37:freechips.rocketchip.system.DefaultRV32Config.fir@180170.4]
  assign tlb__T_2103 = tlb__T_2102[0]; // @[Misc.scala 180:37:freechips.rocketchip.system.DefaultRV32Config.fir@180171.4]
  assign tlb__T_2105 = tlb__T_2102[2:1]; // @[Misc.scala 181:39:freechips.rocketchip.system.DefaultRV32Config.fir@180173.4]
  assign tlb__T_2106 = tlb__T_2105[0]; // @[Misc.scala 180:37:freechips.rocketchip.system.DefaultRV32Config.fir@180174.4]
  assign tlb__T_2108 = tlb__T_2105[1]; // @[Misc.scala 181:39:freechips.rocketchip.system.DefaultRV32Config.fir@180176.4]
  assign tlb__T_2110 = tlb__T_2106 | tlb__T_2108; // @[Misc.scala 182:16:freechips.rocketchip.system.DefaultRV32Config.fir@180178.4]
  assign tlb__T_2112 = tlb__T_2106 & tlb__T_2108; // @[Misc.scala 182:61:freechips.rocketchip.system.DefaultRV32Config.fir@180180.4]
  assign tlb__T_2114 = tlb__T_2103 | tlb__T_2110; // @[Misc.scala 182:16:freechips.rocketchip.system.DefaultRV32Config.fir@180182.4]
  assign tlb__T_2116 = tlb__T_2103 & tlb__T_2110; // @[Misc.scala 182:61:freechips.rocketchip.system.DefaultRV32Config.fir@180184.4]
  assign tlb__T_2117 = tlb__T_2112 | tlb__T_2116; // @[Misc.scala 182:49:freechips.rocketchip.system.DefaultRV32Config.fir@180185.4]
  assign tlb__T_2118 = tlb__T_2101[5:3]; // @[Misc.scala 181:39:freechips.rocketchip.system.DefaultRV32Config.fir@180186.4]
  assign tlb__T_2119 = tlb__T_2118[0]; // @[Misc.scala 180:37:freechips.rocketchip.system.DefaultRV32Config.fir@180187.4]
  assign tlb__T_2121 = tlb__T_2118[2:1]; // @[Misc.scala 181:39:freechips.rocketchip.system.DefaultRV32Config.fir@180189.4]
  assign tlb__T_2122 = tlb__T_2121[0]; // @[Misc.scala 180:37:freechips.rocketchip.system.DefaultRV32Config.fir@180190.4]
  assign tlb__T_2124 = tlb__T_2121[1]; // @[Misc.scala 181:39:freechips.rocketchip.system.DefaultRV32Config.fir@180192.4]
  assign tlb__T_2126 = tlb__T_2122 | tlb__T_2124; // @[Misc.scala 182:16:freechips.rocketchip.system.DefaultRV32Config.fir@180194.4]
  assign tlb__T_2128 = tlb__T_2122 & tlb__T_2124; // @[Misc.scala 182:61:freechips.rocketchip.system.DefaultRV32Config.fir@180196.4]
  assign tlb__T_2130 = tlb__T_2119 | tlb__T_2126; // @[Misc.scala 182:16:freechips.rocketchip.system.DefaultRV32Config.fir@180198.4]
  assign tlb__T_2132 = tlb__T_2119 & tlb__T_2126; // @[Misc.scala 182:61:freechips.rocketchip.system.DefaultRV32Config.fir@180200.4]
  assign tlb__T_2133 = tlb__T_2128 | tlb__T_2132; // @[Misc.scala 182:49:freechips.rocketchip.system.DefaultRV32Config.fir@180201.4]
  assign tlb__T_2134 = tlb__T_2114 | tlb__T_2130; // @[Misc.scala 182:16:freechips.rocketchip.system.DefaultRV32Config.fir@180202.4]
  assign tlb__T_2135 = tlb__T_2117 | tlb__T_2133; // @[Misc.scala 182:37:freechips.rocketchip.system.DefaultRV32Config.fir@180203.4]
  assign tlb__T_2136 = tlb__T_2114 & tlb__T_2130; // @[Misc.scala 182:61:freechips.rocketchip.system.DefaultRV32Config.fir@180204.4]
  assign tlb__T_2137 = tlb__T_2135 | tlb__T_2136; // @[Misc.scala 182:49:freechips.rocketchip.system.DefaultRV32Config.fir@180205.4]
  assign tlb__T_2138 = tlb_real_hits[12:6]; // @[Misc.scala 181:39:freechips.rocketchip.system.DefaultRV32Config.fir@180206.4]
  assign tlb__T_2139 = tlb__T_2138[2:0]; // @[Misc.scala 180:37:freechips.rocketchip.system.DefaultRV32Config.fir@180207.4]
  assign tlb__T_2140 = tlb__T_2139[0]; // @[Misc.scala 180:37:freechips.rocketchip.system.DefaultRV32Config.fir@180208.4]
  assign tlb__T_2142 = tlb__T_2139[2:1]; // @[Misc.scala 181:39:freechips.rocketchip.system.DefaultRV32Config.fir@180210.4]
  assign tlb__T_2143 = tlb__T_2142[0]; // @[Misc.scala 180:37:freechips.rocketchip.system.DefaultRV32Config.fir@180211.4]
  assign tlb__T_2145 = tlb__T_2142[1]; // @[Misc.scala 181:39:freechips.rocketchip.system.DefaultRV32Config.fir@180213.4]
  assign tlb__T_2147 = tlb__T_2143 | tlb__T_2145; // @[Misc.scala 182:16:freechips.rocketchip.system.DefaultRV32Config.fir@180215.4]
  assign tlb__T_2149 = tlb__T_2143 & tlb__T_2145; // @[Misc.scala 182:61:freechips.rocketchip.system.DefaultRV32Config.fir@180217.4]
  assign tlb__T_2151 = tlb__T_2140 | tlb__T_2147; // @[Misc.scala 182:16:freechips.rocketchip.system.DefaultRV32Config.fir@180219.4]
  assign tlb__T_2153 = tlb__T_2140 & tlb__T_2147; // @[Misc.scala 182:61:freechips.rocketchip.system.DefaultRV32Config.fir@180221.4]
  assign tlb__T_2154 = tlb__T_2149 | tlb__T_2153; // @[Misc.scala 182:49:freechips.rocketchip.system.DefaultRV32Config.fir@180222.4]
  assign tlb__T_2155 = tlb__T_2138[6:3]; // @[Misc.scala 181:39:freechips.rocketchip.system.DefaultRV32Config.fir@180223.4]
  assign tlb__T_2156 = tlb__T_2155[1:0]; // @[Misc.scala 180:37:freechips.rocketchip.system.DefaultRV32Config.fir@180224.4]
  assign tlb__T_2157 = tlb__T_2156[0]; // @[Misc.scala 180:37:freechips.rocketchip.system.DefaultRV32Config.fir@180225.4]
  assign tlb__T_2159 = tlb__T_2156[1]; // @[Misc.scala 181:39:freechips.rocketchip.system.DefaultRV32Config.fir@180227.4]
  assign tlb__T_2161 = tlb__T_2157 | tlb__T_2159; // @[Misc.scala 182:16:freechips.rocketchip.system.DefaultRV32Config.fir@180229.4]
  assign tlb__T_2163 = tlb__T_2157 & tlb__T_2159; // @[Misc.scala 182:61:freechips.rocketchip.system.DefaultRV32Config.fir@180231.4]
  assign tlb__T_2165 = tlb__T_2155[3:2]; // @[Misc.scala 181:39:freechips.rocketchip.system.DefaultRV32Config.fir@180233.4]
  assign tlb__T_2166 = tlb__T_2165[0]; // @[Misc.scala 180:37:freechips.rocketchip.system.DefaultRV32Config.fir@180234.4]
  assign tlb__T_2168 = tlb__T_2165[1]; // @[Misc.scala 181:39:freechips.rocketchip.system.DefaultRV32Config.fir@180236.4]
  assign tlb__T_2170 = tlb__T_2166 | tlb__T_2168; // @[Misc.scala 182:16:freechips.rocketchip.system.DefaultRV32Config.fir@180238.4]
  assign tlb__T_2172 = tlb__T_2166 & tlb__T_2168; // @[Misc.scala 182:61:freechips.rocketchip.system.DefaultRV32Config.fir@180240.4]
  assign tlb__T_2174 = tlb__T_2161 | tlb__T_2170; // @[Misc.scala 182:16:freechips.rocketchip.system.DefaultRV32Config.fir@180242.4]
  assign tlb__T_2175 = tlb__T_2163 | tlb__T_2172; // @[Misc.scala 182:37:freechips.rocketchip.system.DefaultRV32Config.fir@180243.4]
  assign tlb__T_2176 = tlb__T_2161 & tlb__T_2170; // @[Misc.scala 182:61:freechips.rocketchip.system.DefaultRV32Config.fir@180244.4]
  assign tlb__T_2177 = tlb__T_2175 | tlb__T_2176; // @[Misc.scala 182:49:freechips.rocketchip.system.DefaultRV32Config.fir@180245.4]
  assign tlb__T_2178 = tlb__T_2151 | tlb__T_2174; // @[Misc.scala 182:16:freechips.rocketchip.system.DefaultRV32Config.fir@180246.4]
  assign tlb__T_2179 = tlb__T_2154 | tlb__T_2177; // @[Misc.scala 182:37:freechips.rocketchip.system.DefaultRV32Config.fir@180247.4]
  assign tlb__T_2180 = tlb__T_2151 & tlb__T_2174; // @[Misc.scala 182:61:freechips.rocketchip.system.DefaultRV32Config.fir@180248.4]
  assign tlb__T_2181 = tlb__T_2179 | tlb__T_2180; // @[Misc.scala 182:49:freechips.rocketchip.system.DefaultRV32Config.fir@180249.4]
  assign tlb__T_2183 = tlb__T_2137 | tlb__T_2181; // @[Misc.scala 182:37:freechips.rocketchip.system.DefaultRV32Config.fir@180251.4]
  assign tlb__T_2184 = tlb__T_2134 & tlb__T_2178; // @[Misc.scala 182:61:freechips.rocketchip.system.DefaultRV32Config.fir@180252.4]
  assign tlb_multipleHits = tlb__T_2183 | tlb__T_2184; // @[Misc.scala 182:49:freechips.rocketchip.system.DefaultRV32Config.fir@180253.4]
  assign tlb__T_2187 = tlb_pf_ld_array & tlb_hits; // @[TLB.scala 333:57:freechips.rocketchip.system.DefaultRV32Config.fir@180257.4]
  assign tlb__T_2191 = tlb_pf_st_array & tlb_hits; // @[TLB.scala 334:64:freechips.rocketchip.system.DefaultRV32Config.fir@180262.4]
  assign tlb__T_2197 = tlb_ae_ld_array & tlb_hits; // @[TLB.scala 336:33:freechips.rocketchip.system.DefaultRV32Config.fir@180270.4]
  assign tlb__T_2199 = tlb_ae_st_array & tlb_hits; // @[TLB.scala 337:33:freechips.rocketchip.system.DefaultRV32Config.fir@180273.4]
  assign tlb__T_2204 = tlb_ma_ld_array & tlb_hits; // @[TLB.scala 339:33:freechips.rocketchip.system.DefaultRV32Config.fir@180280.4]
  assign tlb__T_2206 = tlb_ma_st_array & tlb_hits; // @[TLB.scala 340:33:freechips.rocketchip.system.DefaultRV32Config.fir@180283.4]
  assign tlb__T_2208 = tlb_c_array & tlb_hits; // @[TLB.scala 342:33:freechips.rocketchip.system.DefaultRV32Config.fir@180287.4]
  assign tlb__T_2215 = tlb_io_ptw_resp_valid | tlb_tlb_miss; // @[TLB.scala 345:29:freechips.rocketchip.system.DefaultRV32Config.fir@180297.4]
  assign tlb__T_2221 = tlb_io_req_ready & tlb_io_req_valid; // @[Decoupled.scala 40:37:freechips.rocketchip.system.DefaultRV32Config.fir@180308.4]
  assign tlb__T_2222 = tlb__T_2221 & tlb_tlb_miss; // @[TLB.scala 354:25:freechips.rocketchip.system.DefaultRV32Config.fir@180309.4]
  assign tlb__T_2223 = tlb__T_2008[2]; // @[Replacement.scala 233:38:freechips.rocketchip.system.DefaultRV32Config.fir@180313.6]
  assign tlb__T_2228 = tlb__T_2223 ? tlb__T_2089 : tlb__T_2090; // @[Replacement.scala 240:16:freechips.rocketchip.system.DefaultRV32Config.fir@180318.6]
  assign tlb__T_2229 = {tlb__T_2223,tlb__T_2228}; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@180319.6]
  assign tlb__T_2232 = {tlb_superpage_entries_3_valid_0,tlb_superpage_entries_2_valid_0,tlb_superpage_entries_1_valid_0,tlb_superpage_entries_0_valid_0}; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@180322.6]
  assign tlb__T_2233 = &tlb__T_2232; // @[TLB.scala 402:16:freechips.rocketchip.system.DefaultRV32Config.fir@180323.6]
  assign tlb__T_2234 = ~tlb__T_2232; // @[TLB.scala 402:43:freechips.rocketchip.system.DefaultRV32Config.fir@180324.6]
  assign tlb__T_2235 = tlb__T_2234[0]; // @[OneHot.scala 47:40:freechips.rocketchip.system.DefaultRV32Config.fir@180325.6]
  assign tlb__T_2236 = tlb__T_2234[1]; // @[OneHot.scala 47:40:freechips.rocketchip.system.DefaultRV32Config.fir@180326.6]
  assign tlb__T_2237 = tlb__T_2234[2]; // @[OneHot.scala 47:40:freechips.rocketchip.system.DefaultRV32Config.fir@180327.6]
  assign tlb__T_2243 = tlb__T_2007[6]; // @[Replacement.scala 233:38:freechips.rocketchip.system.DefaultRV32Config.fir@180334.6]
  assign tlb__T_2246 = tlb__T_2038[2]; // @[Replacement.scala 233:38:freechips.rocketchip.system.DefaultRV32Config.fir@180337.6]
  assign tlb__T_2251 = tlb__T_2246 ? tlb__T_2043 : tlb__T_2044; // @[Replacement.scala 240:16:freechips.rocketchip.system.DefaultRV32Config.fir@180342.6]
  assign tlb__T_2252 = {tlb__T_2246,tlb__T_2251}; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@180343.6]
  assign tlb__T_2253 = tlb__T_2039[2]; // @[Replacement.scala 233:38:freechips.rocketchip.system.DefaultRV32Config.fir@180344.6]
  assign tlb__T_2258 = tlb__T_2253 ? tlb__T_2059 : tlb__T_2060; // @[Replacement.scala 240:16:freechips.rocketchip.system.DefaultRV32Config.fir@180349.6]
  assign tlb__T_2259 = {tlb__T_2253,tlb__T_2258}; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@180350.6]
  assign tlb__T_2260 = tlb__T_2243 ? tlb__T_2252 : tlb__T_2259; // @[Replacement.scala 240:16:freechips.rocketchip.system.DefaultRV32Config.fir@180351.6]
  assign tlb__T_2261 = {tlb__T_2243,tlb__T_2260}; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@180352.6]
  assign tlb__T_2292 = {tlb__T_454,tlb__T_448,tlb__T_442,tlb__T_436,tlb__T_430,tlb__T_424,tlb__T_418,tlb__T_412}; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@180383.6]
  assign tlb__T_2293 = &tlb__T_2292; // @[TLB.scala 402:16:freechips.rocketchip.system.DefaultRV32Config.fir@180384.6]
  assign tlb__T_2294 = ~tlb__T_2292; // @[TLB.scala 402:43:freechips.rocketchip.system.DefaultRV32Config.fir@180385.6]
  assign tlb__T_2295 = tlb__T_2294[0]; // @[OneHot.scala 47:40:freechips.rocketchip.system.DefaultRV32Config.fir@180386.6]
  assign tlb__T_2296 = tlb__T_2294[1]; // @[OneHot.scala 47:40:freechips.rocketchip.system.DefaultRV32Config.fir@180387.6]
  assign tlb__T_2297 = tlb__T_2294[2]; // @[OneHot.scala 47:40:freechips.rocketchip.system.DefaultRV32Config.fir@180388.6]
  assign tlb__T_2298 = tlb__T_2294[3]; // @[OneHot.scala 47:40:freechips.rocketchip.system.DefaultRV32Config.fir@180389.6]
  assign tlb__T_2299 = tlb__T_2294[4]; // @[OneHot.scala 47:40:freechips.rocketchip.system.DefaultRV32Config.fir@180390.6]
  assign tlb__T_2300 = tlb__T_2294[5]; // @[OneHot.scala 47:40:freechips.rocketchip.system.DefaultRV32Config.fir@180391.6]
  assign tlb__T_2301 = tlb__T_2294[6]; // @[OneHot.scala 47:40:freechips.rocketchip.system.DefaultRV32Config.fir@180392.6]
  assign tlb__T_2338 = tlb_state == 2'h2; // @[TLB.scala 368:17:freechips.rocketchip.system.DefaultRV32Config.fir@180444.4]
  assign tlb__T_2339 = tlb__T_2338 & tlb_io_sfence_valid; // @[TLB.scala 368:28:freechips.rocketchip.system.DefaultRV32Config.fir@180445.4]
  assign tlb__T_2340 = ~tlb_io_sfence_bits_rs1; // @[TLB.scala 376:14:freechips.rocketchip.system.DefaultRV32Config.fir@180453.6]
  assign tlb__T_2341 = tlb_io_sfence_bits_addr[31:12]; // @[TLB.scala 376:58:freechips.rocketchip.system.DefaultRV32Config.fir@180454.6]
  assign tlb__T_2342 = tlb__T_2341 == tlb_vpn; // @[TLB.scala 376:72:freechips.rocketchip.system.DefaultRV32Config.fir@180455.6]
  assign tlb__T_2343 = tlb__T_2340 | tlb__T_2342; // @[TLB.scala 376:34:freechips.rocketchip.system.DefaultRV32Config.fir@180456.6]
  assign tlb__T_2345 = tlb__T_2343 | tlb_reset; // @[TLB.scala 376:13:freechips.rocketchip.system.DefaultRV32Config.fir@180458.6]
  assign tlb__T_2346 = ~tlb__T_2345; // @[TLB.scala 376:13:freechips.rocketchip.system.DefaultRV32Config.fir@180459.6]
  assign tlb__T_2352 = tlb__T_413[19:10]; // @[TLB.scala 135:26:freechips.rocketchip.system.DefaultRV32Config.fir@180473.8]
  assign tlb__T_2353 = tlb__T_2352 == 10'h0; // @[TLB.scala 135:61:freechips.rocketchip.system.DefaultRV32Config.fir@180474.8]
  assign tlb__T_2356 = tlb_sectored_entries_0_data_0[0]; // @[TLB.scala 83:39:freechips.rocketchip.system.DefaultRV32Config.fir@180481.10]
  assign tlb__T_2369 = tlb_sectored_entries_0_data_0[13]; // @[TLB.scala 83:39:freechips.rocketchip.system.DefaultRV32Config.fir@180507.10]
  assign tlb__T_2374 = tlb_sectored_entries_0_data_1[0]; // @[TLB.scala 83:39:freechips.rocketchip.system.DefaultRV32Config.fir@180518.10]
  assign tlb__T_2387 = tlb_sectored_entries_0_data_1[13]; // @[TLB.scala 83:39:freechips.rocketchip.system.DefaultRV32Config.fir@180544.10]
  assign tlb__T_2392 = tlb_sectored_entries_0_data_2[0]; // @[TLB.scala 83:39:freechips.rocketchip.system.DefaultRV32Config.fir@180555.10]
  assign tlb__T_2405 = tlb_sectored_entries_0_data_2[13]; // @[TLB.scala 83:39:freechips.rocketchip.system.DefaultRV32Config.fir@180581.10]
  assign tlb__T_2410 = tlb_sectored_entries_0_data_3[0]; // @[TLB.scala 83:39:freechips.rocketchip.system.DefaultRV32Config.fir@180592.10]
  assign tlb__T_2423 = tlb_sectored_entries_0_data_3[13]; // @[TLB.scala 83:39:freechips.rocketchip.system.DefaultRV32Config.fir@180618.10]
  assign tlb__T_2498 = ~tlb__T_2369; // @[TLB.scala 143:13:freechips.rocketchip.system.DefaultRV32Config.fir@180788.10]
  assign tlb__GEN_648 = tlb__T_2498 ? 1'h0 : tlb__GEN_472; // @[TLB.scala 143:19:freechips.rocketchip.system.DefaultRV32Config.fir@180789.10]
  assign tlb__T_2499 = ~tlb__T_2387; // @[TLB.scala 143:13:freechips.rocketchip.system.DefaultRV32Config.fir@180792.10]
  assign tlb__GEN_649 = tlb__T_2499 ? 1'h0 : tlb__GEN_473; // @[TLB.scala 143:19:freechips.rocketchip.system.DefaultRV32Config.fir@180793.10]
  assign tlb__T_2500 = ~tlb__T_2405; // @[TLB.scala 143:13:freechips.rocketchip.system.DefaultRV32Config.fir@180796.10]
  assign tlb__GEN_650 = tlb__T_2500 ? 1'h0 : tlb__GEN_474; // @[TLB.scala 143:19:freechips.rocketchip.system.DefaultRV32Config.fir@180797.10]
  assign tlb__T_2501 = ~tlb__T_2423; // @[TLB.scala 143:13:freechips.rocketchip.system.DefaultRV32Config.fir@180800.10]
  assign tlb__GEN_651 = tlb__T_2501 ? 1'h0 : tlb__GEN_475; // @[TLB.scala 143:19:freechips.rocketchip.system.DefaultRV32Config.fir@180801.10]
  assign tlb__GEN_652 = tlb_io_sfence_bits_rs2 & tlb__GEN_648; // @[TLB.scala 379:40:freechips.rocketchip.system.DefaultRV32Config.fir@180639.8]
  assign tlb__GEN_653 = tlb_io_sfence_bits_rs2 & tlb__GEN_649; // @[TLB.scala 379:40:freechips.rocketchip.system.DefaultRV32Config.fir@180639.8]
  assign tlb__GEN_654 = tlb_io_sfence_bits_rs2 & tlb__GEN_650; // @[TLB.scala 379:40:freechips.rocketchip.system.DefaultRV32Config.fir@180639.8]
  assign tlb__GEN_655 = tlb_io_sfence_bits_rs2 & tlb__GEN_651; // @[TLB.scala 379:40:freechips.rocketchip.system.DefaultRV32Config.fir@180639.8]
  assign tlb__T_2507 = tlb__T_419[19:10]; // @[TLB.scala 135:26:freechips.rocketchip.system.DefaultRV32Config.fir@180820.8]
  assign tlb__T_2508 = tlb__T_2507 == 10'h0; // @[TLB.scala 135:61:freechips.rocketchip.system.DefaultRV32Config.fir@180821.8]
  assign tlb__T_2511 = tlb_sectored_entries_1_data_0[0]; // @[TLB.scala 83:39:freechips.rocketchip.system.DefaultRV32Config.fir@180828.10]
  assign tlb__T_2524 = tlb_sectored_entries_1_data_0[13]; // @[TLB.scala 83:39:freechips.rocketchip.system.DefaultRV32Config.fir@180854.10]
  assign tlb__T_2529 = tlb_sectored_entries_1_data_1[0]; // @[TLB.scala 83:39:freechips.rocketchip.system.DefaultRV32Config.fir@180865.10]
  assign tlb__T_2542 = tlb_sectored_entries_1_data_1[13]; // @[TLB.scala 83:39:freechips.rocketchip.system.DefaultRV32Config.fir@180891.10]
  assign tlb__T_2547 = tlb_sectored_entries_1_data_2[0]; // @[TLB.scala 83:39:freechips.rocketchip.system.DefaultRV32Config.fir@180902.10]
  assign tlb__T_2560 = tlb_sectored_entries_1_data_2[13]; // @[TLB.scala 83:39:freechips.rocketchip.system.DefaultRV32Config.fir@180928.10]
  assign tlb__T_2565 = tlb_sectored_entries_1_data_3[0]; // @[TLB.scala 83:39:freechips.rocketchip.system.DefaultRV32Config.fir@180939.10]
  assign tlb__T_2578 = tlb_sectored_entries_1_data_3[13]; // @[TLB.scala 83:39:freechips.rocketchip.system.DefaultRV32Config.fir@180965.10]
  assign tlb__T_2653 = ~tlb__T_2524; // @[TLB.scala 143:13:freechips.rocketchip.system.DefaultRV32Config.fir@181135.10]
  assign tlb__GEN_676 = tlb__T_2653 ? 1'h0 : tlb__GEN_482; // @[TLB.scala 143:19:freechips.rocketchip.system.DefaultRV32Config.fir@181136.10]
  assign tlb__T_2654 = ~tlb__T_2542; // @[TLB.scala 143:13:freechips.rocketchip.system.DefaultRV32Config.fir@181139.10]
  assign tlb__GEN_677 = tlb__T_2654 ? 1'h0 : tlb__GEN_483; // @[TLB.scala 143:19:freechips.rocketchip.system.DefaultRV32Config.fir@181140.10]
  assign tlb__T_2655 = ~tlb__T_2560; // @[TLB.scala 143:13:freechips.rocketchip.system.DefaultRV32Config.fir@181143.10]
  assign tlb__GEN_678 = tlb__T_2655 ? 1'h0 : tlb__GEN_484; // @[TLB.scala 143:19:freechips.rocketchip.system.DefaultRV32Config.fir@181144.10]
  assign tlb__T_2656 = ~tlb__T_2578; // @[TLB.scala 143:13:freechips.rocketchip.system.DefaultRV32Config.fir@181147.10]
  assign tlb__GEN_679 = tlb__T_2656 ? 1'h0 : tlb__GEN_485; // @[TLB.scala 143:19:freechips.rocketchip.system.DefaultRV32Config.fir@181148.10]
  assign tlb__GEN_680 = tlb_io_sfence_bits_rs2 & tlb__GEN_676; // @[TLB.scala 379:40:freechips.rocketchip.system.DefaultRV32Config.fir@180986.8]
  assign tlb__GEN_681 = tlb_io_sfence_bits_rs2 & tlb__GEN_677; // @[TLB.scala 379:40:freechips.rocketchip.system.DefaultRV32Config.fir@180986.8]
  assign tlb__GEN_682 = tlb_io_sfence_bits_rs2 & tlb__GEN_678; // @[TLB.scala 379:40:freechips.rocketchip.system.DefaultRV32Config.fir@180986.8]
  assign tlb__GEN_683 = tlb_io_sfence_bits_rs2 & tlb__GEN_679; // @[TLB.scala 379:40:freechips.rocketchip.system.DefaultRV32Config.fir@180986.8]
  assign tlb__T_2662 = tlb__T_425[19:10]; // @[TLB.scala 135:26:freechips.rocketchip.system.DefaultRV32Config.fir@181167.8]
  assign tlb__T_2663 = tlb__T_2662 == 10'h0; // @[TLB.scala 135:61:freechips.rocketchip.system.DefaultRV32Config.fir@181168.8]
  assign tlb__T_2666 = tlb_sectored_entries_2_data_0[0]; // @[TLB.scala 83:39:freechips.rocketchip.system.DefaultRV32Config.fir@181175.10]
  assign tlb__T_2679 = tlb_sectored_entries_2_data_0[13]; // @[TLB.scala 83:39:freechips.rocketchip.system.DefaultRV32Config.fir@181201.10]
  assign tlb__T_2684 = tlb_sectored_entries_2_data_1[0]; // @[TLB.scala 83:39:freechips.rocketchip.system.DefaultRV32Config.fir@181212.10]
  assign tlb__T_2697 = tlb_sectored_entries_2_data_1[13]; // @[TLB.scala 83:39:freechips.rocketchip.system.DefaultRV32Config.fir@181238.10]
  assign tlb__T_2702 = tlb_sectored_entries_2_data_2[0]; // @[TLB.scala 83:39:freechips.rocketchip.system.DefaultRV32Config.fir@181249.10]
  assign tlb__T_2715 = tlb_sectored_entries_2_data_2[13]; // @[TLB.scala 83:39:freechips.rocketchip.system.DefaultRV32Config.fir@181275.10]
  assign tlb__T_2720 = tlb_sectored_entries_2_data_3[0]; // @[TLB.scala 83:39:freechips.rocketchip.system.DefaultRV32Config.fir@181286.10]
  assign tlb__T_2733 = tlb_sectored_entries_2_data_3[13]; // @[TLB.scala 83:39:freechips.rocketchip.system.DefaultRV32Config.fir@181312.10]
  assign tlb__T_2808 = ~tlb__T_2679; // @[TLB.scala 143:13:freechips.rocketchip.system.DefaultRV32Config.fir@181482.10]
  assign tlb__GEN_704 = tlb__T_2808 ? 1'h0 : tlb__GEN_492; // @[TLB.scala 143:19:freechips.rocketchip.system.DefaultRV32Config.fir@181483.10]
  assign tlb__T_2809 = ~tlb__T_2697; // @[TLB.scala 143:13:freechips.rocketchip.system.DefaultRV32Config.fir@181486.10]
  assign tlb__GEN_705 = tlb__T_2809 ? 1'h0 : tlb__GEN_493; // @[TLB.scala 143:19:freechips.rocketchip.system.DefaultRV32Config.fir@181487.10]
  assign tlb__T_2810 = ~tlb__T_2715; // @[TLB.scala 143:13:freechips.rocketchip.system.DefaultRV32Config.fir@181490.10]
  assign tlb__GEN_706 = tlb__T_2810 ? 1'h0 : tlb__GEN_494; // @[TLB.scala 143:19:freechips.rocketchip.system.DefaultRV32Config.fir@181491.10]
  assign tlb__T_2811 = ~tlb__T_2733; // @[TLB.scala 143:13:freechips.rocketchip.system.DefaultRV32Config.fir@181494.10]
  assign tlb__GEN_707 = tlb__T_2811 ? 1'h0 : tlb__GEN_495; // @[TLB.scala 143:19:freechips.rocketchip.system.DefaultRV32Config.fir@181495.10]
  assign tlb__GEN_708 = tlb_io_sfence_bits_rs2 & tlb__GEN_704; // @[TLB.scala 379:40:freechips.rocketchip.system.DefaultRV32Config.fir@181333.8]
  assign tlb__GEN_709 = tlb_io_sfence_bits_rs2 & tlb__GEN_705; // @[TLB.scala 379:40:freechips.rocketchip.system.DefaultRV32Config.fir@181333.8]
  assign tlb__GEN_710 = tlb_io_sfence_bits_rs2 & tlb__GEN_706; // @[TLB.scala 379:40:freechips.rocketchip.system.DefaultRV32Config.fir@181333.8]
  assign tlb__GEN_711 = tlb_io_sfence_bits_rs2 & tlb__GEN_707; // @[TLB.scala 379:40:freechips.rocketchip.system.DefaultRV32Config.fir@181333.8]
  assign tlb__T_2817 = tlb__T_431[19:10]; // @[TLB.scala 135:26:freechips.rocketchip.system.DefaultRV32Config.fir@181514.8]
  assign tlb__T_2818 = tlb__T_2817 == 10'h0; // @[TLB.scala 135:61:freechips.rocketchip.system.DefaultRV32Config.fir@181515.8]
  assign tlb__T_2821 = tlb_sectored_entries_3_data_0[0]; // @[TLB.scala 83:39:freechips.rocketchip.system.DefaultRV32Config.fir@181522.10]
  assign tlb__T_2834 = tlb_sectored_entries_3_data_0[13]; // @[TLB.scala 83:39:freechips.rocketchip.system.DefaultRV32Config.fir@181548.10]
  assign tlb__T_2839 = tlb_sectored_entries_3_data_1[0]; // @[TLB.scala 83:39:freechips.rocketchip.system.DefaultRV32Config.fir@181559.10]
  assign tlb__T_2852 = tlb_sectored_entries_3_data_1[13]; // @[TLB.scala 83:39:freechips.rocketchip.system.DefaultRV32Config.fir@181585.10]
  assign tlb__T_2857 = tlb_sectored_entries_3_data_2[0]; // @[TLB.scala 83:39:freechips.rocketchip.system.DefaultRV32Config.fir@181596.10]
  assign tlb__T_2870 = tlb_sectored_entries_3_data_2[13]; // @[TLB.scala 83:39:freechips.rocketchip.system.DefaultRV32Config.fir@181622.10]
  assign tlb__T_2875 = tlb_sectored_entries_3_data_3[0]; // @[TLB.scala 83:39:freechips.rocketchip.system.DefaultRV32Config.fir@181633.10]
  assign tlb__T_2888 = tlb_sectored_entries_3_data_3[13]; // @[TLB.scala 83:39:freechips.rocketchip.system.DefaultRV32Config.fir@181659.10]
  assign tlb__T_2963 = ~tlb__T_2834; // @[TLB.scala 143:13:freechips.rocketchip.system.DefaultRV32Config.fir@181829.10]
  assign tlb__GEN_732 = tlb__T_2963 ? 1'h0 : tlb__GEN_502; // @[TLB.scala 143:19:freechips.rocketchip.system.DefaultRV32Config.fir@181830.10]
  assign tlb__T_2964 = ~tlb__T_2852; // @[TLB.scala 143:13:freechips.rocketchip.system.DefaultRV32Config.fir@181833.10]
  assign tlb__GEN_733 = tlb__T_2964 ? 1'h0 : tlb__GEN_503; // @[TLB.scala 143:19:freechips.rocketchip.system.DefaultRV32Config.fir@181834.10]
  assign tlb__T_2965 = ~tlb__T_2870; // @[TLB.scala 143:13:freechips.rocketchip.system.DefaultRV32Config.fir@181837.10]
  assign tlb__GEN_734 = tlb__T_2965 ? 1'h0 : tlb__GEN_504; // @[TLB.scala 143:19:freechips.rocketchip.system.DefaultRV32Config.fir@181838.10]
  assign tlb__T_2966 = ~tlb__T_2888; // @[TLB.scala 143:13:freechips.rocketchip.system.DefaultRV32Config.fir@181841.10]
  assign tlb__GEN_735 = tlb__T_2966 ? 1'h0 : tlb__GEN_505; // @[TLB.scala 143:19:freechips.rocketchip.system.DefaultRV32Config.fir@181842.10]
  assign tlb__GEN_736 = tlb_io_sfence_bits_rs2 & tlb__GEN_732; // @[TLB.scala 379:40:freechips.rocketchip.system.DefaultRV32Config.fir@181680.8]
  assign tlb__GEN_737 = tlb_io_sfence_bits_rs2 & tlb__GEN_733; // @[TLB.scala 379:40:freechips.rocketchip.system.DefaultRV32Config.fir@181680.8]
  assign tlb__GEN_738 = tlb_io_sfence_bits_rs2 & tlb__GEN_734; // @[TLB.scala 379:40:freechips.rocketchip.system.DefaultRV32Config.fir@181680.8]
  assign tlb__GEN_739 = tlb_io_sfence_bits_rs2 & tlb__GEN_735; // @[TLB.scala 379:40:freechips.rocketchip.system.DefaultRV32Config.fir@181680.8]
  assign tlb__T_2972 = tlb__T_437[19:10]; // @[TLB.scala 135:26:freechips.rocketchip.system.DefaultRV32Config.fir@181861.8]
  assign tlb__T_2973 = tlb__T_2972 == 10'h0; // @[TLB.scala 135:61:freechips.rocketchip.system.DefaultRV32Config.fir@181862.8]
  assign tlb__T_2976 = tlb_sectored_entries_4_data_0[0]; // @[TLB.scala 83:39:freechips.rocketchip.system.DefaultRV32Config.fir@181869.10]
  assign tlb__T_2989 = tlb_sectored_entries_4_data_0[13]; // @[TLB.scala 83:39:freechips.rocketchip.system.DefaultRV32Config.fir@181895.10]
  assign tlb__T_2994 = tlb_sectored_entries_4_data_1[0]; // @[TLB.scala 83:39:freechips.rocketchip.system.DefaultRV32Config.fir@181906.10]
  assign tlb__T_3007 = tlb_sectored_entries_4_data_1[13]; // @[TLB.scala 83:39:freechips.rocketchip.system.DefaultRV32Config.fir@181932.10]
  assign tlb__T_3012 = tlb_sectored_entries_4_data_2[0]; // @[TLB.scala 83:39:freechips.rocketchip.system.DefaultRV32Config.fir@181943.10]
  assign tlb__T_3025 = tlb_sectored_entries_4_data_2[13]; // @[TLB.scala 83:39:freechips.rocketchip.system.DefaultRV32Config.fir@181969.10]
  assign tlb__T_3030 = tlb_sectored_entries_4_data_3[0]; // @[TLB.scala 83:39:freechips.rocketchip.system.DefaultRV32Config.fir@181980.10]
  assign tlb__T_3043 = tlb_sectored_entries_4_data_3[13]; // @[TLB.scala 83:39:freechips.rocketchip.system.DefaultRV32Config.fir@182006.10]
  assign tlb__T_3118 = ~tlb__T_2989; // @[TLB.scala 143:13:freechips.rocketchip.system.DefaultRV32Config.fir@182176.10]
  assign tlb__GEN_760 = tlb__T_3118 ? 1'h0 : tlb__GEN_512; // @[TLB.scala 143:19:freechips.rocketchip.system.DefaultRV32Config.fir@182177.10]
  assign tlb__T_3119 = ~tlb__T_3007; // @[TLB.scala 143:13:freechips.rocketchip.system.DefaultRV32Config.fir@182180.10]
  assign tlb__GEN_761 = tlb__T_3119 ? 1'h0 : tlb__GEN_513; // @[TLB.scala 143:19:freechips.rocketchip.system.DefaultRV32Config.fir@182181.10]
  assign tlb__T_3120 = ~tlb__T_3025; // @[TLB.scala 143:13:freechips.rocketchip.system.DefaultRV32Config.fir@182184.10]
  assign tlb__GEN_762 = tlb__T_3120 ? 1'h0 : tlb__GEN_514; // @[TLB.scala 143:19:freechips.rocketchip.system.DefaultRV32Config.fir@182185.10]
  assign tlb__T_3121 = ~tlb__T_3043; // @[TLB.scala 143:13:freechips.rocketchip.system.DefaultRV32Config.fir@182188.10]
  assign tlb__GEN_763 = tlb__T_3121 ? 1'h0 : tlb__GEN_515; // @[TLB.scala 143:19:freechips.rocketchip.system.DefaultRV32Config.fir@182189.10]
  assign tlb__GEN_764 = tlb_io_sfence_bits_rs2 & tlb__GEN_760; // @[TLB.scala 379:40:freechips.rocketchip.system.DefaultRV32Config.fir@182027.8]
  assign tlb__GEN_765 = tlb_io_sfence_bits_rs2 & tlb__GEN_761; // @[TLB.scala 379:40:freechips.rocketchip.system.DefaultRV32Config.fir@182027.8]
  assign tlb__GEN_766 = tlb_io_sfence_bits_rs2 & tlb__GEN_762; // @[TLB.scala 379:40:freechips.rocketchip.system.DefaultRV32Config.fir@182027.8]
  assign tlb__GEN_767 = tlb_io_sfence_bits_rs2 & tlb__GEN_763; // @[TLB.scala 379:40:freechips.rocketchip.system.DefaultRV32Config.fir@182027.8]
  assign tlb__T_3127 = tlb__T_443[19:10]; // @[TLB.scala 135:26:freechips.rocketchip.system.DefaultRV32Config.fir@182208.8]
  assign tlb__T_3128 = tlb__T_3127 == 10'h0; // @[TLB.scala 135:61:freechips.rocketchip.system.DefaultRV32Config.fir@182209.8]
  assign tlb__T_3131 = tlb_sectored_entries_5_data_0[0]; // @[TLB.scala 83:39:freechips.rocketchip.system.DefaultRV32Config.fir@182216.10]
  assign tlb__T_3144 = tlb_sectored_entries_5_data_0[13]; // @[TLB.scala 83:39:freechips.rocketchip.system.DefaultRV32Config.fir@182242.10]
  assign tlb__T_3149 = tlb_sectored_entries_5_data_1[0]; // @[TLB.scala 83:39:freechips.rocketchip.system.DefaultRV32Config.fir@182253.10]
  assign tlb__T_3162 = tlb_sectored_entries_5_data_1[13]; // @[TLB.scala 83:39:freechips.rocketchip.system.DefaultRV32Config.fir@182279.10]
  assign tlb__T_3167 = tlb_sectored_entries_5_data_2[0]; // @[TLB.scala 83:39:freechips.rocketchip.system.DefaultRV32Config.fir@182290.10]
  assign tlb__T_3180 = tlb_sectored_entries_5_data_2[13]; // @[TLB.scala 83:39:freechips.rocketchip.system.DefaultRV32Config.fir@182316.10]
  assign tlb__T_3185 = tlb_sectored_entries_5_data_3[0]; // @[TLB.scala 83:39:freechips.rocketchip.system.DefaultRV32Config.fir@182327.10]
  assign tlb__T_3198 = tlb_sectored_entries_5_data_3[13]; // @[TLB.scala 83:39:freechips.rocketchip.system.DefaultRV32Config.fir@182353.10]
  assign tlb__T_3273 = ~tlb__T_3144; // @[TLB.scala 143:13:freechips.rocketchip.system.DefaultRV32Config.fir@182523.10]
  assign tlb__GEN_788 = tlb__T_3273 ? 1'h0 : tlb__GEN_522; // @[TLB.scala 143:19:freechips.rocketchip.system.DefaultRV32Config.fir@182524.10]
  assign tlb__T_3274 = ~tlb__T_3162; // @[TLB.scala 143:13:freechips.rocketchip.system.DefaultRV32Config.fir@182527.10]
  assign tlb__GEN_789 = tlb__T_3274 ? 1'h0 : tlb__GEN_523; // @[TLB.scala 143:19:freechips.rocketchip.system.DefaultRV32Config.fir@182528.10]
  assign tlb__T_3275 = ~tlb__T_3180; // @[TLB.scala 143:13:freechips.rocketchip.system.DefaultRV32Config.fir@182531.10]
  assign tlb__GEN_790 = tlb__T_3275 ? 1'h0 : tlb__GEN_524; // @[TLB.scala 143:19:freechips.rocketchip.system.DefaultRV32Config.fir@182532.10]
  assign tlb__T_3276 = ~tlb__T_3198; // @[TLB.scala 143:13:freechips.rocketchip.system.DefaultRV32Config.fir@182535.10]
  assign tlb__GEN_791 = tlb__T_3276 ? 1'h0 : tlb__GEN_525; // @[TLB.scala 143:19:freechips.rocketchip.system.DefaultRV32Config.fir@182536.10]
  assign tlb__GEN_792 = tlb_io_sfence_bits_rs2 & tlb__GEN_788; // @[TLB.scala 379:40:freechips.rocketchip.system.DefaultRV32Config.fir@182374.8]
  assign tlb__GEN_793 = tlb_io_sfence_bits_rs2 & tlb__GEN_789; // @[TLB.scala 379:40:freechips.rocketchip.system.DefaultRV32Config.fir@182374.8]
  assign tlb__GEN_794 = tlb_io_sfence_bits_rs2 & tlb__GEN_790; // @[TLB.scala 379:40:freechips.rocketchip.system.DefaultRV32Config.fir@182374.8]
  assign tlb__GEN_795 = tlb_io_sfence_bits_rs2 & tlb__GEN_791; // @[TLB.scala 379:40:freechips.rocketchip.system.DefaultRV32Config.fir@182374.8]
  assign tlb__T_3282 = tlb__T_449[19:10]; // @[TLB.scala 135:26:freechips.rocketchip.system.DefaultRV32Config.fir@182555.8]
  assign tlb__T_3283 = tlb__T_3282 == 10'h0; // @[TLB.scala 135:61:freechips.rocketchip.system.DefaultRV32Config.fir@182556.8]
  assign tlb__T_3286 = tlb_sectored_entries_6_data_0[0]; // @[TLB.scala 83:39:freechips.rocketchip.system.DefaultRV32Config.fir@182563.10]
  assign tlb__T_3299 = tlb_sectored_entries_6_data_0[13]; // @[TLB.scala 83:39:freechips.rocketchip.system.DefaultRV32Config.fir@182589.10]
  assign tlb__T_3304 = tlb_sectored_entries_6_data_1[0]; // @[TLB.scala 83:39:freechips.rocketchip.system.DefaultRV32Config.fir@182600.10]
  assign tlb__T_3317 = tlb_sectored_entries_6_data_1[13]; // @[TLB.scala 83:39:freechips.rocketchip.system.DefaultRV32Config.fir@182626.10]
  assign tlb__T_3322 = tlb_sectored_entries_6_data_2[0]; // @[TLB.scala 83:39:freechips.rocketchip.system.DefaultRV32Config.fir@182637.10]
  assign tlb__T_3335 = tlb_sectored_entries_6_data_2[13]; // @[TLB.scala 83:39:freechips.rocketchip.system.DefaultRV32Config.fir@182663.10]
  assign tlb__T_3340 = tlb_sectored_entries_6_data_3[0]; // @[TLB.scala 83:39:freechips.rocketchip.system.DefaultRV32Config.fir@182674.10]
  assign tlb__T_3353 = tlb_sectored_entries_6_data_3[13]; // @[TLB.scala 83:39:freechips.rocketchip.system.DefaultRV32Config.fir@182700.10]
  assign tlb__T_3428 = ~tlb__T_3299; // @[TLB.scala 143:13:freechips.rocketchip.system.DefaultRV32Config.fir@182870.10]
  assign tlb__GEN_816 = tlb__T_3428 ? 1'h0 : tlb__GEN_532; // @[TLB.scala 143:19:freechips.rocketchip.system.DefaultRV32Config.fir@182871.10]
  assign tlb__T_3429 = ~tlb__T_3317; // @[TLB.scala 143:13:freechips.rocketchip.system.DefaultRV32Config.fir@182874.10]
  assign tlb__GEN_817 = tlb__T_3429 ? 1'h0 : tlb__GEN_533; // @[TLB.scala 143:19:freechips.rocketchip.system.DefaultRV32Config.fir@182875.10]
  assign tlb__T_3430 = ~tlb__T_3335; // @[TLB.scala 143:13:freechips.rocketchip.system.DefaultRV32Config.fir@182878.10]
  assign tlb__GEN_818 = tlb__T_3430 ? 1'h0 : tlb__GEN_534; // @[TLB.scala 143:19:freechips.rocketchip.system.DefaultRV32Config.fir@182879.10]
  assign tlb__T_3431 = ~tlb__T_3353; // @[TLB.scala 143:13:freechips.rocketchip.system.DefaultRV32Config.fir@182882.10]
  assign tlb__GEN_819 = tlb__T_3431 ? 1'h0 : tlb__GEN_535; // @[TLB.scala 143:19:freechips.rocketchip.system.DefaultRV32Config.fir@182883.10]
  assign tlb__GEN_820 = tlb_io_sfence_bits_rs2 & tlb__GEN_816; // @[TLB.scala 379:40:freechips.rocketchip.system.DefaultRV32Config.fir@182721.8]
  assign tlb__GEN_821 = tlb_io_sfence_bits_rs2 & tlb__GEN_817; // @[TLB.scala 379:40:freechips.rocketchip.system.DefaultRV32Config.fir@182721.8]
  assign tlb__GEN_822 = tlb_io_sfence_bits_rs2 & tlb__GEN_818; // @[TLB.scala 379:40:freechips.rocketchip.system.DefaultRV32Config.fir@182721.8]
  assign tlb__GEN_823 = tlb_io_sfence_bits_rs2 & tlb__GEN_819; // @[TLB.scala 379:40:freechips.rocketchip.system.DefaultRV32Config.fir@182721.8]
  assign tlb__T_3437 = tlb__T_455[19:10]; // @[TLB.scala 135:26:freechips.rocketchip.system.DefaultRV32Config.fir@182902.8]
  assign tlb__T_3438 = tlb__T_3437 == 10'h0; // @[TLB.scala 135:61:freechips.rocketchip.system.DefaultRV32Config.fir@182903.8]
  assign tlb__T_3441 = tlb_sectored_entries_7_data_0[0]; // @[TLB.scala 83:39:freechips.rocketchip.system.DefaultRV32Config.fir@182910.10]
  assign tlb__T_3454 = tlb_sectored_entries_7_data_0[13]; // @[TLB.scala 83:39:freechips.rocketchip.system.DefaultRV32Config.fir@182936.10]
  assign tlb__T_3459 = tlb_sectored_entries_7_data_1[0]; // @[TLB.scala 83:39:freechips.rocketchip.system.DefaultRV32Config.fir@182947.10]
  assign tlb__T_3472 = tlb_sectored_entries_7_data_1[13]; // @[TLB.scala 83:39:freechips.rocketchip.system.DefaultRV32Config.fir@182973.10]
  assign tlb__T_3477 = tlb_sectored_entries_7_data_2[0]; // @[TLB.scala 83:39:freechips.rocketchip.system.DefaultRV32Config.fir@182984.10]
  assign tlb__T_3490 = tlb_sectored_entries_7_data_2[13]; // @[TLB.scala 83:39:freechips.rocketchip.system.DefaultRV32Config.fir@183010.10]
  assign tlb__T_3495 = tlb_sectored_entries_7_data_3[0]; // @[TLB.scala 83:39:freechips.rocketchip.system.DefaultRV32Config.fir@183021.10]
  assign tlb__T_3508 = tlb_sectored_entries_7_data_3[13]; // @[TLB.scala 83:39:freechips.rocketchip.system.DefaultRV32Config.fir@183047.10]
  assign tlb__T_3583 = ~tlb__T_3454; // @[TLB.scala 143:13:freechips.rocketchip.system.DefaultRV32Config.fir@183217.10]
  assign tlb__GEN_844 = tlb__T_3583 ? 1'h0 : tlb__GEN_542; // @[TLB.scala 143:19:freechips.rocketchip.system.DefaultRV32Config.fir@183218.10]
  assign tlb__T_3584 = ~tlb__T_3472; // @[TLB.scala 143:13:freechips.rocketchip.system.DefaultRV32Config.fir@183221.10]
  assign tlb__GEN_845 = tlb__T_3584 ? 1'h0 : tlb__GEN_543; // @[TLB.scala 143:19:freechips.rocketchip.system.DefaultRV32Config.fir@183222.10]
  assign tlb__T_3585 = ~tlb__T_3490; // @[TLB.scala 143:13:freechips.rocketchip.system.DefaultRV32Config.fir@183225.10]
  assign tlb__GEN_846 = tlb__T_3585 ? 1'h0 : tlb__GEN_544; // @[TLB.scala 143:19:freechips.rocketchip.system.DefaultRV32Config.fir@183226.10]
  assign tlb__T_3586 = ~tlb__T_3508; // @[TLB.scala 143:13:freechips.rocketchip.system.DefaultRV32Config.fir@183229.10]
  assign tlb__GEN_847 = tlb__T_3586 ? 1'h0 : tlb__GEN_545; // @[TLB.scala 143:19:freechips.rocketchip.system.DefaultRV32Config.fir@183230.10]
  assign tlb__GEN_848 = tlb_io_sfence_bits_rs2 & tlb__GEN_844; // @[TLB.scala 379:40:freechips.rocketchip.system.DefaultRV32Config.fir@183068.8]
  assign tlb__GEN_849 = tlb_io_sfence_bits_rs2 & tlb__GEN_845; // @[TLB.scala 379:40:freechips.rocketchip.system.DefaultRV32Config.fir@183068.8]
  assign tlb__GEN_850 = tlb_io_sfence_bits_rs2 & tlb__GEN_846; // @[TLB.scala 379:40:freechips.rocketchip.system.DefaultRV32Config.fir@183068.8]
  assign tlb__GEN_851 = tlb_io_sfence_bits_rs2 & tlb__GEN_847; // @[TLB.scala 379:40:freechips.rocketchip.system.DefaultRV32Config.fir@183068.8]
  assign tlb__T_3619 = ~tlb__T_800; // @[TLB.scala 143:13:freechips.rocketchip.system.DefaultRV32Config.fir@183298.10]
  assign tlb__GEN_857 = tlb__T_3619 ? 1'h0 : tlb__GEN_458; // @[TLB.scala 143:19:freechips.rocketchip.system.DefaultRV32Config.fir@183299.10]
  assign tlb__GEN_858 = tlb_io_sfence_bits_rs2 & tlb__GEN_857; // @[TLB.scala 379:40:freechips.rocketchip.system.DefaultRV32Config.fir@183260.8]
  assign tlb__T_3652 = ~tlb__T_825; // @[TLB.scala 143:13:freechips.rocketchip.system.DefaultRV32Config.fir@183364.10]
  assign tlb__GEN_861 = tlb__T_3652 ? 1'h0 : tlb__GEN_462; // @[TLB.scala 143:19:freechips.rocketchip.system.DefaultRV32Config.fir@183365.10]
  assign tlb__GEN_862 = tlb_io_sfence_bits_rs2 & tlb__GEN_861; // @[TLB.scala 379:40:freechips.rocketchip.system.DefaultRV32Config.fir@183326.8]
  assign tlb__T_3685 = ~tlb__T_850; // @[TLB.scala 143:13:freechips.rocketchip.system.DefaultRV32Config.fir@183430.10]
  assign tlb__GEN_865 = tlb__T_3685 ? 1'h0 : tlb__GEN_466; // @[TLB.scala 143:19:freechips.rocketchip.system.DefaultRV32Config.fir@183431.10]
  assign tlb__GEN_866 = tlb_io_sfence_bits_rs2 & tlb__GEN_865; // @[TLB.scala 379:40:freechips.rocketchip.system.DefaultRV32Config.fir@183392.8]
  assign tlb__T_3718 = ~tlb__T_875; // @[TLB.scala 143:13:freechips.rocketchip.system.DefaultRV32Config.fir@183496.10]
  assign tlb__GEN_869 = tlb__T_3718 ? 1'h0 : tlb__GEN_470; // @[TLB.scala 143:19:freechips.rocketchip.system.DefaultRV32Config.fir@183497.10]
  assign tlb__GEN_870 = tlb_io_sfence_bits_rs2 & tlb__GEN_869; // @[TLB.scala 379:40:freechips.rocketchip.system.DefaultRV32Config.fir@183458.8]
  assign tlb__T_3751 = ~tlb__T_22; // @[TLB.scala 143:13:freechips.rocketchip.system.DefaultRV32Config.fir@183562.10]
  assign tlb__GEN_873 = tlb__T_3751 ? 1'h0 : tlb__GEN_454; // @[TLB.scala 143:19:freechips.rocketchip.system.DefaultRV32Config.fir@183563.10]
  assign tlb__GEN_874 = tlb_io_sfence_bits_rs2 & tlb__GEN_873; // @[TLB.scala 379:40:freechips.rocketchip.system.DefaultRV32Config.fir@183524.8]
  assign tlb__T_3753 = tlb_multipleHits | tlb_reset; // @[TLB.scala 383:24:freechips.rocketchip.system.DefaultRV32Config.fir@183572.4]
  assign tlb_io_req_ready = tlb_state == 2'h0; // @[TLB.scala 332:16:freechips.rocketchip.system.DefaultRV32Config.fir@180255.4]
  assign tlb_io_resp_miss = tlb__T_2215 | tlb_multipleHits; // @[TLB.scala 345:16:freechips.rocketchip.system.DefaultRV32Config.fir@180299.4]
  assign tlb_io_resp_paddr = {tlb__T_937,tlb__T_34}; // @[TLB.scala 346:17:freechips.rocketchip.system.DefaultRV32Config.fir@180302.4]
  assign tlb_io_resp_pf_ld = |tlb__T_2187; // @[TLB.scala 333:17:freechips.rocketchip.system.DefaultRV32Config.fir@180260.4]
  assign tlb_io_resp_pf_st = |tlb__T_2191; // @[TLB.scala 334:17:freechips.rocketchip.system.DefaultRV32Config.fir@180265.4]
  assign tlb_io_resp_ae_ld = |tlb__T_2197; // @[TLB.scala 336:17:freechips.rocketchip.system.DefaultRV32Config.fir@180272.4]
  assign tlb_io_resp_ae_st = |tlb__T_2199; // @[TLB.scala 337:17:freechips.rocketchip.system.DefaultRV32Config.fir@180275.4]
  assign tlb_io_resp_ma_ld = |tlb__T_2204; // @[TLB.scala 339:17:freechips.rocketchip.system.DefaultRV32Config.fir@180282.4]
  assign tlb_io_resp_ma_st = |tlb__T_2206; // @[TLB.scala 340:17:freechips.rocketchip.system.DefaultRV32Config.fir@180285.4]
  assign tlb_io_resp_cacheable = |tlb__T_2208; // @[TLB.scala 342:21:freechips.rocketchip.system.DefaultRV32Config.fir@180289.4]
  assign tlb_io_ptw_req_valid = tlb_state == 2'h1; // @[TLB.scala 348:20:freechips.rocketchip.system.DefaultRV32Config.fir@180304.4]
  assign tlb_io_ptw_req_bits_bits_addr = tlb_r_refill_tag; // @[TLB.scala 350:29:freechips.rocketchip.system.DefaultRV32Config.fir@180307.4]
  assign tlb_OptimizationBarrier_io_x_ppn = tlb_special_entry_data_0[34:15]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@176911.4]
  assign tlb_OptimizationBarrier_io_x_u = tlb_special_entry_data_0[14]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@176911.4]
  assign tlb_OptimizationBarrier_io_x_ae = tlb_special_entry_data_0[12]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@176911.4]
  assign tlb_OptimizationBarrier_io_x_sw = tlb_special_entry_data_0[11]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@176911.4]
  assign tlb_OptimizationBarrier_io_x_sx = tlb_special_entry_data_0[10]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@176911.4]
  assign tlb_OptimizationBarrier_io_x_sr = tlb_special_entry_data_0[9]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@176911.4]
  assign tlb_OptimizationBarrier_io_x_pw = tlb_special_entry_data_0[8]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@176911.4]
  assign tlb_OptimizationBarrier_io_x_px = tlb_special_entry_data_0[7]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@176911.4]
  assign tlb_OptimizationBarrier_io_x_pr = tlb_special_entry_data_0[6]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@176911.4]
  assign tlb_OptimizationBarrier_io_x_ppp = tlb_special_entry_data_0[5]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@176911.4]
  assign tlb_OptimizationBarrier_io_x_pal = tlb_special_entry_data_0[4]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@176911.4]
  assign tlb_OptimizationBarrier_io_x_paa = tlb_special_entry_data_0[3]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@176911.4]
  assign tlb_OptimizationBarrier_io_x_eff = tlb_special_entry_data_0[2]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@176911.4]
  assign tlb_OptimizationBarrier_io_x_c = tlb_special_entry_data_0[1]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@176911.4]
  assign tlb_pmp_io_prv = tlb_mpu_priv[1:0]; // @[TLB.scala 194:14:freechips.rocketchip.system.DefaultRV32Config.fir@176942.4]
  assign tlb_pmp_io_pmp_0_cfg_l = tlb_io_ptw_pmp_0_cfg_l; // @[TLB.scala 193:14:freechips.rocketchip.system.DefaultRV32Config.fir@176934.4]
  assign tlb_pmp_io_pmp_0_cfg_a = tlb_io_ptw_pmp_0_cfg_a; // @[TLB.scala 193:14:freechips.rocketchip.system.DefaultRV32Config.fir@176934.4]
  assign tlb_pmp_io_pmp_0_cfg_x = tlb_io_ptw_pmp_0_cfg_x; // @[TLB.scala 193:14:freechips.rocketchip.system.DefaultRV32Config.fir@176934.4]
  assign tlb_pmp_io_pmp_0_cfg_w = tlb_io_ptw_pmp_0_cfg_w; // @[TLB.scala 193:14:freechips.rocketchip.system.DefaultRV32Config.fir@176934.4]
  assign tlb_pmp_io_pmp_0_cfg_r = tlb_io_ptw_pmp_0_cfg_r; // @[TLB.scala 193:14:freechips.rocketchip.system.DefaultRV32Config.fir@176934.4]
  assign tlb_pmp_io_pmp_0_addr = tlb_io_ptw_pmp_0_addr; // @[TLB.scala 193:14:freechips.rocketchip.system.DefaultRV32Config.fir@176934.4]
  assign tlb_pmp_io_pmp_0_mask = tlb_io_ptw_pmp_0_mask; // @[TLB.scala 193:14:freechips.rocketchip.system.DefaultRV32Config.fir@176934.4]
  assign tlb_pmp_io_pmp_1_cfg_l = tlb_io_ptw_pmp_1_cfg_l; // @[TLB.scala 193:14:freechips.rocketchip.system.DefaultRV32Config.fir@176935.4]
  assign tlb_pmp_io_pmp_1_cfg_a = tlb_io_ptw_pmp_1_cfg_a; // @[TLB.scala 193:14:freechips.rocketchip.system.DefaultRV32Config.fir@176935.4]
  assign tlb_pmp_io_pmp_1_cfg_x = tlb_io_ptw_pmp_1_cfg_x; // @[TLB.scala 193:14:freechips.rocketchip.system.DefaultRV32Config.fir@176935.4]
  assign tlb_pmp_io_pmp_1_cfg_w = tlb_io_ptw_pmp_1_cfg_w; // @[TLB.scala 193:14:freechips.rocketchip.system.DefaultRV32Config.fir@176935.4]
  assign tlb_pmp_io_pmp_1_cfg_r = tlb_io_ptw_pmp_1_cfg_r; // @[TLB.scala 193:14:freechips.rocketchip.system.DefaultRV32Config.fir@176935.4]
  assign tlb_pmp_io_pmp_1_addr = tlb_io_ptw_pmp_1_addr; // @[TLB.scala 193:14:freechips.rocketchip.system.DefaultRV32Config.fir@176935.4]
  assign tlb_pmp_io_pmp_1_mask = tlb_io_ptw_pmp_1_mask; // @[TLB.scala 193:14:freechips.rocketchip.system.DefaultRV32Config.fir@176935.4]
  assign tlb_pmp_io_pmp_2_cfg_l = tlb_io_ptw_pmp_2_cfg_l; // @[TLB.scala 193:14:freechips.rocketchip.system.DefaultRV32Config.fir@176936.4]
  assign tlb_pmp_io_pmp_2_cfg_a = tlb_io_ptw_pmp_2_cfg_a; // @[TLB.scala 193:14:freechips.rocketchip.system.DefaultRV32Config.fir@176936.4]
  assign tlb_pmp_io_pmp_2_cfg_x = tlb_io_ptw_pmp_2_cfg_x; // @[TLB.scala 193:14:freechips.rocketchip.system.DefaultRV32Config.fir@176936.4]
  assign tlb_pmp_io_pmp_2_cfg_w = tlb_io_ptw_pmp_2_cfg_w; // @[TLB.scala 193:14:freechips.rocketchip.system.DefaultRV32Config.fir@176936.4]
  assign tlb_pmp_io_pmp_2_cfg_r = tlb_io_ptw_pmp_2_cfg_r; // @[TLB.scala 193:14:freechips.rocketchip.system.DefaultRV32Config.fir@176936.4]
  assign tlb_pmp_io_pmp_2_addr = tlb_io_ptw_pmp_2_addr; // @[TLB.scala 193:14:freechips.rocketchip.system.DefaultRV32Config.fir@176936.4]
  assign tlb_pmp_io_pmp_2_mask = tlb_io_ptw_pmp_2_mask; // @[TLB.scala 193:14:freechips.rocketchip.system.DefaultRV32Config.fir@176936.4]
  assign tlb_pmp_io_pmp_3_cfg_l = tlb_io_ptw_pmp_3_cfg_l; // @[TLB.scala 193:14:freechips.rocketchip.system.DefaultRV32Config.fir@176937.4]
  assign tlb_pmp_io_pmp_3_cfg_a = tlb_io_ptw_pmp_3_cfg_a; // @[TLB.scala 193:14:freechips.rocketchip.system.DefaultRV32Config.fir@176937.4]
  assign tlb_pmp_io_pmp_3_cfg_x = tlb_io_ptw_pmp_3_cfg_x; // @[TLB.scala 193:14:freechips.rocketchip.system.DefaultRV32Config.fir@176937.4]
  assign tlb_pmp_io_pmp_3_cfg_w = tlb_io_ptw_pmp_3_cfg_w; // @[TLB.scala 193:14:freechips.rocketchip.system.DefaultRV32Config.fir@176937.4]
  assign tlb_pmp_io_pmp_3_cfg_r = tlb_io_ptw_pmp_3_cfg_r; // @[TLB.scala 193:14:freechips.rocketchip.system.DefaultRV32Config.fir@176937.4]
  assign tlb_pmp_io_pmp_3_addr = tlb_io_ptw_pmp_3_addr; // @[TLB.scala 193:14:freechips.rocketchip.system.DefaultRV32Config.fir@176937.4]
  assign tlb_pmp_io_pmp_3_mask = tlb_io_ptw_pmp_3_mask; // @[TLB.scala 193:14:freechips.rocketchip.system.DefaultRV32Config.fir@176937.4]
  assign tlb_pmp_io_pmp_4_cfg_l = tlb_io_ptw_pmp_4_cfg_l; // @[TLB.scala 193:14:freechips.rocketchip.system.DefaultRV32Config.fir@176938.4]
  assign tlb_pmp_io_pmp_4_cfg_a = tlb_io_ptw_pmp_4_cfg_a; // @[TLB.scala 193:14:freechips.rocketchip.system.DefaultRV32Config.fir@176938.4]
  assign tlb_pmp_io_pmp_4_cfg_x = tlb_io_ptw_pmp_4_cfg_x; // @[TLB.scala 193:14:freechips.rocketchip.system.DefaultRV32Config.fir@176938.4]
  assign tlb_pmp_io_pmp_4_cfg_w = tlb_io_ptw_pmp_4_cfg_w; // @[TLB.scala 193:14:freechips.rocketchip.system.DefaultRV32Config.fir@176938.4]
  assign tlb_pmp_io_pmp_4_cfg_r = tlb_io_ptw_pmp_4_cfg_r; // @[TLB.scala 193:14:freechips.rocketchip.system.DefaultRV32Config.fir@176938.4]
  assign tlb_pmp_io_pmp_4_addr = tlb_io_ptw_pmp_4_addr; // @[TLB.scala 193:14:freechips.rocketchip.system.DefaultRV32Config.fir@176938.4]
  assign tlb_pmp_io_pmp_4_mask = tlb_io_ptw_pmp_4_mask; // @[TLB.scala 193:14:freechips.rocketchip.system.DefaultRV32Config.fir@176938.4]
  assign tlb_pmp_io_pmp_5_cfg_l = tlb_io_ptw_pmp_5_cfg_l; // @[TLB.scala 193:14:freechips.rocketchip.system.DefaultRV32Config.fir@176939.4]
  assign tlb_pmp_io_pmp_5_cfg_a = tlb_io_ptw_pmp_5_cfg_a; // @[TLB.scala 193:14:freechips.rocketchip.system.DefaultRV32Config.fir@176939.4]
  assign tlb_pmp_io_pmp_5_cfg_x = tlb_io_ptw_pmp_5_cfg_x; // @[TLB.scala 193:14:freechips.rocketchip.system.DefaultRV32Config.fir@176939.4]
  assign tlb_pmp_io_pmp_5_cfg_w = tlb_io_ptw_pmp_5_cfg_w; // @[TLB.scala 193:14:freechips.rocketchip.system.DefaultRV32Config.fir@176939.4]
  assign tlb_pmp_io_pmp_5_cfg_r = tlb_io_ptw_pmp_5_cfg_r; // @[TLB.scala 193:14:freechips.rocketchip.system.DefaultRV32Config.fir@176939.4]
  assign tlb_pmp_io_pmp_5_addr = tlb_io_ptw_pmp_5_addr; // @[TLB.scala 193:14:freechips.rocketchip.system.DefaultRV32Config.fir@176939.4]
  assign tlb_pmp_io_pmp_5_mask = tlb_io_ptw_pmp_5_mask; // @[TLB.scala 193:14:freechips.rocketchip.system.DefaultRV32Config.fir@176939.4]
  assign tlb_pmp_io_pmp_6_cfg_l = tlb_io_ptw_pmp_6_cfg_l; // @[TLB.scala 193:14:freechips.rocketchip.system.DefaultRV32Config.fir@176940.4]
  assign tlb_pmp_io_pmp_6_cfg_a = tlb_io_ptw_pmp_6_cfg_a; // @[TLB.scala 193:14:freechips.rocketchip.system.DefaultRV32Config.fir@176940.4]
  assign tlb_pmp_io_pmp_6_cfg_x = tlb_io_ptw_pmp_6_cfg_x; // @[TLB.scala 193:14:freechips.rocketchip.system.DefaultRV32Config.fir@176940.4]
  assign tlb_pmp_io_pmp_6_cfg_w = tlb_io_ptw_pmp_6_cfg_w; // @[TLB.scala 193:14:freechips.rocketchip.system.DefaultRV32Config.fir@176940.4]
  assign tlb_pmp_io_pmp_6_cfg_r = tlb_io_ptw_pmp_6_cfg_r; // @[TLB.scala 193:14:freechips.rocketchip.system.DefaultRV32Config.fir@176940.4]
  assign tlb_pmp_io_pmp_6_addr = tlb_io_ptw_pmp_6_addr; // @[TLB.scala 193:14:freechips.rocketchip.system.DefaultRV32Config.fir@176940.4]
  assign tlb_pmp_io_pmp_6_mask = tlb_io_ptw_pmp_6_mask; // @[TLB.scala 193:14:freechips.rocketchip.system.DefaultRV32Config.fir@176940.4]
  assign tlb_pmp_io_pmp_7_cfg_l = tlb_io_ptw_pmp_7_cfg_l; // @[TLB.scala 193:14:freechips.rocketchip.system.DefaultRV32Config.fir@176941.4]
  assign tlb_pmp_io_pmp_7_cfg_a = tlb_io_ptw_pmp_7_cfg_a; // @[TLB.scala 193:14:freechips.rocketchip.system.DefaultRV32Config.fir@176941.4]
  assign tlb_pmp_io_pmp_7_cfg_x = tlb_io_ptw_pmp_7_cfg_x; // @[TLB.scala 193:14:freechips.rocketchip.system.DefaultRV32Config.fir@176941.4]
  assign tlb_pmp_io_pmp_7_cfg_w = tlb_io_ptw_pmp_7_cfg_w; // @[TLB.scala 193:14:freechips.rocketchip.system.DefaultRV32Config.fir@176941.4]
  assign tlb_pmp_io_pmp_7_cfg_r = tlb_io_ptw_pmp_7_cfg_r; // @[TLB.scala 193:14:freechips.rocketchip.system.DefaultRV32Config.fir@176941.4]
  assign tlb_pmp_io_pmp_7_addr = tlb_io_ptw_pmp_7_addr; // @[TLB.scala 193:14:freechips.rocketchip.system.DefaultRV32Config.fir@176941.4]
  assign tlb_pmp_io_pmp_7_mask = tlb_io_ptw_pmp_7_mask; // @[TLB.scala 193:14:freechips.rocketchip.system.DefaultRV32Config.fir@176941.4]
  assign tlb_pmp_io_addr = {tlb_mpu_ppn,tlb__T_34}; // @[TLB.scala 191:15:freechips.rocketchip.system.DefaultRV32Config.fir@176932.4]
  assign tlb_OptimizationBarrier_1_io_x_ppn = tlb__GEN_35[34:15]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@177633.4]
  assign tlb_OptimizationBarrier_1_io_x_u = tlb__GEN_35[14]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@177633.4]
  assign tlb_OptimizationBarrier_1_io_x_ae = tlb__GEN_35[12]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@177633.4]
  assign tlb_OptimizationBarrier_1_io_x_sw = tlb__GEN_35[11]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@177633.4]
  assign tlb_OptimizationBarrier_1_io_x_sx = tlb__GEN_35[10]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@177633.4]
  assign tlb_OptimizationBarrier_1_io_x_sr = tlb__GEN_35[9]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@177633.4]
  assign tlb_OptimizationBarrier_1_io_x_pw = tlb__GEN_35[8]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@177633.4]
  assign tlb_OptimizationBarrier_1_io_x_px = tlb__GEN_35[7]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@177633.4]
  assign tlb_OptimizationBarrier_1_io_x_pr = tlb__GEN_35[6]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@177633.4]
  assign tlb_OptimizationBarrier_1_io_x_ppp = tlb__GEN_35[5]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@177633.4]
  assign tlb_OptimizationBarrier_1_io_x_pal = tlb__GEN_35[4]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@177633.4]
  assign tlb_OptimizationBarrier_1_io_x_paa = tlb__GEN_35[3]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@177633.4]
  assign tlb_OptimizationBarrier_1_io_x_eff = tlb__GEN_35[2]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@177633.4]
  assign tlb_OptimizationBarrier_1_io_x_c = tlb__GEN_35[1]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@177633.4]
  assign tlb_OptimizationBarrier_2_io_x_ppn = tlb__GEN_39[34:15]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@177676.4]
  assign tlb_OptimizationBarrier_2_io_x_u = tlb__GEN_39[14]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@177676.4]
  assign tlb_OptimizationBarrier_2_io_x_ae = tlb__GEN_39[12]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@177676.4]
  assign tlb_OptimizationBarrier_2_io_x_sw = tlb__GEN_39[11]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@177676.4]
  assign tlb_OptimizationBarrier_2_io_x_sx = tlb__GEN_39[10]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@177676.4]
  assign tlb_OptimizationBarrier_2_io_x_sr = tlb__GEN_39[9]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@177676.4]
  assign tlb_OptimizationBarrier_2_io_x_pw = tlb__GEN_39[8]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@177676.4]
  assign tlb_OptimizationBarrier_2_io_x_px = tlb__GEN_39[7]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@177676.4]
  assign tlb_OptimizationBarrier_2_io_x_pr = tlb__GEN_39[6]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@177676.4]
  assign tlb_OptimizationBarrier_2_io_x_ppp = tlb__GEN_39[5]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@177676.4]
  assign tlb_OptimizationBarrier_2_io_x_pal = tlb__GEN_39[4]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@177676.4]
  assign tlb_OptimizationBarrier_2_io_x_paa = tlb__GEN_39[3]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@177676.4]
  assign tlb_OptimizationBarrier_2_io_x_eff = tlb__GEN_39[2]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@177676.4]
  assign tlb_OptimizationBarrier_2_io_x_c = tlb__GEN_39[1]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@177676.4]
  assign tlb_OptimizationBarrier_3_io_x_ppn = tlb__GEN_43[34:15]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@177719.4]
  assign tlb_OptimizationBarrier_3_io_x_u = tlb__GEN_43[14]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@177719.4]
  assign tlb_OptimizationBarrier_3_io_x_ae = tlb__GEN_43[12]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@177719.4]
  assign tlb_OptimizationBarrier_3_io_x_sw = tlb__GEN_43[11]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@177719.4]
  assign tlb_OptimizationBarrier_3_io_x_sx = tlb__GEN_43[10]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@177719.4]
  assign tlb_OptimizationBarrier_3_io_x_sr = tlb__GEN_43[9]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@177719.4]
  assign tlb_OptimizationBarrier_3_io_x_pw = tlb__GEN_43[8]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@177719.4]
  assign tlb_OptimizationBarrier_3_io_x_px = tlb__GEN_43[7]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@177719.4]
  assign tlb_OptimizationBarrier_3_io_x_pr = tlb__GEN_43[6]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@177719.4]
  assign tlb_OptimizationBarrier_3_io_x_ppp = tlb__GEN_43[5]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@177719.4]
  assign tlb_OptimizationBarrier_3_io_x_pal = tlb__GEN_43[4]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@177719.4]
  assign tlb_OptimizationBarrier_3_io_x_paa = tlb__GEN_43[3]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@177719.4]
  assign tlb_OptimizationBarrier_3_io_x_eff = tlb__GEN_43[2]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@177719.4]
  assign tlb_OptimizationBarrier_3_io_x_c = tlb__GEN_43[1]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@177719.4]
  assign tlb_OptimizationBarrier_4_io_x_ppn = tlb__GEN_47[34:15]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@177762.4]
  assign tlb_OptimizationBarrier_4_io_x_u = tlb__GEN_47[14]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@177762.4]
  assign tlb_OptimizationBarrier_4_io_x_ae = tlb__GEN_47[12]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@177762.4]
  assign tlb_OptimizationBarrier_4_io_x_sw = tlb__GEN_47[11]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@177762.4]
  assign tlb_OptimizationBarrier_4_io_x_sx = tlb__GEN_47[10]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@177762.4]
  assign tlb_OptimizationBarrier_4_io_x_sr = tlb__GEN_47[9]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@177762.4]
  assign tlb_OptimizationBarrier_4_io_x_pw = tlb__GEN_47[8]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@177762.4]
  assign tlb_OptimizationBarrier_4_io_x_px = tlb__GEN_47[7]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@177762.4]
  assign tlb_OptimizationBarrier_4_io_x_pr = tlb__GEN_47[6]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@177762.4]
  assign tlb_OptimizationBarrier_4_io_x_ppp = tlb__GEN_47[5]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@177762.4]
  assign tlb_OptimizationBarrier_4_io_x_pal = tlb__GEN_47[4]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@177762.4]
  assign tlb_OptimizationBarrier_4_io_x_paa = tlb__GEN_47[3]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@177762.4]
  assign tlb_OptimizationBarrier_4_io_x_eff = tlb__GEN_47[2]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@177762.4]
  assign tlb_OptimizationBarrier_4_io_x_c = tlb__GEN_47[1]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@177762.4]
  assign tlb_OptimizationBarrier_5_io_x_ppn = tlb__GEN_51[34:15]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@177805.4]
  assign tlb_OptimizationBarrier_5_io_x_u = tlb__GEN_51[14]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@177805.4]
  assign tlb_OptimizationBarrier_5_io_x_ae = tlb__GEN_51[12]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@177805.4]
  assign tlb_OptimizationBarrier_5_io_x_sw = tlb__GEN_51[11]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@177805.4]
  assign tlb_OptimizationBarrier_5_io_x_sx = tlb__GEN_51[10]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@177805.4]
  assign tlb_OptimizationBarrier_5_io_x_sr = tlb__GEN_51[9]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@177805.4]
  assign tlb_OptimizationBarrier_5_io_x_pw = tlb__GEN_51[8]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@177805.4]
  assign tlb_OptimizationBarrier_5_io_x_px = tlb__GEN_51[7]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@177805.4]
  assign tlb_OptimizationBarrier_5_io_x_pr = tlb__GEN_51[6]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@177805.4]
  assign tlb_OptimizationBarrier_5_io_x_ppp = tlb__GEN_51[5]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@177805.4]
  assign tlb_OptimizationBarrier_5_io_x_pal = tlb__GEN_51[4]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@177805.4]
  assign tlb_OptimizationBarrier_5_io_x_paa = tlb__GEN_51[3]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@177805.4]
  assign tlb_OptimizationBarrier_5_io_x_eff = tlb__GEN_51[2]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@177805.4]
  assign tlb_OptimizationBarrier_5_io_x_c = tlb__GEN_51[1]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@177805.4]
  assign tlb_OptimizationBarrier_6_io_x_ppn = tlb__GEN_55[34:15]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@177848.4]
  assign tlb_OptimizationBarrier_6_io_x_u = tlb__GEN_55[14]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@177848.4]
  assign tlb_OptimizationBarrier_6_io_x_ae = tlb__GEN_55[12]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@177848.4]
  assign tlb_OptimizationBarrier_6_io_x_sw = tlb__GEN_55[11]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@177848.4]
  assign tlb_OptimizationBarrier_6_io_x_sx = tlb__GEN_55[10]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@177848.4]
  assign tlb_OptimizationBarrier_6_io_x_sr = tlb__GEN_55[9]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@177848.4]
  assign tlb_OptimizationBarrier_6_io_x_pw = tlb__GEN_55[8]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@177848.4]
  assign tlb_OptimizationBarrier_6_io_x_px = tlb__GEN_55[7]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@177848.4]
  assign tlb_OptimizationBarrier_6_io_x_pr = tlb__GEN_55[6]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@177848.4]
  assign tlb_OptimizationBarrier_6_io_x_ppp = tlb__GEN_55[5]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@177848.4]
  assign tlb_OptimizationBarrier_6_io_x_pal = tlb__GEN_55[4]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@177848.4]
  assign tlb_OptimizationBarrier_6_io_x_paa = tlb__GEN_55[3]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@177848.4]
  assign tlb_OptimizationBarrier_6_io_x_eff = tlb__GEN_55[2]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@177848.4]
  assign tlb_OptimizationBarrier_6_io_x_c = tlb__GEN_55[1]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@177848.4]
  assign tlb_OptimizationBarrier_7_io_x_ppn = tlb__GEN_59[34:15]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@177891.4]
  assign tlb_OptimizationBarrier_7_io_x_u = tlb__GEN_59[14]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@177891.4]
  assign tlb_OptimizationBarrier_7_io_x_ae = tlb__GEN_59[12]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@177891.4]
  assign tlb_OptimizationBarrier_7_io_x_sw = tlb__GEN_59[11]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@177891.4]
  assign tlb_OptimizationBarrier_7_io_x_sx = tlb__GEN_59[10]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@177891.4]
  assign tlb_OptimizationBarrier_7_io_x_sr = tlb__GEN_59[9]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@177891.4]
  assign tlb_OptimizationBarrier_7_io_x_pw = tlb__GEN_59[8]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@177891.4]
  assign tlb_OptimizationBarrier_7_io_x_px = tlb__GEN_59[7]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@177891.4]
  assign tlb_OptimizationBarrier_7_io_x_pr = tlb__GEN_59[6]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@177891.4]
  assign tlb_OptimizationBarrier_7_io_x_ppp = tlb__GEN_59[5]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@177891.4]
  assign tlb_OptimizationBarrier_7_io_x_pal = tlb__GEN_59[4]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@177891.4]
  assign tlb_OptimizationBarrier_7_io_x_paa = tlb__GEN_59[3]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@177891.4]
  assign tlb_OptimizationBarrier_7_io_x_eff = tlb__GEN_59[2]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@177891.4]
  assign tlb_OptimizationBarrier_7_io_x_c = tlb__GEN_59[1]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@177891.4]
  assign tlb_OptimizationBarrier_8_io_x_ppn = tlb__GEN_63[34:15]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@177934.4]
  assign tlb_OptimizationBarrier_8_io_x_u = tlb__GEN_63[14]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@177934.4]
  assign tlb_OptimizationBarrier_8_io_x_ae = tlb__GEN_63[12]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@177934.4]
  assign tlb_OptimizationBarrier_8_io_x_sw = tlb__GEN_63[11]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@177934.4]
  assign tlb_OptimizationBarrier_8_io_x_sx = tlb__GEN_63[10]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@177934.4]
  assign tlb_OptimizationBarrier_8_io_x_sr = tlb__GEN_63[9]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@177934.4]
  assign tlb_OptimizationBarrier_8_io_x_pw = tlb__GEN_63[8]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@177934.4]
  assign tlb_OptimizationBarrier_8_io_x_px = tlb__GEN_63[7]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@177934.4]
  assign tlb_OptimizationBarrier_8_io_x_pr = tlb__GEN_63[6]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@177934.4]
  assign tlb_OptimizationBarrier_8_io_x_ppp = tlb__GEN_63[5]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@177934.4]
  assign tlb_OptimizationBarrier_8_io_x_pal = tlb__GEN_63[4]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@177934.4]
  assign tlb_OptimizationBarrier_8_io_x_paa = tlb__GEN_63[3]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@177934.4]
  assign tlb_OptimizationBarrier_8_io_x_eff = tlb__GEN_63[2]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@177934.4]
  assign tlb_OptimizationBarrier_8_io_x_c = tlb__GEN_63[1]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@177934.4]
  assign tlb_OptimizationBarrier_9_io_x_ppn = tlb_superpage_entries_0_data_0[34:15]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@177976.4]
  assign tlb_OptimizationBarrier_9_io_x_u = tlb_superpage_entries_0_data_0[14]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@177976.4]
  assign tlb_OptimizationBarrier_9_io_x_ae = tlb_superpage_entries_0_data_0[12]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@177976.4]
  assign tlb_OptimizationBarrier_9_io_x_sw = tlb_superpage_entries_0_data_0[11]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@177976.4]
  assign tlb_OptimizationBarrier_9_io_x_sx = tlb_superpage_entries_0_data_0[10]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@177976.4]
  assign tlb_OptimizationBarrier_9_io_x_sr = tlb_superpage_entries_0_data_0[9]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@177976.4]
  assign tlb_OptimizationBarrier_9_io_x_pw = tlb_superpage_entries_0_data_0[8]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@177976.4]
  assign tlb_OptimizationBarrier_9_io_x_px = tlb_superpage_entries_0_data_0[7]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@177976.4]
  assign tlb_OptimizationBarrier_9_io_x_pr = tlb_superpage_entries_0_data_0[6]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@177976.4]
  assign tlb_OptimizationBarrier_9_io_x_ppp = tlb_superpage_entries_0_data_0[5]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@177976.4]
  assign tlb_OptimizationBarrier_9_io_x_pal = tlb_superpage_entries_0_data_0[4]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@177976.4]
  assign tlb_OptimizationBarrier_9_io_x_paa = tlb_superpage_entries_0_data_0[3]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@177976.4]
  assign tlb_OptimizationBarrier_9_io_x_eff = tlb_superpage_entries_0_data_0[2]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@177976.4]
  assign tlb_OptimizationBarrier_9_io_x_c = tlb_superpage_entries_0_data_0[1]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@177976.4]
  assign tlb_OptimizationBarrier_10_io_x_ppn = tlb_superpage_entries_1_data_0[34:15]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@178025.4]
  assign tlb_OptimizationBarrier_10_io_x_u = tlb_superpage_entries_1_data_0[14]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@178025.4]
  assign tlb_OptimizationBarrier_10_io_x_ae = tlb_superpage_entries_1_data_0[12]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@178025.4]
  assign tlb_OptimizationBarrier_10_io_x_sw = tlb_superpage_entries_1_data_0[11]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@178025.4]
  assign tlb_OptimizationBarrier_10_io_x_sx = tlb_superpage_entries_1_data_0[10]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@178025.4]
  assign tlb_OptimizationBarrier_10_io_x_sr = tlb_superpage_entries_1_data_0[9]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@178025.4]
  assign tlb_OptimizationBarrier_10_io_x_pw = tlb_superpage_entries_1_data_0[8]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@178025.4]
  assign tlb_OptimizationBarrier_10_io_x_px = tlb_superpage_entries_1_data_0[7]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@178025.4]
  assign tlb_OptimizationBarrier_10_io_x_pr = tlb_superpage_entries_1_data_0[6]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@178025.4]
  assign tlb_OptimizationBarrier_10_io_x_ppp = tlb_superpage_entries_1_data_0[5]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@178025.4]
  assign tlb_OptimizationBarrier_10_io_x_pal = tlb_superpage_entries_1_data_0[4]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@178025.4]
  assign tlb_OptimizationBarrier_10_io_x_paa = tlb_superpage_entries_1_data_0[3]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@178025.4]
  assign tlb_OptimizationBarrier_10_io_x_eff = tlb_superpage_entries_1_data_0[2]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@178025.4]
  assign tlb_OptimizationBarrier_10_io_x_c = tlb_superpage_entries_1_data_0[1]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@178025.4]
  assign tlb_OptimizationBarrier_11_io_x_ppn = tlb_superpage_entries_2_data_0[34:15]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@178074.4]
  assign tlb_OptimizationBarrier_11_io_x_u = tlb_superpage_entries_2_data_0[14]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@178074.4]
  assign tlb_OptimizationBarrier_11_io_x_ae = tlb_superpage_entries_2_data_0[12]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@178074.4]
  assign tlb_OptimizationBarrier_11_io_x_sw = tlb_superpage_entries_2_data_0[11]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@178074.4]
  assign tlb_OptimizationBarrier_11_io_x_sx = tlb_superpage_entries_2_data_0[10]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@178074.4]
  assign tlb_OptimizationBarrier_11_io_x_sr = tlb_superpage_entries_2_data_0[9]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@178074.4]
  assign tlb_OptimizationBarrier_11_io_x_pw = tlb_superpage_entries_2_data_0[8]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@178074.4]
  assign tlb_OptimizationBarrier_11_io_x_px = tlb_superpage_entries_2_data_0[7]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@178074.4]
  assign tlb_OptimizationBarrier_11_io_x_pr = tlb_superpage_entries_2_data_0[6]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@178074.4]
  assign tlb_OptimizationBarrier_11_io_x_ppp = tlb_superpage_entries_2_data_0[5]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@178074.4]
  assign tlb_OptimizationBarrier_11_io_x_pal = tlb_superpage_entries_2_data_0[4]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@178074.4]
  assign tlb_OptimizationBarrier_11_io_x_paa = tlb_superpage_entries_2_data_0[3]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@178074.4]
  assign tlb_OptimizationBarrier_11_io_x_eff = tlb_superpage_entries_2_data_0[2]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@178074.4]
  assign tlb_OptimizationBarrier_11_io_x_c = tlb_superpage_entries_2_data_0[1]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@178074.4]
  assign tlb_OptimizationBarrier_12_io_x_ppn = tlb_superpage_entries_3_data_0[34:15]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@178123.4]
  assign tlb_OptimizationBarrier_12_io_x_u = tlb_superpage_entries_3_data_0[14]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@178123.4]
  assign tlb_OptimizationBarrier_12_io_x_ae = tlb_superpage_entries_3_data_0[12]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@178123.4]
  assign tlb_OptimizationBarrier_12_io_x_sw = tlb_superpage_entries_3_data_0[11]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@178123.4]
  assign tlb_OptimizationBarrier_12_io_x_sx = tlb_superpage_entries_3_data_0[10]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@178123.4]
  assign tlb_OptimizationBarrier_12_io_x_sr = tlb_superpage_entries_3_data_0[9]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@178123.4]
  assign tlb_OptimizationBarrier_12_io_x_pw = tlb_superpage_entries_3_data_0[8]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@178123.4]
  assign tlb_OptimizationBarrier_12_io_x_px = tlb_superpage_entries_3_data_0[7]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@178123.4]
  assign tlb_OptimizationBarrier_12_io_x_pr = tlb_superpage_entries_3_data_0[6]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@178123.4]
  assign tlb_OptimizationBarrier_12_io_x_ppp = tlb_superpage_entries_3_data_0[5]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@178123.4]
  assign tlb_OptimizationBarrier_12_io_x_pal = tlb_superpage_entries_3_data_0[4]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@178123.4]
  assign tlb_OptimizationBarrier_12_io_x_paa = tlb_superpage_entries_3_data_0[3]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@178123.4]
  assign tlb_OptimizationBarrier_12_io_x_eff = tlb_superpage_entries_3_data_0[2]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@178123.4]
  assign tlb_OptimizationBarrier_12_io_x_c = tlb_superpage_entries_3_data_0[1]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@178123.4]
  assign tlb_OptimizationBarrier_13_io_x_ppn = tlb_special_entry_data_0[34:15]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@178172.4]
  assign tlb_OptimizationBarrier_13_io_x_u = tlb_special_entry_data_0[14]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@178172.4]
  assign tlb_OptimizationBarrier_13_io_x_ae = tlb_special_entry_data_0[12]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@178172.4]
  assign tlb_OptimizationBarrier_13_io_x_sw = tlb_special_entry_data_0[11]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@178172.4]
  assign tlb_OptimizationBarrier_13_io_x_sx = tlb_special_entry_data_0[10]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@178172.4]
  assign tlb_OptimizationBarrier_13_io_x_sr = tlb_special_entry_data_0[9]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@178172.4]
  assign tlb_OptimizationBarrier_13_io_x_pw = tlb_special_entry_data_0[8]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@178172.4]
  assign tlb_OptimizationBarrier_13_io_x_px = tlb_special_entry_data_0[7]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@178172.4]
  assign tlb_OptimizationBarrier_13_io_x_pr = tlb_special_entry_data_0[6]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@178172.4]
  assign tlb_OptimizationBarrier_13_io_x_ppp = tlb_special_entry_data_0[5]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@178172.4]
  assign tlb_OptimizationBarrier_13_io_x_pal = tlb_special_entry_data_0[4]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@178172.4]
  assign tlb_OptimizationBarrier_13_io_x_paa = tlb_special_entry_data_0[3]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@178172.4]
  assign tlb_OptimizationBarrier_13_io_x_eff = tlb_special_entry_data_0[2]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@178172.4]
  assign tlb_OptimizationBarrier_13_io_x_c = tlb_special_entry_data_0[1]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@178172.4]
  assign tlb_OptimizationBarrier_14_io_x_ppn = tlb__GEN_35[34:15]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@178653.4]
  assign tlb_OptimizationBarrier_14_io_x_u = tlb__GEN_35[14]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@178653.4]
  assign tlb_OptimizationBarrier_14_io_x_ae = tlb__GEN_35[12]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@178653.4]
  assign tlb_OptimizationBarrier_14_io_x_sw = tlb__GEN_35[11]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@178653.4]
  assign tlb_OptimizationBarrier_14_io_x_sx = tlb__GEN_35[10]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@178653.4]
  assign tlb_OptimizationBarrier_14_io_x_sr = tlb__GEN_35[9]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@178653.4]
  assign tlb_OptimizationBarrier_14_io_x_pw = tlb__GEN_35[8]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@178653.4]
  assign tlb_OptimizationBarrier_14_io_x_px = tlb__GEN_35[7]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@178653.4]
  assign tlb_OptimizationBarrier_14_io_x_pr = tlb__GEN_35[6]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@178653.4]
  assign tlb_OptimizationBarrier_14_io_x_ppp = tlb__GEN_35[5]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@178653.4]
  assign tlb_OptimizationBarrier_14_io_x_pal = tlb__GEN_35[4]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@178653.4]
  assign tlb_OptimizationBarrier_14_io_x_paa = tlb__GEN_35[3]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@178653.4]
  assign tlb_OptimizationBarrier_14_io_x_eff = tlb__GEN_35[2]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@178653.4]
  assign tlb_OptimizationBarrier_14_io_x_c = tlb__GEN_35[1]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@178653.4]
  assign tlb_OptimizationBarrier_15_io_x_ppn = tlb__GEN_39[34:15]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@178696.4]
  assign tlb_OptimizationBarrier_15_io_x_u = tlb__GEN_39[14]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@178696.4]
  assign tlb_OptimizationBarrier_15_io_x_ae = tlb__GEN_39[12]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@178696.4]
  assign tlb_OptimizationBarrier_15_io_x_sw = tlb__GEN_39[11]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@178696.4]
  assign tlb_OptimizationBarrier_15_io_x_sx = tlb__GEN_39[10]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@178696.4]
  assign tlb_OptimizationBarrier_15_io_x_sr = tlb__GEN_39[9]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@178696.4]
  assign tlb_OptimizationBarrier_15_io_x_pw = tlb__GEN_39[8]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@178696.4]
  assign tlb_OptimizationBarrier_15_io_x_px = tlb__GEN_39[7]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@178696.4]
  assign tlb_OptimizationBarrier_15_io_x_pr = tlb__GEN_39[6]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@178696.4]
  assign tlb_OptimizationBarrier_15_io_x_ppp = tlb__GEN_39[5]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@178696.4]
  assign tlb_OptimizationBarrier_15_io_x_pal = tlb__GEN_39[4]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@178696.4]
  assign tlb_OptimizationBarrier_15_io_x_paa = tlb__GEN_39[3]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@178696.4]
  assign tlb_OptimizationBarrier_15_io_x_eff = tlb__GEN_39[2]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@178696.4]
  assign tlb_OptimizationBarrier_15_io_x_c = tlb__GEN_39[1]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@178696.4]
  assign tlb_OptimizationBarrier_16_io_x_ppn = tlb__GEN_43[34:15]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@178739.4]
  assign tlb_OptimizationBarrier_16_io_x_u = tlb__GEN_43[14]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@178739.4]
  assign tlb_OptimizationBarrier_16_io_x_ae = tlb__GEN_43[12]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@178739.4]
  assign tlb_OptimizationBarrier_16_io_x_sw = tlb__GEN_43[11]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@178739.4]
  assign tlb_OptimizationBarrier_16_io_x_sx = tlb__GEN_43[10]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@178739.4]
  assign tlb_OptimizationBarrier_16_io_x_sr = tlb__GEN_43[9]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@178739.4]
  assign tlb_OptimizationBarrier_16_io_x_pw = tlb__GEN_43[8]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@178739.4]
  assign tlb_OptimizationBarrier_16_io_x_px = tlb__GEN_43[7]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@178739.4]
  assign tlb_OptimizationBarrier_16_io_x_pr = tlb__GEN_43[6]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@178739.4]
  assign tlb_OptimizationBarrier_16_io_x_ppp = tlb__GEN_43[5]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@178739.4]
  assign tlb_OptimizationBarrier_16_io_x_pal = tlb__GEN_43[4]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@178739.4]
  assign tlb_OptimizationBarrier_16_io_x_paa = tlb__GEN_43[3]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@178739.4]
  assign tlb_OptimizationBarrier_16_io_x_eff = tlb__GEN_43[2]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@178739.4]
  assign tlb_OptimizationBarrier_16_io_x_c = tlb__GEN_43[1]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@178739.4]
  assign tlb_OptimizationBarrier_17_io_x_ppn = tlb__GEN_47[34:15]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@178782.4]
  assign tlb_OptimizationBarrier_17_io_x_u = tlb__GEN_47[14]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@178782.4]
  assign tlb_OptimizationBarrier_17_io_x_ae = tlb__GEN_47[12]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@178782.4]
  assign tlb_OptimizationBarrier_17_io_x_sw = tlb__GEN_47[11]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@178782.4]
  assign tlb_OptimizationBarrier_17_io_x_sx = tlb__GEN_47[10]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@178782.4]
  assign tlb_OptimizationBarrier_17_io_x_sr = tlb__GEN_47[9]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@178782.4]
  assign tlb_OptimizationBarrier_17_io_x_pw = tlb__GEN_47[8]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@178782.4]
  assign tlb_OptimizationBarrier_17_io_x_px = tlb__GEN_47[7]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@178782.4]
  assign tlb_OptimizationBarrier_17_io_x_pr = tlb__GEN_47[6]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@178782.4]
  assign tlb_OptimizationBarrier_17_io_x_ppp = tlb__GEN_47[5]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@178782.4]
  assign tlb_OptimizationBarrier_17_io_x_pal = tlb__GEN_47[4]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@178782.4]
  assign tlb_OptimizationBarrier_17_io_x_paa = tlb__GEN_47[3]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@178782.4]
  assign tlb_OptimizationBarrier_17_io_x_eff = tlb__GEN_47[2]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@178782.4]
  assign tlb_OptimizationBarrier_17_io_x_c = tlb__GEN_47[1]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@178782.4]
  assign tlb_OptimizationBarrier_18_io_x_ppn = tlb__GEN_51[34:15]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@178825.4]
  assign tlb_OptimizationBarrier_18_io_x_u = tlb__GEN_51[14]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@178825.4]
  assign tlb_OptimizationBarrier_18_io_x_ae = tlb__GEN_51[12]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@178825.4]
  assign tlb_OptimizationBarrier_18_io_x_sw = tlb__GEN_51[11]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@178825.4]
  assign tlb_OptimizationBarrier_18_io_x_sx = tlb__GEN_51[10]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@178825.4]
  assign tlb_OptimizationBarrier_18_io_x_sr = tlb__GEN_51[9]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@178825.4]
  assign tlb_OptimizationBarrier_18_io_x_pw = tlb__GEN_51[8]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@178825.4]
  assign tlb_OptimizationBarrier_18_io_x_px = tlb__GEN_51[7]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@178825.4]
  assign tlb_OptimizationBarrier_18_io_x_pr = tlb__GEN_51[6]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@178825.4]
  assign tlb_OptimizationBarrier_18_io_x_ppp = tlb__GEN_51[5]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@178825.4]
  assign tlb_OptimizationBarrier_18_io_x_pal = tlb__GEN_51[4]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@178825.4]
  assign tlb_OptimizationBarrier_18_io_x_paa = tlb__GEN_51[3]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@178825.4]
  assign tlb_OptimizationBarrier_18_io_x_eff = tlb__GEN_51[2]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@178825.4]
  assign tlb_OptimizationBarrier_18_io_x_c = tlb__GEN_51[1]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@178825.4]
  assign tlb_OptimizationBarrier_19_io_x_ppn = tlb__GEN_55[34:15]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@178868.4]
  assign tlb_OptimizationBarrier_19_io_x_u = tlb__GEN_55[14]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@178868.4]
  assign tlb_OptimizationBarrier_19_io_x_ae = tlb__GEN_55[12]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@178868.4]
  assign tlb_OptimizationBarrier_19_io_x_sw = tlb__GEN_55[11]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@178868.4]
  assign tlb_OptimizationBarrier_19_io_x_sx = tlb__GEN_55[10]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@178868.4]
  assign tlb_OptimizationBarrier_19_io_x_sr = tlb__GEN_55[9]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@178868.4]
  assign tlb_OptimizationBarrier_19_io_x_pw = tlb__GEN_55[8]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@178868.4]
  assign tlb_OptimizationBarrier_19_io_x_px = tlb__GEN_55[7]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@178868.4]
  assign tlb_OptimizationBarrier_19_io_x_pr = tlb__GEN_55[6]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@178868.4]
  assign tlb_OptimizationBarrier_19_io_x_ppp = tlb__GEN_55[5]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@178868.4]
  assign tlb_OptimizationBarrier_19_io_x_pal = tlb__GEN_55[4]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@178868.4]
  assign tlb_OptimizationBarrier_19_io_x_paa = tlb__GEN_55[3]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@178868.4]
  assign tlb_OptimizationBarrier_19_io_x_eff = tlb__GEN_55[2]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@178868.4]
  assign tlb_OptimizationBarrier_19_io_x_c = tlb__GEN_55[1]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@178868.4]
  assign tlb_OptimizationBarrier_20_io_x_ppn = tlb__GEN_59[34:15]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@178911.4]
  assign tlb_OptimizationBarrier_20_io_x_u = tlb__GEN_59[14]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@178911.4]
  assign tlb_OptimizationBarrier_20_io_x_ae = tlb__GEN_59[12]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@178911.4]
  assign tlb_OptimizationBarrier_20_io_x_sw = tlb__GEN_59[11]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@178911.4]
  assign tlb_OptimizationBarrier_20_io_x_sx = tlb__GEN_59[10]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@178911.4]
  assign tlb_OptimizationBarrier_20_io_x_sr = tlb__GEN_59[9]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@178911.4]
  assign tlb_OptimizationBarrier_20_io_x_pw = tlb__GEN_59[8]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@178911.4]
  assign tlb_OptimizationBarrier_20_io_x_px = tlb__GEN_59[7]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@178911.4]
  assign tlb_OptimizationBarrier_20_io_x_pr = tlb__GEN_59[6]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@178911.4]
  assign tlb_OptimizationBarrier_20_io_x_ppp = tlb__GEN_59[5]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@178911.4]
  assign tlb_OptimizationBarrier_20_io_x_pal = tlb__GEN_59[4]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@178911.4]
  assign tlb_OptimizationBarrier_20_io_x_paa = tlb__GEN_59[3]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@178911.4]
  assign tlb_OptimizationBarrier_20_io_x_eff = tlb__GEN_59[2]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@178911.4]
  assign tlb_OptimizationBarrier_20_io_x_c = tlb__GEN_59[1]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@178911.4]
  assign tlb_OptimizationBarrier_21_io_x_ppn = tlb__GEN_63[34:15]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@178954.4]
  assign tlb_OptimizationBarrier_21_io_x_u = tlb__GEN_63[14]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@178954.4]
  assign tlb_OptimizationBarrier_21_io_x_ae = tlb__GEN_63[12]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@178954.4]
  assign tlb_OptimizationBarrier_21_io_x_sw = tlb__GEN_63[11]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@178954.4]
  assign tlb_OptimizationBarrier_21_io_x_sx = tlb__GEN_63[10]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@178954.4]
  assign tlb_OptimizationBarrier_21_io_x_sr = tlb__GEN_63[9]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@178954.4]
  assign tlb_OptimizationBarrier_21_io_x_pw = tlb__GEN_63[8]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@178954.4]
  assign tlb_OptimizationBarrier_21_io_x_px = tlb__GEN_63[7]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@178954.4]
  assign tlb_OptimizationBarrier_21_io_x_pr = tlb__GEN_63[6]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@178954.4]
  assign tlb_OptimizationBarrier_21_io_x_ppp = tlb__GEN_63[5]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@178954.4]
  assign tlb_OptimizationBarrier_21_io_x_pal = tlb__GEN_63[4]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@178954.4]
  assign tlb_OptimizationBarrier_21_io_x_paa = tlb__GEN_63[3]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@178954.4]
  assign tlb_OptimizationBarrier_21_io_x_eff = tlb__GEN_63[2]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@178954.4]
  assign tlb_OptimizationBarrier_21_io_x_c = tlb__GEN_63[1]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@178954.4]
  assign tlb_OptimizationBarrier_22_io_x_ppn = tlb_superpage_entries_0_data_0[34:15]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@178996.4]
  assign tlb_OptimizationBarrier_22_io_x_u = tlb_superpage_entries_0_data_0[14]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@178996.4]
  assign tlb_OptimizationBarrier_22_io_x_ae = tlb_superpage_entries_0_data_0[12]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@178996.4]
  assign tlb_OptimizationBarrier_22_io_x_sw = tlb_superpage_entries_0_data_0[11]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@178996.4]
  assign tlb_OptimizationBarrier_22_io_x_sx = tlb_superpage_entries_0_data_0[10]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@178996.4]
  assign tlb_OptimizationBarrier_22_io_x_sr = tlb_superpage_entries_0_data_0[9]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@178996.4]
  assign tlb_OptimizationBarrier_22_io_x_pw = tlb_superpage_entries_0_data_0[8]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@178996.4]
  assign tlb_OptimizationBarrier_22_io_x_px = tlb_superpage_entries_0_data_0[7]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@178996.4]
  assign tlb_OptimizationBarrier_22_io_x_pr = tlb_superpage_entries_0_data_0[6]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@178996.4]
  assign tlb_OptimizationBarrier_22_io_x_ppp = tlb_superpage_entries_0_data_0[5]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@178996.4]
  assign tlb_OptimizationBarrier_22_io_x_pal = tlb_superpage_entries_0_data_0[4]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@178996.4]
  assign tlb_OptimizationBarrier_22_io_x_paa = tlb_superpage_entries_0_data_0[3]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@178996.4]
  assign tlb_OptimizationBarrier_22_io_x_eff = tlb_superpage_entries_0_data_0[2]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@178996.4]
  assign tlb_OptimizationBarrier_22_io_x_c = tlb_superpage_entries_0_data_0[1]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@178996.4]
  assign tlb_OptimizationBarrier_23_io_x_ppn = tlb_superpage_entries_1_data_0[34:15]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@179038.4]
  assign tlb_OptimizationBarrier_23_io_x_u = tlb_superpage_entries_1_data_0[14]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@179038.4]
  assign tlb_OptimizationBarrier_23_io_x_ae = tlb_superpage_entries_1_data_0[12]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@179038.4]
  assign tlb_OptimizationBarrier_23_io_x_sw = tlb_superpage_entries_1_data_0[11]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@179038.4]
  assign tlb_OptimizationBarrier_23_io_x_sx = tlb_superpage_entries_1_data_0[10]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@179038.4]
  assign tlb_OptimizationBarrier_23_io_x_sr = tlb_superpage_entries_1_data_0[9]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@179038.4]
  assign tlb_OptimizationBarrier_23_io_x_pw = tlb_superpage_entries_1_data_0[8]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@179038.4]
  assign tlb_OptimizationBarrier_23_io_x_px = tlb_superpage_entries_1_data_0[7]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@179038.4]
  assign tlb_OptimizationBarrier_23_io_x_pr = tlb_superpage_entries_1_data_0[6]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@179038.4]
  assign tlb_OptimizationBarrier_23_io_x_ppp = tlb_superpage_entries_1_data_0[5]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@179038.4]
  assign tlb_OptimizationBarrier_23_io_x_pal = tlb_superpage_entries_1_data_0[4]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@179038.4]
  assign tlb_OptimizationBarrier_23_io_x_paa = tlb_superpage_entries_1_data_0[3]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@179038.4]
  assign tlb_OptimizationBarrier_23_io_x_eff = tlb_superpage_entries_1_data_0[2]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@179038.4]
  assign tlb_OptimizationBarrier_23_io_x_c = tlb_superpage_entries_1_data_0[1]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@179038.4]
  assign tlb_OptimizationBarrier_24_io_x_ppn = tlb_superpage_entries_2_data_0[34:15]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@179080.4]
  assign tlb_OptimizationBarrier_24_io_x_u = tlb_superpage_entries_2_data_0[14]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@179080.4]
  assign tlb_OptimizationBarrier_24_io_x_ae = tlb_superpage_entries_2_data_0[12]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@179080.4]
  assign tlb_OptimizationBarrier_24_io_x_sw = tlb_superpage_entries_2_data_0[11]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@179080.4]
  assign tlb_OptimizationBarrier_24_io_x_sx = tlb_superpage_entries_2_data_0[10]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@179080.4]
  assign tlb_OptimizationBarrier_24_io_x_sr = tlb_superpage_entries_2_data_0[9]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@179080.4]
  assign tlb_OptimizationBarrier_24_io_x_pw = tlb_superpage_entries_2_data_0[8]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@179080.4]
  assign tlb_OptimizationBarrier_24_io_x_px = tlb_superpage_entries_2_data_0[7]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@179080.4]
  assign tlb_OptimizationBarrier_24_io_x_pr = tlb_superpage_entries_2_data_0[6]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@179080.4]
  assign tlb_OptimizationBarrier_24_io_x_ppp = tlb_superpage_entries_2_data_0[5]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@179080.4]
  assign tlb_OptimizationBarrier_24_io_x_pal = tlb_superpage_entries_2_data_0[4]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@179080.4]
  assign tlb_OptimizationBarrier_24_io_x_paa = tlb_superpage_entries_2_data_0[3]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@179080.4]
  assign tlb_OptimizationBarrier_24_io_x_eff = tlb_superpage_entries_2_data_0[2]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@179080.4]
  assign tlb_OptimizationBarrier_24_io_x_c = tlb_superpage_entries_2_data_0[1]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@179080.4]
  assign tlb_OptimizationBarrier_25_io_x_ppn = tlb_superpage_entries_3_data_0[34:15]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@179122.4]
  assign tlb_OptimizationBarrier_25_io_x_u = tlb_superpage_entries_3_data_0[14]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@179122.4]
  assign tlb_OptimizationBarrier_25_io_x_ae = tlb_superpage_entries_3_data_0[12]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@179122.4]
  assign tlb_OptimizationBarrier_25_io_x_sw = tlb_superpage_entries_3_data_0[11]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@179122.4]
  assign tlb_OptimizationBarrier_25_io_x_sx = tlb_superpage_entries_3_data_0[10]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@179122.4]
  assign tlb_OptimizationBarrier_25_io_x_sr = tlb_superpage_entries_3_data_0[9]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@179122.4]
  assign tlb_OptimizationBarrier_25_io_x_pw = tlb_superpage_entries_3_data_0[8]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@179122.4]
  assign tlb_OptimizationBarrier_25_io_x_px = tlb_superpage_entries_3_data_0[7]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@179122.4]
  assign tlb_OptimizationBarrier_25_io_x_pr = tlb_superpage_entries_3_data_0[6]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@179122.4]
  assign tlb_OptimizationBarrier_25_io_x_ppp = tlb_superpage_entries_3_data_0[5]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@179122.4]
  assign tlb_OptimizationBarrier_25_io_x_pal = tlb_superpage_entries_3_data_0[4]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@179122.4]
  assign tlb_OptimizationBarrier_25_io_x_paa = tlb_superpage_entries_3_data_0[3]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@179122.4]
  assign tlb_OptimizationBarrier_25_io_x_eff = tlb_superpage_entries_3_data_0[2]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@179122.4]
  assign tlb_OptimizationBarrier_25_io_x_c = tlb_superpage_entries_3_data_0[1]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@179122.4]
  assign tlb_OptimizationBarrier_26_io_x_ppn = tlb_special_entry_data_0[34:15]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@179164.4]
  assign tlb_OptimizationBarrier_26_io_x_u = tlb_special_entry_data_0[14]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@179164.4]
  assign tlb_OptimizationBarrier_26_io_x_ae = tlb_special_entry_data_0[12]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@179164.4]
  assign tlb_OptimizationBarrier_26_io_x_sw = tlb_special_entry_data_0[11]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@179164.4]
  assign tlb_OptimizationBarrier_26_io_x_sx = tlb_special_entry_data_0[10]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@179164.4]
  assign tlb_OptimizationBarrier_26_io_x_sr = tlb_special_entry_data_0[9]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@179164.4]
  assign tlb_OptimizationBarrier_26_io_x_pw = tlb_special_entry_data_0[8]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@179164.4]
  assign tlb_OptimizationBarrier_26_io_x_px = tlb_special_entry_data_0[7]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@179164.4]
  assign tlb_OptimizationBarrier_26_io_x_pr = tlb_special_entry_data_0[6]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@179164.4]
  assign tlb_OptimizationBarrier_26_io_x_ppp = tlb_special_entry_data_0[5]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@179164.4]
  assign tlb_OptimizationBarrier_26_io_x_pal = tlb_special_entry_data_0[4]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@179164.4]
  assign tlb_OptimizationBarrier_26_io_x_paa = tlb_special_entry_data_0[3]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@179164.4]
  assign tlb_OptimizationBarrier_26_io_x_eff = tlb_special_entry_data_0[2]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@179164.4]
  assign tlb_OptimizationBarrier_26_io_x_c = tlb_special_entry_data_0[1]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@179164.4]
  assign tlb_OptimizationBarrier_27_io_x_ppn = tlb__GEN_35[34:15]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@179207.4]
  assign tlb_OptimizationBarrier_27_io_x_u = tlb__GEN_35[14]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@179207.4]
  assign tlb_OptimizationBarrier_27_io_x_ae = tlb__GEN_35[12]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@179207.4]
  assign tlb_OptimizationBarrier_27_io_x_sw = tlb__GEN_35[11]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@179207.4]
  assign tlb_OptimizationBarrier_27_io_x_sx = tlb__GEN_35[10]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@179207.4]
  assign tlb_OptimizationBarrier_27_io_x_sr = tlb__GEN_35[9]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@179207.4]
  assign tlb_OptimizationBarrier_27_io_x_pw = tlb__GEN_35[8]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@179207.4]
  assign tlb_OptimizationBarrier_27_io_x_px = tlb__GEN_35[7]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@179207.4]
  assign tlb_OptimizationBarrier_27_io_x_pr = tlb__GEN_35[6]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@179207.4]
  assign tlb_OptimizationBarrier_27_io_x_ppp = tlb__GEN_35[5]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@179207.4]
  assign tlb_OptimizationBarrier_27_io_x_pal = tlb__GEN_35[4]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@179207.4]
  assign tlb_OptimizationBarrier_27_io_x_paa = tlb__GEN_35[3]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@179207.4]
  assign tlb_OptimizationBarrier_27_io_x_eff = tlb__GEN_35[2]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@179207.4]
  assign tlb_OptimizationBarrier_27_io_x_c = tlb__GEN_35[1]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@179207.4]
  assign tlb_OptimizationBarrier_28_io_x_ppn = tlb__GEN_39[34:15]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@179250.4]
  assign tlb_OptimizationBarrier_28_io_x_u = tlb__GEN_39[14]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@179250.4]
  assign tlb_OptimizationBarrier_28_io_x_ae = tlb__GEN_39[12]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@179250.4]
  assign tlb_OptimizationBarrier_28_io_x_sw = tlb__GEN_39[11]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@179250.4]
  assign tlb_OptimizationBarrier_28_io_x_sx = tlb__GEN_39[10]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@179250.4]
  assign tlb_OptimizationBarrier_28_io_x_sr = tlb__GEN_39[9]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@179250.4]
  assign tlb_OptimizationBarrier_28_io_x_pw = tlb__GEN_39[8]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@179250.4]
  assign tlb_OptimizationBarrier_28_io_x_px = tlb__GEN_39[7]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@179250.4]
  assign tlb_OptimizationBarrier_28_io_x_pr = tlb__GEN_39[6]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@179250.4]
  assign tlb_OptimizationBarrier_28_io_x_ppp = tlb__GEN_39[5]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@179250.4]
  assign tlb_OptimizationBarrier_28_io_x_pal = tlb__GEN_39[4]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@179250.4]
  assign tlb_OptimizationBarrier_28_io_x_paa = tlb__GEN_39[3]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@179250.4]
  assign tlb_OptimizationBarrier_28_io_x_eff = tlb__GEN_39[2]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@179250.4]
  assign tlb_OptimizationBarrier_28_io_x_c = tlb__GEN_39[1]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@179250.4]
  assign tlb_OptimizationBarrier_29_io_x_ppn = tlb__GEN_43[34:15]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@179293.4]
  assign tlb_OptimizationBarrier_29_io_x_u = tlb__GEN_43[14]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@179293.4]
  assign tlb_OptimizationBarrier_29_io_x_ae = tlb__GEN_43[12]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@179293.4]
  assign tlb_OptimizationBarrier_29_io_x_sw = tlb__GEN_43[11]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@179293.4]
  assign tlb_OptimizationBarrier_29_io_x_sx = tlb__GEN_43[10]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@179293.4]
  assign tlb_OptimizationBarrier_29_io_x_sr = tlb__GEN_43[9]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@179293.4]
  assign tlb_OptimizationBarrier_29_io_x_pw = tlb__GEN_43[8]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@179293.4]
  assign tlb_OptimizationBarrier_29_io_x_px = tlb__GEN_43[7]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@179293.4]
  assign tlb_OptimizationBarrier_29_io_x_pr = tlb__GEN_43[6]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@179293.4]
  assign tlb_OptimizationBarrier_29_io_x_ppp = tlb__GEN_43[5]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@179293.4]
  assign tlb_OptimizationBarrier_29_io_x_pal = tlb__GEN_43[4]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@179293.4]
  assign tlb_OptimizationBarrier_29_io_x_paa = tlb__GEN_43[3]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@179293.4]
  assign tlb_OptimizationBarrier_29_io_x_eff = tlb__GEN_43[2]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@179293.4]
  assign tlb_OptimizationBarrier_29_io_x_c = tlb__GEN_43[1]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@179293.4]
  assign tlb_OptimizationBarrier_30_io_x_ppn = tlb__GEN_47[34:15]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@179336.4]
  assign tlb_OptimizationBarrier_30_io_x_u = tlb__GEN_47[14]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@179336.4]
  assign tlb_OptimizationBarrier_30_io_x_ae = tlb__GEN_47[12]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@179336.4]
  assign tlb_OptimizationBarrier_30_io_x_sw = tlb__GEN_47[11]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@179336.4]
  assign tlb_OptimizationBarrier_30_io_x_sx = tlb__GEN_47[10]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@179336.4]
  assign tlb_OptimizationBarrier_30_io_x_sr = tlb__GEN_47[9]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@179336.4]
  assign tlb_OptimizationBarrier_30_io_x_pw = tlb__GEN_47[8]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@179336.4]
  assign tlb_OptimizationBarrier_30_io_x_px = tlb__GEN_47[7]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@179336.4]
  assign tlb_OptimizationBarrier_30_io_x_pr = tlb__GEN_47[6]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@179336.4]
  assign tlb_OptimizationBarrier_30_io_x_ppp = tlb__GEN_47[5]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@179336.4]
  assign tlb_OptimizationBarrier_30_io_x_pal = tlb__GEN_47[4]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@179336.4]
  assign tlb_OptimizationBarrier_30_io_x_paa = tlb__GEN_47[3]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@179336.4]
  assign tlb_OptimizationBarrier_30_io_x_eff = tlb__GEN_47[2]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@179336.4]
  assign tlb_OptimizationBarrier_30_io_x_c = tlb__GEN_47[1]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@179336.4]
  assign tlb_OptimizationBarrier_31_io_x_ppn = tlb__GEN_51[34:15]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@179379.4]
  assign tlb_OptimizationBarrier_31_io_x_u = tlb__GEN_51[14]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@179379.4]
  assign tlb_OptimizationBarrier_31_io_x_ae = tlb__GEN_51[12]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@179379.4]
  assign tlb_OptimizationBarrier_31_io_x_sw = tlb__GEN_51[11]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@179379.4]
  assign tlb_OptimizationBarrier_31_io_x_sx = tlb__GEN_51[10]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@179379.4]
  assign tlb_OptimizationBarrier_31_io_x_sr = tlb__GEN_51[9]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@179379.4]
  assign tlb_OptimizationBarrier_31_io_x_pw = tlb__GEN_51[8]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@179379.4]
  assign tlb_OptimizationBarrier_31_io_x_px = tlb__GEN_51[7]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@179379.4]
  assign tlb_OptimizationBarrier_31_io_x_pr = tlb__GEN_51[6]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@179379.4]
  assign tlb_OptimizationBarrier_31_io_x_ppp = tlb__GEN_51[5]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@179379.4]
  assign tlb_OptimizationBarrier_31_io_x_pal = tlb__GEN_51[4]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@179379.4]
  assign tlb_OptimizationBarrier_31_io_x_paa = tlb__GEN_51[3]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@179379.4]
  assign tlb_OptimizationBarrier_31_io_x_eff = tlb__GEN_51[2]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@179379.4]
  assign tlb_OptimizationBarrier_31_io_x_c = tlb__GEN_51[1]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@179379.4]
  assign tlb_OptimizationBarrier_32_io_x_ppn = tlb__GEN_55[34:15]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@179422.4]
  assign tlb_OptimizationBarrier_32_io_x_u = tlb__GEN_55[14]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@179422.4]
  assign tlb_OptimizationBarrier_32_io_x_ae = tlb__GEN_55[12]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@179422.4]
  assign tlb_OptimizationBarrier_32_io_x_sw = tlb__GEN_55[11]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@179422.4]
  assign tlb_OptimizationBarrier_32_io_x_sx = tlb__GEN_55[10]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@179422.4]
  assign tlb_OptimizationBarrier_32_io_x_sr = tlb__GEN_55[9]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@179422.4]
  assign tlb_OptimizationBarrier_32_io_x_pw = tlb__GEN_55[8]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@179422.4]
  assign tlb_OptimizationBarrier_32_io_x_px = tlb__GEN_55[7]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@179422.4]
  assign tlb_OptimizationBarrier_32_io_x_pr = tlb__GEN_55[6]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@179422.4]
  assign tlb_OptimizationBarrier_32_io_x_ppp = tlb__GEN_55[5]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@179422.4]
  assign tlb_OptimizationBarrier_32_io_x_pal = tlb__GEN_55[4]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@179422.4]
  assign tlb_OptimizationBarrier_32_io_x_paa = tlb__GEN_55[3]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@179422.4]
  assign tlb_OptimizationBarrier_32_io_x_eff = tlb__GEN_55[2]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@179422.4]
  assign tlb_OptimizationBarrier_32_io_x_c = tlb__GEN_55[1]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@179422.4]
  assign tlb_OptimizationBarrier_33_io_x_ppn = tlb__GEN_59[34:15]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@179465.4]
  assign tlb_OptimizationBarrier_33_io_x_u = tlb__GEN_59[14]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@179465.4]
  assign tlb_OptimizationBarrier_33_io_x_ae = tlb__GEN_59[12]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@179465.4]
  assign tlb_OptimizationBarrier_33_io_x_sw = tlb__GEN_59[11]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@179465.4]
  assign tlb_OptimizationBarrier_33_io_x_sx = tlb__GEN_59[10]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@179465.4]
  assign tlb_OptimizationBarrier_33_io_x_sr = tlb__GEN_59[9]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@179465.4]
  assign tlb_OptimizationBarrier_33_io_x_pw = tlb__GEN_59[8]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@179465.4]
  assign tlb_OptimizationBarrier_33_io_x_px = tlb__GEN_59[7]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@179465.4]
  assign tlb_OptimizationBarrier_33_io_x_pr = tlb__GEN_59[6]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@179465.4]
  assign tlb_OptimizationBarrier_33_io_x_ppp = tlb__GEN_59[5]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@179465.4]
  assign tlb_OptimizationBarrier_33_io_x_pal = tlb__GEN_59[4]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@179465.4]
  assign tlb_OptimizationBarrier_33_io_x_paa = tlb__GEN_59[3]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@179465.4]
  assign tlb_OptimizationBarrier_33_io_x_eff = tlb__GEN_59[2]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@179465.4]
  assign tlb_OptimizationBarrier_33_io_x_c = tlb__GEN_59[1]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@179465.4]
  assign tlb_OptimizationBarrier_34_io_x_ppn = tlb__GEN_63[34:15]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@179508.4]
  assign tlb_OptimizationBarrier_34_io_x_u = tlb__GEN_63[14]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@179508.4]
  assign tlb_OptimizationBarrier_34_io_x_ae = tlb__GEN_63[12]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@179508.4]
  assign tlb_OptimizationBarrier_34_io_x_sw = tlb__GEN_63[11]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@179508.4]
  assign tlb_OptimizationBarrier_34_io_x_sx = tlb__GEN_63[10]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@179508.4]
  assign tlb_OptimizationBarrier_34_io_x_sr = tlb__GEN_63[9]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@179508.4]
  assign tlb_OptimizationBarrier_34_io_x_pw = tlb__GEN_63[8]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@179508.4]
  assign tlb_OptimizationBarrier_34_io_x_px = tlb__GEN_63[7]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@179508.4]
  assign tlb_OptimizationBarrier_34_io_x_pr = tlb__GEN_63[6]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@179508.4]
  assign tlb_OptimizationBarrier_34_io_x_ppp = tlb__GEN_63[5]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@179508.4]
  assign tlb_OptimizationBarrier_34_io_x_pal = tlb__GEN_63[4]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@179508.4]
  assign tlb_OptimizationBarrier_34_io_x_paa = tlb__GEN_63[3]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@179508.4]
  assign tlb_OptimizationBarrier_34_io_x_eff = tlb__GEN_63[2]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@179508.4]
  assign tlb_OptimizationBarrier_34_io_x_c = tlb__GEN_63[1]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@179508.4]
  assign tlb_OptimizationBarrier_35_io_x_ppn = tlb_superpage_entries_0_data_0[34:15]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@179550.4]
  assign tlb_OptimizationBarrier_35_io_x_u = tlb_superpage_entries_0_data_0[14]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@179550.4]
  assign tlb_OptimizationBarrier_35_io_x_ae = tlb_superpage_entries_0_data_0[12]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@179550.4]
  assign tlb_OptimizationBarrier_35_io_x_sw = tlb_superpage_entries_0_data_0[11]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@179550.4]
  assign tlb_OptimizationBarrier_35_io_x_sx = tlb_superpage_entries_0_data_0[10]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@179550.4]
  assign tlb_OptimizationBarrier_35_io_x_sr = tlb_superpage_entries_0_data_0[9]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@179550.4]
  assign tlb_OptimizationBarrier_35_io_x_pw = tlb_superpage_entries_0_data_0[8]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@179550.4]
  assign tlb_OptimizationBarrier_35_io_x_px = tlb_superpage_entries_0_data_0[7]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@179550.4]
  assign tlb_OptimizationBarrier_35_io_x_pr = tlb_superpage_entries_0_data_0[6]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@179550.4]
  assign tlb_OptimizationBarrier_35_io_x_ppp = tlb_superpage_entries_0_data_0[5]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@179550.4]
  assign tlb_OptimizationBarrier_35_io_x_pal = tlb_superpage_entries_0_data_0[4]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@179550.4]
  assign tlb_OptimizationBarrier_35_io_x_paa = tlb_superpage_entries_0_data_0[3]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@179550.4]
  assign tlb_OptimizationBarrier_35_io_x_eff = tlb_superpage_entries_0_data_0[2]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@179550.4]
  assign tlb_OptimizationBarrier_35_io_x_c = tlb_superpage_entries_0_data_0[1]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@179550.4]
  assign tlb_OptimizationBarrier_36_io_x_ppn = tlb_superpage_entries_1_data_0[34:15]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@179592.4]
  assign tlb_OptimizationBarrier_36_io_x_u = tlb_superpage_entries_1_data_0[14]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@179592.4]
  assign tlb_OptimizationBarrier_36_io_x_ae = tlb_superpage_entries_1_data_0[12]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@179592.4]
  assign tlb_OptimizationBarrier_36_io_x_sw = tlb_superpage_entries_1_data_0[11]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@179592.4]
  assign tlb_OptimizationBarrier_36_io_x_sx = tlb_superpage_entries_1_data_0[10]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@179592.4]
  assign tlb_OptimizationBarrier_36_io_x_sr = tlb_superpage_entries_1_data_0[9]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@179592.4]
  assign tlb_OptimizationBarrier_36_io_x_pw = tlb_superpage_entries_1_data_0[8]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@179592.4]
  assign tlb_OptimizationBarrier_36_io_x_px = tlb_superpage_entries_1_data_0[7]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@179592.4]
  assign tlb_OptimizationBarrier_36_io_x_pr = tlb_superpage_entries_1_data_0[6]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@179592.4]
  assign tlb_OptimizationBarrier_36_io_x_ppp = tlb_superpage_entries_1_data_0[5]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@179592.4]
  assign tlb_OptimizationBarrier_36_io_x_pal = tlb_superpage_entries_1_data_0[4]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@179592.4]
  assign tlb_OptimizationBarrier_36_io_x_paa = tlb_superpage_entries_1_data_0[3]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@179592.4]
  assign tlb_OptimizationBarrier_36_io_x_eff = tlb_superpage_entries_1_data_0[2]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@179592.4]
  assign tlb_OptimizationBarrier_36_io_x_c = tlb_superpage_entries_1_data_0[1]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@179592.4]
  assign tlb_OptimizationBarrier_37_io_x_ppn = tlb_superpage_entries_2_data_0[34:15]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@179634.4]
  assign tlb_OptimizationBarrier_37_io_x_u = tlb_superpage_entries_2_data_0[14]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@179634.4]
  assign tlb_OptimizationBarrier_37_io_x_ae = tlb_superpage_entries_2_data_0[12]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@179634.4]
  assign tlb_OptimizationBarrier_37_io_x_sw = tlb_superpage_entries_2_data_0[11]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@179634.4]
  assign tlb_OptimizationBarrier_37_io_x_sx = tlb_superpage_entries_2_data_0[10]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@179634.4]
  assign tlb_OptimizationBarrier_37_io_x_sr = tlb_superpage_entries_2_data_0[9]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@179634.4]
  assign tlb_OptimizationBarrier_37_io_x_pw = tlb_superpage_entries_2_data_0[8]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@179634.4]
  assign tlb_OptimizationBarrier_37_io_x_px = tlb_superpage_entries_2_data_0[7]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@179634.4]
  assign tlb_OptimizationBarrier_37_io_x_pr = tlb_superpage_entries_2_data_0[6]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@179634.4]
  assign tlb_OptimizationBarrier_37_io_x_ppp = tlb_superpage_entries_2_data_0[5]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@179634.4]
  assign tlb_OptimizationBarrier_37_io_x_pal = tlb_superpage_entries_2_data_0[4]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@179634.4]
  assign tlb_OptimizationBarrier_37_io_x_paa = tlb_superpage_entries_2_data_0[3]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@179634.4]
  assign tlb_OptimizationBarrier_37_io_x_eff = tlb_superpage_entries_2_data_0[2]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@179634.4]
  assign tlb_OptimizationBarrier_37_io_x_c = tlb_superpage_entries_2_data_0[1]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@179634.4]
  assign tlb_OptimizationBarrier_38_io_x_ppn = tlb_superpage_entries_3_data_0[34:15]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@179676.4]
  assign tlb_OptimizationBarrier_38_io_x_u = tlb_superpage_entries_3_data_0[14]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@179676.4]
  assign tlb_OptimizationBarrier_38_io_x_ae = tlb_superpage_entries_3_data_0[12]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@179676.4]
  assign tlb_OptimizationBarrier_38_io_x_sw = tlb_superpage_entries_3_data_0[11]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@179676.4]
  assign tlb_OptimizationBarrier_38_io_x_sx = tlb_superpage_entries_3_data_0[10]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@179676.4]
  assign tlb_OptimizationBarrier_38_io_x_sr = tlb_superpage_entries_3_data_0[9]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@179676.4]
  assign tlb_OptimizationBarrier_38_io_x_pw = tlb_superpage_entries_3_data_0[8]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@179676.4]
  assign tlb_OptimizationBarrier_38_io_x_px = tlb_superpage_entries_3_data_0[7]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@179676.4]
  assign tlb_OptimizationBarrier_38_io_x_pr = tlb_superpage_entries_3_data_0[6]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@179676.4]
  assign tlb_OptimizationBarrier_38_io_x_ppp = tlb_superpage_entries_3_data_0[5]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@179676.4]
  assign tlb_OptimizationBarrier_38_io_x_pal = tlb_superpage_entries_3_data_0[4]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@179676.4]
  assign tlb_OptimizationBarrier_38_io_x_paa = tlb_superpage_entries_3_data_0[3]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@179676.4]
  assign tlb_OptimizationBarrier_38_io_x_eff = tlb_superpage_entries_3_data_0[2]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@179676.4]
  assign tlb_OptimizationBarrier_38_io_x_c = tlb_superpage_entries_3_data_0[1]; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@179676.4]
  assign pma_checker__T_2026 = |4'h0; // @[OneHot.scala 32:14:freechips.rocketchip.system.DefaultRV32Config.fir@180088.8]
  assign pma_checker_OptimizationBarrier_io_x_ppn = 20'h0; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@176911.4]
  assign pma_checker_OptimizationBarrier_io_x_u = 1'h0; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@176911.4]
  assign pma_checker_OptimizationBarrier_io_x_ae = 1'h0; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@176911.4]
  assign pma_checker_OptimizationBarrier_io_x_sw = 1'h0; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@176911.4]
  assign pma_checker_OptimizationBarrier_io_x_sx = 1'h0; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@176911.4]
  assign pma_checker_OptimizationBarrier_io_x_sr = 1'h0; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@176911.4]
  assign pma_checker_OptimizationBarrier_io_x_pw = 1'h0; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@176911.4]
  assign pma_checker_OptimizationBarrier_io_x_px = 1'h0; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@176911.4]
  assign pma_checker_OptimizationBarrier_io_x_pr = 1'h0; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@176911.4]
  assign pma_checker_OptimizationBarrier_io_x_ppp = 1'h0; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@176911.4]
  assign pma_checker_OptimizationBarrier_io_x_pal = 1'h0; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@176911.4]
  assign pma_checker_OptimizationBarrier_io_x_paa = 1'h0; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@176911.4]
  assign pma_checker_OptimizationBarrier_io_x_eff = 1'h0; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@176911.4]
  assign pma_checker_OptimizationBarrier_io_x_c = 1'h0; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@176911.4]
  assign pma_checker_pmp_io_prv = 2'h1; // @[TLB.scala 194:14:freechips.rocketchip.system.DefaultRV32Config.fir@176942.4]
  assign pma_checker_pmp_io_pmp_0_cfg_l = 1'h0; // @[TLB.scala 193:14:freechips.rocketchip.system.DefaultRV32Config.fir@176934.4]
  assign pma_checker_pmp_io_pmp_0_cfg_a = 2'h0; // @[TLB.scala 193:14:freechips.rocketchip.system.DefaultRV32Config.fir@176934.4]
  assign pma_checker_pmp_io_pmp_0_cfg_x = 1'h0; // @[TLB.scala 193:14:freechips.rocketchip.system.DefaultRV32Config.fir@176934.4]
  assign pma_checker_pmp_io_pmp_0_cfg_w = 1'h0; // @[TLB.scala 193:14:freechips.rocketchip.system.DefaultRV32Config.fir@176934.4]
  assign pma_checker_pmp_io_pmp_0_cfg_r = 1'h0; // @[TLB.scala 193:14:freechips.rocketchip.system.DefaultRV32Config.fir@176934.4]
  assign pma_checker_pmp_io_pmp_0_addr = 30'h0; // @[TLB.scala 193:14:freechips.rocketchip.system.DefaultRV32Config.fir@176934.4]
  assign pma_checker_pmp_io_pmp_0_mask = 32'h0; // @[TLB.scala 193:14:freechips.rocketchip.system.DefaultRV32Config.fir@176934.4]
  assign pma_checker_pmp_io_pmp_1_cfg_l = 1'h0; // @[TLB.scala 193:14:freechips.rocketchip.system.DefaultRV32Config.fir@176935.4]
  assign pma_checker_pmp_io_pmp_1_cfg_a = 2'h0; // @[TLB.scala 193:14:freechips.rocketchip.system.DefaultRV32Config.fir@176935.4]
  assign pma_checker_pmp_io_pmp_1_cfg_x = 1'h0; // @[TLB.scala 193:14:freechips.rocketchip.system.DefaultRV32Config.fir@176935.4]
  assign pma_checker_pmp_io_pmp_1_cfg_w = 1'h0; // @[TLB.scala 193:14:freechips.rocketchip.system.DefaultRV32Config.fir@176935.4]
  assign pma_checker_pmp_io_pmp_1_cfg_r = 1'h0; // @[TLB.scala 193:14:freechips.rocketchip.system.DefaultRV32Config.fir@176935.4]
  assign pma_checker_pmp_io_pmp_1_addr = 30'h0; // @[TLB.scala 193:14:freechips.rocketchip.system.DefaultRV32Config.fir@176935.4]
  assign pma_checker_pmp_io_pmp_1_mask = 32'h0; // @[TLB.scala 193:14:freechips.rocketchip.system.DefaultRV32Config.fir@176935.4]
  assign pma_checker_pmp_io_pmp_2_cfg_l = 1'h0; // @[TLB.scala 193:14:freechips.rocketchip.system.DefaultRV32Config.fir@176936.4]
  assign pma_checker_pmp_io_pmp_2_cfg_a = 2'h0; // @[TLB.scala 193:14:freechips.rocketchip.system.DefaultRV32Config.fir@176936.4]
  assign pma_checker_pmp_io_pmp_2_cfg_x = 1'h0; // @[TLB.scala 193:14:freechips.rocketchip.system.DefaultRV32Config.fir@176936.4]
  assign pma_checker_pmp_io_pmp_2_cfg_w = 1'h0; // @[TLB.scala 193:14:freechips.rocketchip.system.DefaultRV32Config.fir@176936.4]
  assign pma_checker_pmp_io_pmp_2_cfg_r = 1'h0; // @[TLB.scala 193:14:freechips.rocketchip.system.DefaultRV32Config.fir@176936.4]
  assign pma_checker_pmp_io_pmp_2_addr = 30'h0; // @[TLB.scala 193:14:freechips.rocketchip.system.DefaultRV32Config.fir@176936.4]
  assign pma_checker_pmp_io_pmp_2_mask = 32'h0; // @[TLB.scala 193:14:freechips.rocketchip.system.DefaultRV32Config.fir@176936.4]
  assign pma_checker_pmp_io_pmp_3_cfg_l = 1'h0; // @[TLB.scala 193:14:freechips.rocketchip.system.DefaultRV32Config.fir@176937.4]
  assign pma_checker_pmp_io_pmp_3_cfg_a = 2'h0; // @[TLB.scala 193:14:freechips.rocketchip.system.DefaultRV32Config.fir@176937.4]
  assign pma_checker_pmp_io_pmp_3_cfg_x = 1'h0; // @[TLB.scala 193:14:freechips.rocketchip.system.DefaultRV32Config.fir@176937.4]
  assign pma_checker_pmp_io_pmp_3_cfg_w = 1'h0; // @[TLB.scala 193:14:freechips.rocketchip.system.DefaultRV32Config.fir@176937.4]
  assign pma_checker_pmp_io_pmp_3_cfg_r = 1'h0; // @[TLB.scala 193:14:freechips.rocketchip.system.DefaultRV32Config.fir@176937.4]
  assign pma_checker_pmp_io_pmp_3_addr = 30'h0; // @[TLB.scala 193:14:freechips.rocketchip.system.DefaultRV32Config.fir@176937.4]
  assign pma_checker_pmp_io_pmp_3_mask = 32'h0; // @[TLB.scala 193:14:freechips.rocketchip.system.DefaultRV32Config.fir@176937.4]
  assign pma_checker_pmp_io_pmp_4_cfg_l = 1'h0; // @[TLB.scala 193:14:freechips.rocketchip.system.DefaultRV32Config.fir@176938.4]
  assign pma_checker_pmp_io_pmp_4_cfg_a = 2'h0; // @[TLB.scala 193:14:freechips.rocketchip.system.DefaultRV32Config.fir@176938.4]
  assign pma_checker_pmp_io_pmp_4_cfg_x = 1'h0; // @[TLB.scala 193:14:freechips.rocketchip.system.DefaultRV32Config.fir@176938.4]
  assign pma_checker_pmp_io_pmp_4_cfg_w = 1'h0; // @[TLB.scala 193:14:freechips.rocketchip.system.DefaultRV32Config.fir@176938.4]
  assign pma_checker_pmp_io_pmp_4_cfg_r = 1'h0; // @[TLB.scala 193:14:freechips.rocketchip.system.DefaultRV32Config.fir@176938.4]
  assign pma_checker_pmp_io_pmp_4_addr = 30'h0; // @[TLB.scala 193:14:freechips.rocketchip.system.DefaultRV32Config.fir@176938.4]
  assign pma_checker_pmp_io_pmp_4_mask = 32'h0; // @[TLB.scala 193:14:freechips.rocketchip.system.DefaultRV32Config.fir@176938.4]
  assign pma_checker_pmp_io_pmp_5_cfg_l = 1'h0; // @[TLB.scala 193:14:freechips.rocketchip.system.DefaultRV32Config.fir@176939.4]
  assign pma_checker_pmp_io_pmp_5_cfg_a = 2'h0; // @[TLB.scala 193:14:freechips.rocketchip.system.DefaultRV32Config.fir@176939.4]
  assign pma_checker_pmp_io_pmp_5_cfg_x = 1'h0; // @[TLB.scala 193:14:freechips.rocketchip.system.DefaultRV32Config.fir@176939.4]
  assign pma_checker_pmp_io_pmp_5_cfg_w = 1'h0; // @[TLB.scala 193:14:freechips.rocketchip.system.DefaultRV32Config.fir@176939.4]
  assign pma_checker_pmp_io_pmp_5_cfg_r = 1'h0; // @[TLB.scala 193:14:freechips.rocketchip.system.DefaultRV32Config.fir@176939.4]
  assign pma_checker_pmp_io_pmp_5_addr = 30'h0; // @[TLB.scala 193:14:freechips.rocketchip.system.DefaultRV32Config.fir@176939.4]
  assign pma_checker_pmp_io_pmp_5_mask = 32'h0; // @[TLB.scala 193:14:freechips.rocketchip.system.DefaultRV32Config.fir@176939.4]
  assign pma_checker_pmp_io_pmp_6_cfg_l = 1'h0; // @[TLB.scala 193:14:freechips.rocketchip.system.DefaultRV32Config.fir@176940.4]
  assign pma_checker_pmp_io_pmp_6_cfg_a = 2'h0; // @[TLB.scala 193:14:freechips.rocketchip.system.DefaultRV32Config.fir@176940.4]
  assign pma_checker_pmp_io_pmp_6_cfg_x = 1'h0; // @[TLB.scala 193:14:freechips.rocketchip.system.DefaultRV32Config.fir@176940.4]
  assign pma_checker_pmp_io_pmp_6_cfg_w = 1'h0; // @[TLB.scala 193:14:freechips.rocketchip.system.DefaultRV32Config.fir@176940.4]
  assign pma_checker_pmp_io_pmp_6_cfg_r = 1'h0; // @[TLB.scala 193:14:freechips.rocketchip.system.DefaultRV32Config.fir@176940.4]
  assign pma_checker_pmp_io_pmp_6_addr = 30'h0; // @[TLB.scala 193:14:freechips.rocketchip.system.DefaultRV32Config.fir@176940.4]
  assign pma_checker_pmp_io_pmp_6_mask = 32'h0; // @[TLB.scala 193:14:freechips.rocketchip.system.DefaultRV32Config.fir@176940.4]
  assign pma_checker_pmp_io_pmp_7_cfg_l = 1'h0; // @[TLB.scala 193:14:freechips.rocketchip.system.DefaultRV32Config.fir@176941.4]
  assign pma_checker_pmp_io_pmp_7_cfg_a = 2'h0; // @[TLB.scala 193:14:freechips.rocketchip.system.DefaultRV32Config.fir@176941.4]
  assign pma_checker_pmp_io_pmp_7_cfg_x = 1'h0; // @[TLB.scala 193:14:freechips.rocketchip.system.DefaultRV32Config.fir@176941.4]
  assign pma_checker_pmp_io_pmp_7_cfg_w = 1'h0; // @[TLB.scala 193:14:freechips.rocketchip.system.DefaultRV32Config.fir@176941.4]
  assign pma_checker_pmp_io_pmp_7_cfg_r = 1'h0; // @[TLB.scala 193:14:freechips.rocketchip.system.DefaultRV32Config.fir@176941.4]
  assign pma_checker_pmp_io_pmp_7_addr = 30'h0; // @[TLB.scala 193:14:freechips.rocketchip.system.DefaultRV32Config.fir@176941.4]
  assign pma_checker_pmp_io_pmp_7_mask = 32'h0; // @[TLB.scala 193:14:freechips.rocketchip.system.DefaultRV32Config.fir@176941.4]
  assign pma_checker_pmp_io_addr = 32'h0; // @[TLB.scala 191:15:freechips.rocketchip.system.DefaultRV32Config.fir@176932.4]
  assign pma_checker_OptimizationBarrier_1_io_x_ppn = 20'h0; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@177633.4]
  assign pma_checker_OptimizationBarrier_1_io_x_u = 1'h0; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@177633.4]
  assign pma_checker_OptimizationBarrier_1_io_x_ae = 1'h0; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@177633.4]
  assign pma_checker_OptimizationBarrier_1_io_x_sw = 1'h0; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@177633.4]
  assign pma_checker_OptimizationBarrier_1_io_x_sx = 1'h0; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@177633.4]
  assign pma_checker_OptimizationBarrier_1_io_x_sr = 1'h0; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@177633.4]
  assign pma_checker_OptimizationBarrier_1_io_x_pw = 1'h0; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@177633.4]
  assign pma_checker_OptimizationBarrier_1_io_x_px = 1'h0; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@177633.4]
  assign pma_checker_OptimizationBarrier_1_io_x_pr = 1'h0; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@177633.4]
  assign pma_checker_OptimizationBarrier_1_io_x_ppp = 1'h0; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@177633.4]
  assign pma_checker_OptimizationBarrier_1_io_x_pal = 1'h0; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@177633.4]
  assign pma_checker_OptimizationBarrier_1_io_x_paa = 1'h0; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@177633.4]
  assign pma_checker_OptimizationBarrier_1_io_x_eff = 1'h0; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@177633.4]
  assign pma_checker_OptimizationBarrier_1_io_x_c = 1'h0; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@177633.4]
  assign pma_checker_OptimizationBarrier_2_io_x_ppn = 20'h0; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@177676.4]
  assign pma_checker_OptimizationBarrier_2_io_x_u = 1'h0; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@177676.4]
  assign pma_checker_OptimizationBarrier_2_io_x_ae = 1'h0; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@177676.4]
  assign pma_checker_OptimizationBarrier_2_io_x_sw = 1'h0; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@177676.4]
  assign pma_checker_OptimizationBarrier_2_io_x_sx = 1'h0; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@177676.4]
  assign pma_checker_OptimizationBarrier_2_io_x_sr = 1'h0; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@177676.4]
  assign pma_checker_OptimizationBarrier_2_io_x_pw = 1'h0; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@177676.4]
  assign pma_checker_OptimizationBarrier_2_io_x_px = 1'h0; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@177676.4]
  assign pma_checker_OptimizationBarrier_2_io_x_pr = 1'h0; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@177676.4]
  assign pma_checker_OptimizationBarrier_2_io_x_ppp = 1'h0; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@177676.4]
  assign pma_checker_OptimizationBarrier_2_io_x_pal = 1'h0; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@177676.4]
  assign pma_checker_OptimizationBarrier_2_io_x_paa = 1'h0; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@177676.4]
  assign pma_checker_OptimizationBarrier_2_io_x_eff = 1'h0; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@177676.4]
  assign pma_checker_OptimizationBarrier_2_io_x_c = 1'h0; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@177676.4]
  assign pma_checker_OptimizationBarrier_3_io_x_ppn = 20'h0; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@177719.4]
  assign pma_checker_OptimizationBarrier_3_io_x_u = 1'h0; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@177719.4]
  assign pma_checker_OptimizationBarrier_3_io_x_ae = 1'h0; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@177719.4]
  assign pma_checker_OptimizationBarrier_3_io_x_sw = 1'h0; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@177719.4]
  assign pma_checker_OptimizationBarrier_3_io_x_sx = 1'h0; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@177719.4]
  assign pma_checker_OptimizationBarrier_3_io_x_sr = 1'h0; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@177719.4]
  assign pma_checker_OptimizationBarrier_3_io_x_pw = 1'h0; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@177719.4]
  assign pma_checker_OptimizationBarrier_3_io_x_px = 1'h0; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@177719.4]
  assign pma_checker_OptimizationBarrier_3_io_x_pr = 1'h0; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@177719.4]
  assign pma_checker_OptimizationBarrier_3_io_x_ppp = 1'h0; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@177719.4]
  assign pma_checker_OptimizationBarrier_3_io_x_pal = 1'h0; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@177719.4]
  assign pma_checker_OptimizationBarrier_3_io_x_paa = 1'h0; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@177719.4]
  assign pma_checker_OptimizationBarrier_3_io_x_eff = 1'h0; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@177719.4]
  assign pma_checker_OptimizationBarrier_3_io_x_c = 1'h0; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@177719.4]
  assign pma_checker_OptimizationBarrier_4_io_x_ppn = 20'h0; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@177762.4]
  assign pma_checker_OptimizationBarrier_4_io_x_u = 1'h0; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@177762.4]
  assign pma_checker_OptimizationBarrier_4_io_x_ae = 1'h0; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@177762.4]
  assign pma_checker_OptimizationBarrier_4_io_x_sw = 1'h0; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@177762.4]
  assign pma_checker_OptimizationBarrier_4_io_x_sx = 1'h0; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@177762.4]
  assign pma_checker_OptimizationBarrier_4_io_x_sr = 1'h0; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@177762.4]
  assign pma_checker_OptimizationBarrier_4_io_x_pw = 1'h0; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@177762.4]
  assign pma_checker_OptimizationBarrier_4_io_x_px = 1'h0; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@177762.4]
  assign pma_checker_OptimizationBarrier_4_io_x_pr = 1'h0; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@177762.4]
  assign pma_checker_OptimizationBarrier_4_io_x_ppp = 1'h0; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@177762.4]
  assign pma_checker_OptimizationBarrier_4_io_x_pal = 1'h0; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@177762.4]
  assign pma_checker_OptimizationBarrier_4_io_x_paa = 1'h0; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@177762.4]
  assign pma_checker_OptimizationBarrier_4_io_x_eff = 1'h0; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@177762.4]
  assign pma_checker_OptimizationBarrier_4_io_x_c = 1'h0; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@177762.4]
  assign pma_checker_OptimizationBarrier_5_io_x_ppn = 20'h0; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@177805.4]
  assign pma_checker_OptimizationBarrier_5_io_x_u = 1'h0; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@177805.4]
  assign pma_checker_OptimizationBarrier_5_io_x_ae = 1'h0; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@177805.4]
  assign pma_checker_OptimizationBarrier_5_io_x_sw = 1'h0; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@177805.4]
  assign pma_checker_OptimizationBarrier_5_io_x_sx = 1'h0; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@177805.4]
  assign pma_checker_OptimizationBarrier_5_io_x_sr = 1'h0; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@177805.4]
  assign pma_checker_OptimizationBarrier_5_io_x_pw = 1'h0; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@177805.4]
  assign pma_checker_OptimizationBarrier_5_io_x_px = 1'h0; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@177805.4]
  assign pma_checker_OptimizationBarrier_5_io_x_pr = 1'h0; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@177805.4]
  assign pma_checker_OptimizationBarrier_5_io_x_ppp = 1'h0; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@177805.4]
  assign pma_checker_OptimizationBarrier_5_io_x_pal = 1'h0; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@177805.4]
  assign pma_checker_OptimizationBarrier_5_io_x_paa = 1'h0; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@177805.4]
  assign pma_checker_OptimizationBarrier_5_io_x_eff = 1'h0; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@177805.4]
  assign pma_checker_OptimizationBarrier_5_io_x_c = 1'h0; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@177805.4]
  assign pma_checker_OptimizationBarrier_6_io_x_ppn = 20'h0; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@177848.4]
  assign pma_checker_OptimizationBarrier_6_io_x_u = 1'h0; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@177848.4]
  assign pma_checker_OptimizationBarrier_6_io_x_ae = 1'h0; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@177848.4]
  assign pma_checker_OptimizationBarrier_6_io_x_sw = 1'h0; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@177848.4]
  assign pma_checker_OptimizationBarrier_6_io_x_sx = 1'h0; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@177848.4]
  assign pma_checker_OptimizationBarrier_6_io_x_sr = 1'h0; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@177848.4]
  assign pma_checker_OptimizationBarrier_6_io_x_pw = 1'h0; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@177848.4]
  assign pma_checker_OptimizationBarrier_6_io_x_px = 1'h0; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@177848.4]
  assign pma_checker_OptimizationBarrier_6_io_x_pr = 1'h0; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@177848.4]
  assign pma_checker_OptimizationBarrier_6_io_x_ppp = 1'h0; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@177848.4]
  assign pma_checker_OptimizationBarrier_6_io_x_pal = 1'h0; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@177848.4]
  assign pma_checker_OptimizationBarrier_6_io_x_paa = 1'h0; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@177848.4]
  assign pma_checker_OptimizationBarrier_6_io_x_eff = 1'h0; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@177848.4]
  assign pma_checker_OptimizationBarrier_6_io_x_c = 1'h0; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@177848.4]
  assign pma_checker_OptimizationBarrier_7_io_x_ppn = 20'h0; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@177891.4]
  assign pma_checker_OptimizationBarrier_7_io_x_u = 1'h0; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@177891.4]
  assign pma_checker_OptimizationBarrier_7_io_x_ae = 1'h0; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@177891.4]
  assign pma_checker_OptimizationBarrier_7_io_x_sw = 1'h0; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@177891.4]
  assign pma_checker_OptimizationBarrier_7_io_x_sx = 1'h0; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@177891.4]
  assign pma_checker_OptimizationBarrier_7_io_x_sr = 1'h0; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@177891.4]
  assign pma_checker_OptimizationBarrier_7_io_x_pw = 1'h0; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@177891.4]
  assign pma_checker_OptimizationBarrier_7_io_x_px = 1'h0; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@177891.4]
  assign pma_checker_OptimizationBarrier_7_io_x_pr = 1'h0; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@177891.4]
  assign pma_checker_OptimizationBarrier_7_io_x_ppp = 1'h0; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@177891.4]
  assign pma_checker_OptimizationBarrier_7_io_x_pal = 1'h0; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@177891.4]
  assign pma_checker_OptimizationBarrier_7_io_x_paa = 1'h0; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@177891.4]
  assign pma_checker_OptimizationBarrier_7_io_x_eff = 1'h0; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@177891.4]
  assign pma_checker_OptimizationBarrier_7_io_x_c = 1'h0; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@177891.4]
  assign pma_checker_OptimizationBarrier_8_io_x_ppn = 20'h0; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@177934.4]
  assign pma_checker_OptimizationBarrier_8_io_x_u = 1'h0; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@177934.4]
  assign pma_checker_OptimizationBarrier_8_io_x_ae = 1'h0; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@177934.4]
  assign pma_checker_OptimizationBarrier_8_io_x_sw = 1'h0; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@177934.4]
  assign pma_checker_OptimizationBarrier_8_io_x_sx = 1'h0; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@177934.4]
  assign pma_checker_OptimizationBarrier_8_io_x_sr = 1'h0; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@177934.4]
  assign pma_checker_OptimizationBarrier_8_io_x_pw = 1'h0; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@177934.4]
  assign pma_checker_OptimizationBarrier_8_io_x_px = 1'h0; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@177934.4]
  assign pma_checker_OptimizationBarrier_8_io_x_pr = 1'h0; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@177934.4]
  assign pma_checker_OptimizationBarrier_8_io_x_ppp = 1'h0; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@177934.4]
  assign pma_checker_OptimizationBarrier_8_io_x_pal = 1'h0; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@177934.4]
  assign pma_checker_OptimizationBarrier_8_io_x_paa = 1'h0; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@177934.4]
  assign pma_checker_OptimizationBarrier_8_io_x_eff = 1'h0; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@177934.4]
  assign pma_checker_OptimizationBarrier_8_io_x_c = 1'h0; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@177934.4]
  assign pma_checker_OptimizationBarrier_9_io_x_ppn = 20'h0; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@177976.4]
  assign pma_checker_OptimizationBarrier_9_io_x_u = 1'h0; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@177976.4]
  assign pma_checker_OptimizationBarrier_9_io_x_ae = 1'h0; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@177976.4]
  assign pma_checker_OptimizationBarrier_9_io_x_sw = 1'h0; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@177976.4]
  assign pma_checker_OptimizationBarrier_9_io_x_sx = 1'h0; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@177976.4]
  assign pma_checker_OptimizationBarrier_9_io_x_sr = 1'h0; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@177976.4]
  assign pma_checker_OptimizationBarrier_9_io_x_pw = 1'h0; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@177976.4]
  assign pma_checker_OptimizationBarrier_9_io_x_px = 1'h0; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@177976.4]
  assign pma_checker_OptimizationBarrier_9_io_x_pr = 1'h0; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@177976.4]
  assign pma_checker_OptimizationBarrier_9_io_x_ppp = 1'h0; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@177976.4]
  assign pma_checker_OptimizationBarrier_9_io_x_pal = 1'h0; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@177976.4]
  assign pma_checker_OptimizationBarrier_9_io_x_paa = 1'h0; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@177976.4]
  assign pma_checker_OptimizationBarrier_9_io_x_eff = 1'h0; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@177976.4]
  assign pma_checker_OptimizationBarrier_9_io_x_c = 1'h0; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@177976.4]
  assign pma_checker_OptimizationBarrier_10_io_x_ppn = 20'h0; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@178025.4]
  assign pma_checker_OptimizationBarrier_10_io_x_u = 1'h0; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@178025.4]
  assign pma_checker_OptimizationBarrier_10_io_x_ae = 1'h0; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@178025.4]
  assign pma_checker_OptimizationBarrier_10_io_x_sw = 1'h0; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@178025.4]
  assign pma_checker_OptimizationBarrier_10_io_x_sx = 1'h0; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@178025.4]
  assign pma_checker_OptimizationBarrier_10_io_x_sr = 1'h0; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@178025.4]
  assign pma_checker_OptimizationBarrier_10_io_x_pw = 1'h0; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@178025.4]
  assign pma_checker_OptimizationBarrier_10_io_x_px = 1'h0; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@178025.4]
  assign pma_checker_OptimizationBarrier_10_io_x_pr = 1'h0; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@178025.4]
  assign pma_checker_OptimizationBarrier_10_io_x_ppp = 1'h0; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@178025.4]
  assign pma_checker_OptimizationBarrier_10_io_x_pal = 1'h0; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@178025.4]
  assign pma_checker_OptimizationBarrier_10_io_x_paa = 1'h0; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@178025.4]
  assign pma_checker_OptimizationBarrier_10_io_x_eff = 1'h0; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@178025.4]
  assign pma_checker_OptimizationBarrier_10_io_x_c = 1'h0; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@178025.4]
  assign pma_checker_OptimizationBarrier_11_io_x_ppn = 20'h0; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@178074.4]
  assign pma_checker_OptimizationBarrier_11_io_x_u = 1'h0; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@178074.4]
  assign pma_checker_OptimizationBarrier_11_io_x_ae = 1'h0; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@178074.4]
  assign pma_checker_OptimizationBarrier_11_io_x_sw = 1'h0; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@178074.4]
  assign pma_checker_OptimizationBarrier_11_io_x_sx = 1'h0; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@178074.4]
  assign pma_checker_OptimizationBarrier_11_io_x_sr = 1'h0; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@178074.4]
  assign pma_checker_OptimizationBarrier_11_io_x_pw = 1'h0; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@178074.4]
  assign pma_checker_OptimizationBarrier_11_io_x_px = 1'h0; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@178074.4]
  assign pma_checker_OptimizationBarrier_11_io_x_pr = 1'h0; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@178074.4]
  assign pma_checker_OptimizationBarrier_11_io_x_ppp = 1'h0; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@178074.4]
  assign pma_checker_OptimizationBarrier_11_io_x_pal = 1'h0; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@178074.4]
  assign pma_checker_OptimizationBarrier_11_io_x_paa = 1'h0; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@178074.4]
  assign pma_checker_OptimizationBarrier_11_io_x_eff = 1'h0; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@178074.4]
  assign pma_checker_OptimizationBarrier_11_io_x_c = 1'h0; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@178074.4]
  assign pma_checker_OptimizationBarrier_12_io_x_ppn = 20'h0; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@178123.4]
  assign pma_checker_OptimizationBarrier_12_io_x_u = 1'h0; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@178123.4]
  assign pma_checker_OptimizationBarrier_12_io_x_ae = 1'h0; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@178123.4]
  assign pma_checker_OptimizationBarrier_12_io_x_sw = 1'h0; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@178123.4]
  assign pma_checker_OptimizationBarrier_12_io_x_sx = 1'h0; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@178123.4]
  assign pma_checker_OptimizationBarrier_12_io_x_sr = 1'h0; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@178123.4]
  assign pma_checker_OptimizationBarrier_12_io_x_pw = 1'h0; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@178123.4]
  assign pma_checker_OptimizationBarrier_12_io_x_px = 1'h0; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@178123.4]
  assign pma_checker_OptimizationBarrier_12_io_x_pr = 1'h0; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@178123.4]
  assign pma_checker_OptimizationBarrier_12_io_x_ppp = 1'h0; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@178123.4]
  assign pma_checker_OptimizationBarrier_12_io_x_pal = 1'h0; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@178123.4]
  assign pma_checker_OptimizationBarrier_12_io_x_paa = 1'h0; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@178123.4]
  assign pma_checker_OptimizationBarrier_12_io_x_eff = 1'h0; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@178123.4]
  assign pma_checker_OptimizationBarrier_12_io_x_c = 1'h0; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@178123.4]
  assign pma_checker_OptimizationBarrier_13_io_x_ppn = 20'h0; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@178172.4]
  assign pma_checker_OptimizationBarrier_13_io_x_u = 1'h0; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@178172.4]
  assign pma_checker_OptimizationBarrier_13_io_x_ae = 1'h0; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@178172.4]
  assign pma_checker_OptimizationBarrier_13_io_x_sw = 1'h0; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@178172.4]
  assign pma_checker_OptimizationBarrier_13_io_x_sx = 1'h0; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@178172.4]
  assign pma_checker_OptimizationBarrier_13_io_x_sr = 1'h0; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@178172.4]
  assign pma_checker_OptimizationBarrier_13_io_x_pw = 1'h0; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@178172.4]
  assign pma_checker_OptimizationBarrier_13_io_x_px = 1'h0; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@178172.4]
  assign pma_checker_OptimizationBarrier_13_io_x_pr = 1'h0; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@178172.4]
  assign pma_checker_OptimizationBarrier_13_io_x_ppp = 1'h0; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@178172.4]
  assign pma_checker_OptimizationBarrier_13_io_x_pal = 1'h0; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@178172.4]
  assign pma_checker_OptimizationBarrier_13_io_x_paa = 1'h0; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@178172.4]
  assign pma_checker_OptimizationBarrier_13_io_x_eff = 1'h0; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@178172.4]
  assign pma_checker_OptimizationBarrier_13_io_x_c = 1'h0; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@178172.4]
  assign pma_checker_OptimizationBarrier_14_io_x_ppn = 20'h0; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@178653.4]
  assign pma_checker_OptimizationBarrier_14_io_x_u = 1'h0; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@178653.4]
  assign pma_checker_OptimizationBarrier_14_io_x_ae = 1'h0; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@178653.4]
  assign pma_checker_OptimizationBarrier_14_io_x_sw = 1'h0; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@178653.4]
  assign pma_checker_OptimizationBarrier_14_io_x_sx = 1'h0; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@178653.4]
  assign pma_checker_OptimizationBarrier_14_io_x_sr = 1'h0; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@178653.4]
  assign pma_checker_OptimizationBarrier_14_io_x_pw = 1'h0; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@178653.4]
  assign pma_checker_OptimizationBarrier_14_io_x_px = 1'h0; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@178653.4]
  assign pma_checker_OptimizationBarrier_14_io_x_pr = 1'h0; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@178653.4]
  assign pma_checker_OptimizationBarrier_14_io_x_ppp = 1'h0; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@178653.4]
  assign pma_checker_OptimizationBarrier_14_io_x_pal = 1'h0; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@178653.4]
  assign pma_checker_OptimizationBarrier_14_io_x_paa = 1'h0; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@178653.4]
  assign pma_checker_OptimizationBarrier_14_io_x_eff = 1'h0; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@178653.4]
  assign pma_checker_OptimizationBarrier_14_io_x_c = 1'h0; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@178653.4]
  assign pma_checker_OptimizationBarrier_15_io_x_ppn = 20'h0; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@178696.4]
  assign pma_checker_OptimizationBarrier_15_io_x_u = 1'h0; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@178696.4]
  assign pma_checker_OptimizationBarrier_15_io_x_ae = 1'h0; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@178696.4]
  assign pma_checker_OptimizationBarrier_15_io_x_sw = 1'h0; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@178696.4]
  assign pma_checker_OptimizationBarrier_15_io_x_sx = 1'h0; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@178696.4]
  assign pma_checker_OptimizationBarrier_15_io_x_sr = 1'h0; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@178696.4]
  assign pma_checker_OptimizationBarrier_15_io_x_pw = 1'h0; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@178696.4]
  assign pma_checker_OptimizationBarrier_15_io_x_px = 1'h0; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@178696.4]
  assign pma_checker_OptimizationBarrier_15_io_x_pr = 1'h0; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@178696.4]
  assign pma_checker_OptimizationBarrier_15_io_x_ppp = 1'h0; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@178696.4]
  assign pma_checker_OptimizationBarrier_15_io_x_pal = 1'h0; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@178696.4]
  assign pma_checker_OptimizationBarrier_15_io_x_paa = 1'h0; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@178696.4]
  assign pma_checker_OptimizationBarrier_15_io_x_eff = 1'h0; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@178696.4]
  assign pma_checker_OptimizationBarrier_15_io_x_c = 1'h0; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@178696.4]
  assign pma_checker_OptimizationBarrier_16_io_x_ppn = 20'h0; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@178739.4]
  assign pma_checker_OptimizationBarrier_16_io_x_u = 1'h0; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@178739.4]
  assign pma_checker_OptimizationBarrier_16_io_x_ae = 1'h0; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@178739.4]
  assign pma_checker_OptimizationBarrier_16_io_x_sw = 1'h0; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@178739.4]
  assign pma_checker_OptimizationBarrier_16_io_x_sx = 1'h0; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@178739.4]
  assign pma_checker_OptimizationBarrier_16_io_x_sr = 1'h0; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@178739.4]
  assign pma_checker_OptimizationBarrier_16_io_x_pw = 1'h0; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@178739.4]
  assign pma_checker_OptimizationBarrier_16_io_x_px = 1'h0; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@178739.4]
  assign pma_checker_OptimizationBarrier_16_io_x_pr = 1'h0; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@178739.4]
  assign pma_checker_OptimizationBarrier_16_io_x_ppp = 1'h0; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@178739.4]
  assign pma_checker_OptimizationBarrier_16_io_x_pal = 1'h0; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@178739.4]
  assign pma_checker_OptimizationBarrier_16_io_x_paa = 1'h0; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@178739.4]
  assign pma_checker_OptimizationBarrier_16_io_x_eff = 1'h0; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@178739.4]
  assign pma_checker_OptimizationBarrier_16_io_x_c = 1'h0; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@178739.4]
  assign pma_checker_OptimizationBarrier_17_io_x_ppn = 20'h0; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@178782.4]
  assign pma_checker_OptimizationBarrier_17_io_x_u = 1'h0; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@178782.4]
  assign pma_checker_OptimizationBarrier_17_io_x_ae = 1'h0; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@178782.4]
  assign pma_checker_OptimizationBarrier_17_io_x_sw = 1'h0; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@178782.4]
  assign pma_checker_OptimizationBarrier_17_io_x_sx = 1'h0; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@178782.4]
  assign pma_checker_OptimizationBarrier_17_io_x_sr = 1'h0; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@178782.4]
  assign pma_checker_OptimizationBarrier_17_io_x_pw = 1'h0; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@178782.4]
  assign pma_checker_OptimizationBarrier_17_io_x_px = 1'h0; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@178782.4]
  assign pma_checker_OptimizationBarrier_17_io_x_pr = 1'h0; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@178782.4]
  assign pma_checker_OptimizationBarrier_17_io_x_ppp = 1'h0; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@178782.4]
  assign pma_checker_OptimizationBarrier_17_io_x_pal = 1'h0; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@178782.4]
  assign pma_checker_OptimizationBarrier_17_io_x_paa = 1'h0; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@178782.4]
  assign pma_checker_OptimizationBarrier_17_io_x_eff = 1'h0; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@178782.4]
  assign pma_checker_OptimizationBarrier_17_io_x_c = 1'h0; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@178782.4]
  assign pma_checker_OptimizationBarrier_18_io_x_ppn = 20'h0; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@178825.4]
  assign pma_checker_OptimizationBarrier_18_io_x_u = 1'h0; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@178825.4]
  assign pma_checker_OptimizationBarrier_18_io_x_ae = 1'h0; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@178825.4]
  assign pma_checker_OptimizationBarrier_18_io_x_sw = 1'h0; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@178825.4]
  assign pma_checker_OptimizationBarrier_18_io_x_sx = 1'h0; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@178825.4]
  assign pma_checker_OptimizationBarrier_18_io_x_sr = 1'h0; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@178825.4]
  assign pma_checker_OptimizationBarrier_18_io_x_pw = 1'h0; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@178825.4]
  assign pma_checker_OptimizationBarrier_18_io_x_px = 1'h0; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@178825.4]
  assign pma_checker_OptimizationBarrier_18_io_x_pr = 1'h0; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@178825.4]
  assign pma_checker_OptimizationBarrier_18_io_x_ppp = 1'h0; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@178825.4]
  assign pma_checker_OptimizationBarrier_18_io_x_pal = 1'h0; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@178825.4]
  assign pma_checker_OptimizationBarrier_18_io_x_paa = 1'h0; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@178825.4]
  assign pma_checker_OptimizationBarrier_18_io_x_eff = 1'h0; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@178825.4]
  assign pma_checker_OptimizationBarrier_18_io_x_c = 1'h0; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@178825.4]
  assign pma_checker_OptimizationBarrier_19_io_x_ppn = 20'h0; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@178868.4]
  assign pma_checker_OptimizationBarrier_19_io_x_u = 1'h0; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@178868.4]
  assign pma_checker_OptimizationBarrier_19_io_x_ae = 1'h0; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@178868.4]
  assign pma_checker_OptimizationBarrier_19_io_x_sw = 1'h0; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@178868.4]
  assign pma_checker_OptimizationBarrier_19_io_x_sx = 1'h0; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@178868.4]
  assign pma_checker_OptimizationBarrier_19_io_x_sr = 1'h0; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@178868.4]
  assign pma_checker_OptimizationBarrier_19_io_x_pw = 1'h0; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@178868.4]
  assign pma_checker_OptimizationBarrier_19_io_x_px = 1'h0; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@178868.4]
  assign pma_checker_OptimizationBarrier_19_io_x_pr = 1'h0; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@178868.4]
  assign pma_checker_OptimizationBarrier_19_io_x_ppp = 1'h0; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@178868.4]
  assign pma_checker_OptimizationBarrier_19_io_x_pal = 1'h0; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@178868.4]
  assign pma_checker_OptimizationBarrier_19_io_x_paa = 1'h0; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@178868.4]
  assign pma_checker_OptimizationBarrier_19_io_x_eff = 1'h0; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@178868.4]
  assign pma_checker_OptimizationBarrier_19_io_x_c = 1'h0; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@178868.4]
  assign pma_checker_OptimizationBarrier_20_io_x_ppn = 20'h0; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@178911.4]
  assign pma_checker_OptimizationBarrier_20_io_x_u = 1'h0; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@178911.4]
  assign pma_checker_OptimizationBarrier_20_io_x_ae = 1'h0; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@178911.4]
  assign pma_checker_OptimizationBarrier_20_io_x_sw = 1'h0; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@178911.4]
  assign pma_checker_OptimizationBarrier_20_io_x_sx = 1'h0; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@178911.4]
  assign pma_checker_OptimizationBarrier_20_io_x_sr = 1'h0; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@178911.4]
  assign pma_checker_OptimizationBarrier_20_io_x_pw = 1'h0; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@178911.4]
  assign pma_checker_OptimizationBarrier_20_io_x_px = 1'h0; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@178911.4]
  assign pma_checker_OptimizationBarrier_20_io_x_pr = 1'h0; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@178911.4]
  assign pma_checker_OptimizationBarrier_20_io_x_ppp = 1'h0; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@178911.4]
  assign pma_checker_OptimizationBarrier_20_io_x_pal = 1'h0; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@178911.4]
  assign pma_checker_OptimizationBarrier_20_io_x_paa = 1'h0; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@178911.4]
  assign pma_checker_OptimizationBarrier_20_io_x_eff = 1'h0; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@178911.4]
  assign pma_checker_OptimizationBarrier_20_io_x_c = 1'h0; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@178911.4]
  assign pma_checker_OptimizationBarrier_21_io_x_ppn = 20'h0; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@178954.4]
  assign pma_checker_OptimizationBarrier_21_io_x_u = 1'h0; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@178954.4]
  assign pma_checker_OptimizationBarrier_21_io_x_ae = 1'h0; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@178954.4]
  assign pma_checker_OptimizationBarrier_21_io_x_sw = 1'h0; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@178954.4]
  assign pma_checker_OptimizationBarrier_21_io_x_sx = 1'h0; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@178954.4]
  assign pma_checker_OptimizationBarrier_21_io_x_sr = 1'h0; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@178954.4]
  assign pma_checker_OptimizationBarrier_21_io_x_pw = 1'h0; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@178954.4]
  assign pma_checker_OptimizationBarrier_21_io_x_px = 1'h0; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@178954.4]
  assign pma_checker_OptimizationBarrier_21_io_x_pr = 1'h0; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@178954.4]
  assign pma_checker_OptimizationBarrier_21_io_x_ppp = 1'h0; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@178954.4]
  assign pma_checker_OptimizationBarrier_21_io_x_pal = 1'h0; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@178954.4]
  assign pma_checker_OptimizationBarrier_21_io_x_paa = 1'h0; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@178954.4]
  assign pma_checker_OptimizationBarrier_21_io_x_eff = 1'h0; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@178954.4]
  assign pma_checker_OptimizationBarrier_21_io_x_c = 1'h0; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@178954.4]
  assign pma_checker_OptimizationBarrier_22_io_x_ppn = 20'h0; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@178996.4]
  assign pma_checker_OptimizationBarrier_22_io_x_u = 1'h0; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@178996.4]
  assign pma_checker_OptimizationBarrier_22_io_x_ae = 1'h0; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@178996.4]
  assign pma_checker_OptimizationBarrier_22_io_x_sw = 1'h0; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@178996.4]
  assign pma_checker_OptimizationBarrier_22_io_x_sx = 1'h0; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@178996.4]
  assign pma_checker_OptimizationBarrier_22_io_x_sr = 1'h0; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@178996.4]
  assign pma_checker_OptimizationBarrier_22_io_x_pw = 1'h0; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@178996.4]
  assign pma_checker_OptimizationBarrier_22_io_x_px = 1'h0; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@178996.4]
  assign pma_checker_OptimizationBarrier_22_io_x_pr = 1'h0; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@178996.4]
  assign pma_checker_OptimizationBarrier_22_io_x_ppp = 1'h0; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@178996.4]
  assign pma_checker_OptimizationBarrier_22_io_x_pal = 1'h0; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@178996.4]
  assign pma_checker_OptimizationBarrier_22_io_x_paa = 1'h0; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@178996.4]
  assign pma_checker_OptimizationBarrier_22_io_x_eff = 1'h0; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@178996.4]
  assign pma_checker_OptimizationBarrier_22_io_x_c = 1'h0; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@178996.4]
  assign pma_checker_OptimizationBarrier_23_io_x_ppn = 20'h0; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@179038.4]
  assign pma_checker_OptimizationBarrier_23_io_x_u = 1'h0; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@179038.4]
  assign pma_checker_OptimizationBarrier_23_io_x_ae = 1'h0; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@179038.4]
  assign pma_checker_OptimizationBarrier_23_io_x_sw = 1'h0; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@179038.4]
  assign pma_checker_OptimizationBarrier_23_io_x_sx = 1'h0; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@179038.4]
  assign pma_checker_OptimizationBarrier_23_io_x_sr = 1'h0; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@179038.4]
  assign pma_checker_OptimizationBarrier_23_io_x_pw = 1'h0; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@179038.4]
  assign pma_checker_OptimizationBarrier_23_io_x_px = 1'h0; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@179038.4]
  assign pma_checker_OptimizationBarrier_23_io_x_pr = 1'h0; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@179038.4]
  assign pma_checker_OptimizationBarrier_23_io_x_ppp = 1'h0; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@179038.4]
  assign pma_checker_OptimizationBarrier_23_io_x_pal = 1'h0; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@179038.4]
  assign pma_checker_OptimizationBarrier_23_io_x_paa = 1'h0; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@179038.4]
  assign pma_checker_OptimizationBarrier_23_io_x_eff = 1'h0; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@179038.4]
  assign pma_checker_OptimizationBarrier_23_io_x_c = 1'h0; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@179038.4]
  assign pma_checker_OptimizationBarrier_24_io_x_ppn = 20'h0; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@179080.4]
  assign pma_checker_OptimizationBarrier_24_io_x_u = 1'h0; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@179080.4]
  assign pma_checker_OptimizationBarrier_24_io_x_ae = 1'h0; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@179080.4]
  assign pma_checker_OptimizationBarrier_24_io_x_sw = 1'h0; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@179080.4]
  assign pma_checker_OptimizationBarrier_24_io_x_sx = 1'h0; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@179080.4]
  assign pma_checker_OptimizationBarrier_24_io_x_sr = 1'h0; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@179080.4]
  assign pma_checker_OptimizationBarrier_24_io_x_pw = 1'h0; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@179080.4]
  assign pma_checker_OptimizationBarrier_24_io_x_px = 1'h0; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@179080.4]
  assign pma_checker_OptimizationBarrier_24_io_x_pr = 1'h0; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@179080.4]
  assign pma_checker_OptimizationBarrier_24_io_x_ppp = 1'h0; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@179080.4]
  assign pma_checker_OptimizationBarrier_24_io_x_pal = 1'h0; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@179080.4]
  assign pma_checker_OptimizationBarrier_24_io_x_paa = 1'h0; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@179080.4]
  assign pma_checker_OptimizationBarrier_24_io_x_eff = 1'h0; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@179080.4]
  assign pma_checker_OptimizationBarrier_24_io_x_c = 1'h0; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@179080.4]
  assign pma_checker_OptimizationBarrier_25_io_x_ppn = 20'h0; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@179122.4]
  assign pma_checker_OptimizationBarrier_25_io_x_u = 1'h0; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@179122.4]
  assign pma_checker_OptimizationBarrier_25_io_x_ae = 1'h0; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@179122.4]
  assign pma_checker_OptimizationBarrier_25_io_x_sw = 1'h0; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@179122.4]
  assign pma_checker_OptimizationBarrier_25_io_x_sx = 1'h0; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@179122.4]
  assign pma_checker_OptimizationBarrier_25_io_x_sr = 1'h0; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@179122.4]
  assign pma_checker_OptimizationBarrier_25_io_x_pw = 1'h0; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@179122.4]
  assign pma_checker_OptimizationBarrier_25_io_x_px = 1'h0; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@179122.4]
  assign pma_checker_OptimizationBarrier_25_io_x_pr = 1'h0; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@179122.4]
  assign pma_checker_OptimizationBarrier_25_io_x_ppp = 1'h0; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@179122.4]
  assign pma_checker_OptimizationBarrier_25_io_x_pal = 1'h0; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@179122.4]
  assign pma_checker_OptimizationBarrier_25_io_x_paa = 1'h0; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@179122.4]
  assign pma_checker_OptimizationBarrier_25_io_x_eff = 1'h0; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@179122.4]
  assign pma_checker_OptimizationBarrier_25_io_x_c = 1'h0; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@179122.4]
  assign pma_checker_OptimizationBarrier_26_io_x_ppn = 20'h0; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@179164.4]
  assign pma_checker_OptimizationBarrier_26_io_x_u = 1'h0; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@179164.4]
  assign pma_checker_OptimizationBarrier_26_io_x_ae = 1'h0; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@179164.4]
  assign pma_checker_OptimizationBarrier_26_io_x_sw = 1'h0; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@179164.4]
  assign pma_checker_OptimizationBarrier_26_io_x_sx = 1'h0; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@179164.4]
  assign pma_checker_OptimizationBarrier_26_io_x_sr = 1'h0; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@179164.4]
  assign pma_checker_OptimizationBarrier_26_io_x_pw = 1'h0; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@179164.4]
  assign pma_checker_OptimizationBarrier_26_io_x_px = 1'h0; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@179164.4]
  assign pma_checker_OptimizationBarrier_26_io_x_pr = 1'h0; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@179164.4]
  assign pma_checker_OptimizationBarrier_26_io_x_ppp = 1'h0; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@179164.4]
  assign pma_checker_OptimizationBarrier_26_io_x_pal = 1'h0; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@179164.4]
  assign pma_checker_OptimizationBarrier_26_io_x_paa = 1'h0; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@179164.4]
  assign pma_checker_OptimizationBarrier_26_io_x_eff = 1'h0; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@179164.4]
  assign pma_checker_OptimizationBarrier_26_io_x_c = 1'h0; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@179164.4]
  assign pma_checker_OptimizationBarrier_27_io_x_ppn = 20'h0; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@179207.4]
  assign pma_checker_OptimizationBarrier_27_io_x_u = 1'h0; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@179207.4]
  assign pma_checker_OptimizationBarrier_27_io_x_ae = 1'h0; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@179207.4]
  assign pma_checker_OptimizationBarrier_27_io_x_sw = 1'h0; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@179207.4]
  assign pma_checker_OptimizationBarrier_27_io_x_sx = 1'h0; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@179207.4]
  assign pma_checker_OptimizationBarrier_27_io_x_sr = 1'h0; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@179207.4]
  assign pma_checker_OptimizationBarrier_27_io_x_pw = 1'h0; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@179207.4]
  assign pma_checker_OptimizationBarrier_27_io_x_px = 1'h0; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@179207.4]
  assign pma_checker_OptimizationBarrier_27_io_x_pr = 1'h0; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@179207.4]
  assign pma_checker_OptimizationBarrier_27_io_x_ppp = 1'h0; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@179207.4]
  assign pma_checker_OptimizationBarrier_27_io_x_pal = 1'h0; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@179207.4]
  assign pma_checker_OptimizationBarrier_27_io_x_paa = 1'h0; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@179207.4]
  assign pma_checker_OptimizationBarrier_27_io_x_eff = 1'h0; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@179207.4]
  assign pma_checker_OptimizationBarrier_27_io_x_c = 1'h0; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@179207.4]
  assign pma_checker_OptimizationBarrier_28_io_x_ppn = 20'h0; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@179250.4]
  assign pma_checker_OptimizationBarrier_28_io_x_u = 1'h0; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@179250.4]
  assign pma_checker_OptimizationBarrier_28_io_x_ae = 1'h0; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@179250.4]
  assign pma_checker_OptimizationBarrier_28_io_x_sw = 1'h0; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@179250.4]
  assign pma_checker_OptimizationBarrier_28_io_x_sx = 1'h0; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@179250.4]
  assign pma_checker_OptimizationBarrier_28_io_x_sr = 1'h0; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@179250.4]
  assign pma_checker_OptimizationBarrier_28_io_x_pw = 1'h0; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@179250.4]
  assign pma_checker_OptimizationBarrier_28_io_x_px = 1'h0; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@179250.4]
  assign pma_checker_OptimizationBarrier_28_io_x_pr = 1'h0; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@179250.4]
  assign pma_checker_OptimizationBarrier_28_io_x_ppp = 1'h0; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@179250.4]
  assign pma_checker_OptimizationBarrier_28_io_x_pal = 1'h0; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@179250.4]
  assign pma_checker_OptimizationBarrier_28_io_x_paa = 1'h0; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@179250.4]
  assign pma_checker_OptimizationBarrier_28_io_x_eff = 1'h0; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@179250.4]
  assign pma_checker_OptimizationBarrier_28_io_x_c = 1'h0; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@179250.4]
  assign pma_checker_OptimizationBarrier_29_io_x_ppn = 20'h0; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@179293.4]
  assign pma_checker_OptimizationBarrier_29_io_x_u = 1'h0; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@179293.4]
  assign pma_checker_OptimizationBarrier_29_io_x_ae = 1'h0; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@179293.4]
  assign pma_checker_OptimizationBarrier_29_io_x_sw = 1'h0; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@179293.4]
  assign pma_checker_OptimizationBarrier_29_io_x_sx = 1'h0; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@179293.4]
  assign pma_checker_OptimizationBarrier_29_io_x_sr = 1'h0; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@179293.4]
  assign pma_checker_OptimizationBarrier_29_io_x_pw = 1'h0; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@179293.4]
  assign pma_checker_OptimizationBarrier_29_io_x_px = 1'h0; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@179293.4]
  assign pma_checker_OptimizationBarrier_29_io_x_pr = 1'h0; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@179293.4]
  assign pma_checker_OptimizationBarrier_29_io_x_ppp = 1'h0; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@179293.4]
  assign pma_checker_OptimizationBarrier_29_io_x_pal = 1'h0; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@179293.4]
  assign pma_checker_OptimizationBarrier_29_io_x_paa = 1'h0; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@179293.4]
  assign pma_checker_OptimizationBarrier_29_io_x_eff = 1'h0; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@179293.4]
  assign pma_checker_OptimizationBarrier_29_io_x_c = 1'h0; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@179293.4]
  assign pma_checker_OptimizationBarrier_30_io_x_ppn = 20'h0; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@179336.4]
  assign pma_checker_OptimizationBarrier_30_io_x_u = 1'h0; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@179336.4]
  assign pma_checker_OptimizationBarrier_30_io_x_ae = 1'h0; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@179336.4]
  assign pma_checker_OptimizationBarrier_30_io_x_sw = 1'h0; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@179336.4]
  assign pma_checker_OptimizationBarrier_30_io_x_sx = 1'h0; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@179336.4]
  assign pma_checker_OptimizationBarrier_30_io_x_sr = 1'h0; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@179336.4]
  assign pma_checker_OptimizationBarrier_30_io_x_pw = 1'h0; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@179336.4]
  assign pma_checker_OptimizationBarrier_30_io_x_px = 1'h0; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@179336.4]
  assign pma_checker_OptimizationBarrier_30_io_x_pr = 1'h0; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@179336.4]
  assign pma_checker_OptimizationBarrier_30_io_x_ppp = 1'h0; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@179336.4]
  assign pma_checker_OptimizationBarrier_30_io_x_pal = 1'h0; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@179336.4]
  assign pma_checker_OptimizationBarrier_30_io_x_paa = 1'h0; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@179336.4]
  assign pma_checker_OptimizationBarrier_30_io_x_eff = 1'h0; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@179336.4]
  assign pma_checker_OptimizationBarrier_30_io_x_c = 1'h0; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@179336.4]
  assign pma_checker_OptimizationBarrier_31_io_x_ppn = 20'h0; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@179379.4]
  assign pma_checker_OptimizationBarrier_31_io_x_u = 1'h0; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@179379.4]
  assign pma_checker_OptimizationBarrier_31_io_x_ae = 1'h0; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@179379.4]
  assign pma_checker_OptimizationBarrier_31_io_x_sw = 1'h0; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@179379.4]
  assign pma_checker_OptimizationBarrier_31_io_x_sx = 1'h0; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@179379.4]
  assign pma_checker_OptimizationBarrier_31_io_x_sr = 1'h0; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@179379.4]
  assign pma_checker_OptimizationBarrier_31_io_x_pw = 1'h0; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@179379.4]
  assign pma_checker_OptimizationBarrier_31_io_x_px = 1'h0; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@179379.4]
  assign pma_checker_OptimizationBarrier_31_io_x_pr = 1'h0; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@179379.4]
  assign pma_checker_OptimizationBarrier_31_io_x_ppp = 1'h0; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@179379.4]
  assign pma_checker_OptimizationBarrier_31_io_x_pal = 1'h0; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@179379.4]
  assign pma_checker_OptimizationBarrier_31_io_x_paa = 1'h0; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@179379.4]
  assign pma_checker_OptimizationBarrier_31_io_x_eff = 1'h0; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@179379.4]
  assign pma_checker_OptimizationBarrier_31_io_x_c = 1'h0; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@179379.4]
  assign pma_checker_OptimizationBarrier_32_io_x_ppn = 20'h0; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@179422.4]
  assign pma_checker_OptimizationBarrier_32_io_x_u = 1'h0; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@179422.4]
  assign pma_checker_OptimizationBarrier_32_io_x_ae = 1'h0; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@179422.4]
  assign pma_checker_OptimizationBarrier_32_io_x_sw = 1'h0; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@179422.4]
  assign pma_checker_OptimizationBarrier_32_io_x_sx = 1'h0; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@179422.4]
  assign pma_checker_OptimizationBarrier_32_io_x_sr = 1'h0; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@179422.4]
  assign pma_checker_OptimizationBarrier_32_io_x_pw = 1'h0; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@179422.4]
  assign pma_checker_OptimizationBarrier_32_io_x_px = 1'h0; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@179422.4]
  assign pma_checker_OptimizationBarrier_32_io_x_pr = 1'h0; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@179422.4]
  assign pma_checker_OptimizationBarrier_32_io_x_ppp = 1'h0; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@179422.4]
  assign pma_checker_OptimizationBarrier_32_io_x_pal = 1'h0; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@179422.4]
  assign pma_checker_OptimizationBarrier_32_io_x_paa = 1'h0; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@179422.4]
  assign pma_checker_OptimizationBarrier_32_io_x_eff = 1'h0; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@179422.4]
  assign pma_checker_OptimizationBarrier_32_io_x_c = 1'h0; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@179422.4]
  assign pma_checker_OptimizationBarrier_33_io_x_ppn = 20'h0; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@179465.4]
  assign pma_checker_OptimizationBarrier_33_io_x_u = 1'h0; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@179465.4]
  assign pma_checker_OptimizationBarrier_33_io_x_ae = 1'h0; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@179465.4]
  assign pma_checker_OptimizationBarrier_33_io_x_sw = 1'h0; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@179465.4]
  assign pma_checker_OptimizationBarrier_33_io_x_sx = 1'h0; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@179465.4]
  assign pma_checker_OptimizationBarrier_33_io_x_sr = 1'h0; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@179465.4]
  assign pma_checker_OptimizationBarrier_33_io_x_pw = 1'h0; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@179465.4]
  assign pma_checker_OptimizationBarrier_33_io_x_px = 1'h0; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@179465.4]
  assign pma_checker_OptimizationBarrier_33_io_x_pr = 1'h0; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@179465.4]
  assign pma_checker_OptimizationBarrier_33_io_x_ppp = 1'h0; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@179465.4]
  assign pma_checker_OptimizationBarrier_33_io_x_pal = 1'h0; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@179465.4]
  assign pma_checker_OptimizationBarrier_33_io_x_paa = 1'h0; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@179465.4]
  assign pma_checker_OptimizationBarrier_33_io_x_eff = 1'h0; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@179465.4]
  assign pma_checker_OptimizationBarrier_33_io_x_c = 1'h0; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@179465.4]
  assign pma_checker_OptimizationBarrier_34_io_x_ppn = 20'h0; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@179508.4]
  assign pma_checker_OptimizationBarrier_34_io_x_u = 1'h0; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@179508.4]
  assign pma_checker_OptimizationBarrier_34_io_x_ae = 1'h0; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@179508.4]
  assign pma_checker_OptimizationBarrier_34_io_x_sw = 1'h0; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@179508.4]
  assign pma_checker_OptimizationBarrier_34_io_x_sx = 1'h0; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@179508.4]
  assign pma_checker_OptimizationBarrier_34_io_x_sr = 1'h0; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@179508.4]
  assign pma_checker_OptimizationBarrier_34_io_x_pw = 1'h0; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@179508.4]
  assign pma_checker_OptimizationBarrier_34_io_x_px = 1'h0; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@179508.4]
  assign pma_checker_OptimizationBarrier_34_io_x_pr = 1'h0; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@179508.4]
  assign pma_checker_OptimizationBarrier_34_io_x_ppp = 1'h0; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@179508.4]
  assign pma_checker_OptimizationBarrier_34_io_x_pal = 1'h0; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@179508.4]
  assign pma_checker_OptimizationBarrier_34_io_x_paa = 1'h0; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@179508.4]
  assign pma_checker_OptimizationBarrier_34_io_x_eff = 1'h0; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@179508.4]
  assign pma_checker_OptimizationBarrier_34_io_x_c = 1'h0; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@179508.4]
  assign pma_checker_OptimizationBarrier_35_io_x_ppn = 20'h0; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@179550.4]
  assign pma_checker_OptimizationBarrier_35_io_x_u = 1'h0; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@179550.4]
  assign pma_checker_OptimizationBarrier_35_io_x_ae = 1'h0; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@179550.4]
  assign pma_checker_OptimizationBarrier_35_io_x_sw = 1'h0; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@179550.4]
  assign pma_checker_OptimizationBarrier_35_io_x_sx = 1'h0; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@179550.4]
  assign pma_checker_OptimizationBarrier_35_io_x_sr = 1'h0; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@179550.4]
  assign pma_checker_OptimizationBarrier_35_io_x_pw = 1'h0; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@179550.4]
  assign pma_checker_OptimizationBarrier_35_io_x_px = 1'h0; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@179550.4]
  assign pma_checker_OptimizationBarrier_35_io_x_pr = 1'h0; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@179550.4]
  assign pma_checker_OptimizationBarrier_35_io_x_ppp = 1'h0; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@179550.4]
  assign pma_checker_OptimizationBarrier_35_io_x_pal = 1'h0; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@179550.4]
  assign pma_checker_OptimizationBarrier_35_io_x_paa = 1'h0; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@179550.4]
  assign pma_checker_OptimizationBarrier_35_io_x_eff = 1'h0; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@179550.4]
  assign pma_checker_OptimizationBarrier_35_io_x_c = 1'h0; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@179550.4]
  assign pma_checker_OptimizationBarrier_36_io_x_ppn = 20'h0; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@179592.4]
  assign pma_checker_OptimizationBarrier_36_io_x_u = 1'h0; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@179592.4]
  assign pma_checker_OptimizationBarrier_36_io_x_ae = 1'h0; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@179592.4]
  assign pma_checker_OptimizationBarrier_36_io_x_sw = 1'h0; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@179592.4]
  assign pma_checker_OptimizationBarrier_36_io_x_sx = 1'h0; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@179592.4]
  assign pma_checker_OptimizationBarrier_36_io_x_sr = 1'h0; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@179592.4]
  assign pma_checker_OptimizationBarrier_36_io_x_pw = 1'h0; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@179592.4]
  assign pma_checker_OptimizationBarrier_36_io_x_px = 1'h0; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@179592.4]
  assign pma_checker_OptimizationBarrier_36_io_x_pr = 1'h0; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@179592.4]
  assign pma_checker_OptimizationBarrier_36_io_x_ppp = 1'h0; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@179592.4]
  assign pma_checker_OptimizationBarrier_36_io_x_pal = 1'h0; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@179592.4]
  assign pma_checker_OptimizationBarrier_36_io_x_paa = 1'h0; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@179592.4]
  assign pma_checker_OptimizationBarrier_36_io_x_eff = 1'h0; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@179592.4]
  assign pma_checker_OptimizationBarrier_36_io_x_c = 1'h0; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@179592.4]
  assign pma_checker_OptimizationBarrier_37_io_x_ppn = 20'h0; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@179634.4]
  assign pma_checker_OptimizationBarrier_37_io_x_u = 1'h0; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@179634.4]
  assign pma_checker_OptimizationBarrier_37_io_x_ae = 1'h0; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@179634.4]
  assign pma_checker_OptimizationBarrier_37_io_x_sw = 1'h0; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@179634.4]
  assign pma_checker_OptimizationBarrier_37_io_x_sx = 1'h0; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@179634.4]
  assign pma_checker_OptimizationBarrier_37_io_x_sr = 1'h0; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@179634.4]
  assign pma_checker_OptimizationBarrier_37_io_x_pw = 1'h0; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@179634.4]
  assign pma_checker_OptimizationBarrier_37_io_x_px = 1'h0; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@179634.4]
  assign pma_checker_OptimizationBarrier_37_io_x_pr = 1'h0; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@179634.4]
  assign pma_checker_OptimizationBarrier_37_io_x_ppp = 1'h0; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@179634.4]
  assign pma_checker_OptimizationBarrier_37_io_x_pal = 1'h0; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@179634.4]
  assign pma_checker_OptimizationBarrier_37_io_x_paa = 1'h0; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@179634.4]
  assign pma_checker_OptimizationBarrier_37_io_x_eff = 1'h0; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@179634.4]
  assign pma_checker_OptimizationBarrier_37_io_x_c = 1'h0; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@179634.4]
  assign pma_checker_OptimizationBarrier_38_io_x_ppn = 20'h0; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@179676.4]
  assign pma_checker_OptimizationBarrier_38_io_x_u = 1'h0; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@179676.4]
  assign pma_checker_OptimizationBarrier_38_io_x_ae = 1'h0; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@179676.4]
  assign pma_checker_OptimizationBarrier_38_io_x_sw = 1'h0; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@179676.4]
  assign pma_checker_OptimizationBarrier_38_io_x_sx = 1'h0; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@179676.4]
  assign pma_checker_OptimizationBarrier_38_io_x_sr = 1'h0; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@179676.4]
  assign pma_checker_OptimizationBarrier_38_io_x_pw = 1'h0; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@179676.4]
  assign pma_checker_OptimizationBarrier_38_io_x_px = 1'h0; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@179676.4]
  assign pma_checker_OptimizationBarrier_38_io_x_pr = 1'h0; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@179676.4]
  assign pma_checker_OptimizationBarrier_38_io_x_ppp = 1'h0; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@179676.4]
  assign pma_checker_OptimizationBarrier_38_io_x_pal = 1'h0; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@179676.4]
  assign pma_checker_OptimizationBarrier_38_io_x_paa = 1'h0; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@179676.4]
  assign pma_checker_OptimizationBarrier_38_io_x_eff = 1'h0; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@179676.4]
  assign pma_checker_OptimizationBarrier_38_io_x_c = 1'h0; // @[package.scala 239:18:freechips.rocketchip.system.DefaultRV32Config.fir@179676.4]
  assign metaArb__GEN_1 = metaArb_io_in_6_valid ? metaArb_io_in_6_bits_data : metaArb_io_in_7_bits_data; // @[Arbiter.scala 126:27:freechips.rocketchip.system.DefaultRV32Config.fir@191722.4]
  assign metaArb__GEN_2 = metaArb_io_in_6_valid ? metaArb_io_in_6_bits_way_en : metaArb_io_in_7_bits_way_en; // @[Arbiter.scala 126:27:freechips.rocketchip.system.DefaultRV32Config.fir@191722.4]
  assign metaArb__GEN_3 = metaArb_io_in_6_valid ? metaArb_io_in_6_bits_idx : metaArb_io_in_7_bits_idx; // @[Arbiter.scala 126:27:freechips.rocketchip.system.DefaultRV32Config.fir@191722.4]
  assign metaArb__GEN_4 = metaArb_io_in_6_valid ? metaArb_io_in_6_bits_addr : metaArb_io_in_7_bits_addr; // @[Arbiter.scala 126:27:freechips.rocketchip.system.DefaultRV32Config.fir@191722.4]
  assign metaArb__GEN_13 = metaArb_io_in_4_valid ? metaArb_io_in_4_bits_data : metaArb__GEN_1; // @[Arbiter.scala 126:27:freechips.rocketchip.system.DefaultRV32Config.fir@191738.4]
  assign metaArb__GEN_14 = metaArb_io_in_4_valid ? metaArb_io_in_4_bits_way_en : metaArb__GEN_2; // @[Arbiter.scala 126:27:freechips.rocketchip.system.DefaultRV32Config.fir@191738.4]
  assign metaArb__GEN_15 = metaArb_io_in_4_valid ? metaArb_io_in_4_bits_idx : metaArb__GEN_3; // @[Arbiter.scala 126:27:freechips.rocketchip.system.DefaultRV32Config.fir@191738.4]
  assign metaArb__GEN_16 = metaArb_io_in_4_valid ? metaArb_io_in_4_bits_addr : metaArb__GEN_4; // @[Arbiter.scala 126:27:freechips.rocketchip.system.DefaultRV32Config.fir@191738.4]
  assign metaArb__GEN_19 = metaArb_io_in_3_valid ? metaArb_io_in_3_bits_data : metaArb__GEN_13; // @[Arbiter.scala 126:27:freechips.rocketchip.system.DefaultRV32Config.fir@191746.4]
  assign metaArb__GEN_20 = metaArb_io_in_3_valid ? metaArb_io_in_3_bits_way_en : metaArb__GEN_14; // @[Arbiter.scala 126:27:freechips.rocketchip.system.DefaultRV32Config.fir@191746.4]
  assign metaArb__GEN_21 = metaArb_io_in_3_valid ? metaArb_io_in_3_bits_idx : metaArb__GEN_15; // @[Arbiter.scala 126:27:freechips.rocketchip.system.DefaultRV32Config.fir@191746.4]
  assign metaArb__GEN_22 = metaArb_io_in_3_valid ? metaArb_io_in_3_bits_addr : metaArb__GEN_16; // @[Arbiter.scala 126:27:freechips.rocketchip.system.DefaultRV32Config.fir@191746.4]
  assign metaArb__GEN_23 = metaArb_io_in_3_valid | metaArb_io_in_4_valid; // @[Arbiter.scala 126:27:freechips.rocketchip.system.DefaultRV32Config.fir@191746.4]
  assign metaArb__GEN_25 = metaArb_io_in_2_valid ? metaArb_io_in_2_bits_data : metaArb__GEN_19; // @[Arbiter.scala 126:27:freechips.rocketchip.system.DefaultRV32Config.fir@191754.4]
  assign metaArb__GEN_26 = metaArb_io_in_2_valid ? metaArb_io_in_2_bits_way_en : metaArb__GEN_20; // @[Arbiter.scala 126:27:freechips.rocketchip.system.DefaultRV32Config.fir@191754.4]
  assign metaArb__GEN_27 = metaArb_io_in_2_valid ? metaArb_io_in_2_bits_idx : metaArb__GEN_21; // @[Arbiter.scala 126:27:freechips.rocketchip.system.DefaultRV32Config.fir@191754.4]
  assign metaArb__GEN_28 = metaArb_io_in_2_valid ? metaArb_io_in_2_bits_addr : metaArb__GEN_22; // @[Arbiter.scala 126:27:freechips.rocketchip.system.DefaultRV32Config.fir@191754.4]
  assign metaArb__GEN_29 = metaArb_io_in_2_valid | metaArb__GEN_23; // @[Arbiter.scala 126:27:freechips.rocketchip.system.DefaultRV32Config.fir@191754.4]
  assign metaArb__GEN_31 = metaArb_io_in_1_valid ? metaArb_io_in_1_bits_data : metaArb__GEN_25; // @[Arbiter.scala 126:27:freechips.rocketchip.system.DefaultRV32Config.fir@191762.4]
  assign metaArb__GEN_32 = metaArb_io_in_1_valid ? 4'h0 : metaArb__GEN_26; // @[Arbiter.scala 126:27:freechips.rocketchip.system.DefaultRV32Config.fir@191762.4]
  assign metaArb__GEN_33 = metaArb_io_in_1_valid ? metaArb_io_in_1_bits_idx : metaArb__GEN_27; // @[Arbiter.scala 126:27:freechips.rocketchip.system.DefaultRV32Config.fir@191762.4]
  assign metaArb__GEN_34 = metaArb_io_in_1_valid ? metaArb_io_in_1_bits_addr : metaArb__GEN_28; // @[Arbiter.scala 126:27:freechips.rocketchip.system.DefaultRV32Config.fir@191762.4]
  assign metaArb__GEN_35 = metaArb_io_in_1_valid | metaArb__GEN_29; // @[Arbiter.scala 126:27:freechips.rocketchip.system.DefaultRV32Config.fir@191762.4]
  assign metaArb__T = metaArb_io_in_0_valid | metaArb_io_in_1_valid; // @[Arbiter.scala 31:68:freechips.rocketchip.system.DefaultRV32Config.fir@191778.4]
  assign metaArb__T_1 = metaArb__T | metaArb_io_in_2_valid; // @[Arbiter.scala 31:68:freechips.rocketchip.system.DefaultRV32Config.fir@191779.4]
  assign metaArb__T_2 = metaArb__T_1 | metaArb_io_in_3_valid; // @[Arbiter.scala 31:68:freechips.rocketchip.system.DefaultRV32Config.fir@191780.4]
  assign metaArb__T_3 = metaArb__T_2 | metaArb_io_in_4_valid; // @[Arbiter.scala 31:68:freechips.rocketchip.system.DefaultRV32Config.fir@191781.4]
  assign metaArb__T_5 = metaArb__T_3 | metaArb_io_in_6_valid; // @[Arbiter.scala 31:68:freechips.rocketchip.system.DefaultRV32Config.fir@191783.4]
  assign metaArb_grant_7 = ~metaArb__T_5; // @[Arbiter.scala 31:78:freechips.rocketchip.system.DefaultRV32Config.fir@191790.4]
  assign metaArb__T_14 = ~metaArb_grant_7; // @[Arbiter.scala 135:19:freechips.rocketchip.system.DefaultRV32Config.fir@191807.4]
  assign metaArb_io_in_4_ready = ~metaArb__T_2; // @[Arbiter.scala 134:14:freechips.rocketchip.system.DefaultRV32Config.fir@191800.4]
  assign metaArb_io_in_6_ready = ~metaArb__T_3; // @[Arbiter.scala 134:14:freechips.rocketchip.system.DefaultRV32Config.fir@191804.4]
  assign metaArb_io_in_7_ready = ~metaArb__T_5; // @[Arbiter.scala 134:14:freechips.rocketchip.system.DefaultRV32Config.fir@191806.4]
  assign metaArb_io_out_valid = metaArb__T_14 | metaArb_io_in_7_valid; // @[Arbiter.scala 135:16:freechips.rocketchip.system.DefaultRV32Config.fir@191809.4]
  assign metaArb_io_out_bits_write = metaArb_io_in_0_valid | metaArb__GEN_35; // @[Arbiter.scala 124:15:freechips.rocketchip.system.DefaultRV32Config.fir@191721.4 Arbiter.scala 128:19:freechips.rocketchip.system.DefaultRV32Config.fir@191728.6 Arbiter.scala 128:19:freechips.rocketchip.system.DefaultRV32Config.fir@191736.6 Arbiter.scala 128:19:freechips.rocketchip.system.DefaultRV32Config.fir@191744.6 Arbiter.scala 128:19:freechips.rocketchip.system.DefaultRV32Config.fir@191752.6 Arbiter.scala 128:19:freechips.rocketchip.system.DefaultRV32Config.fir@191760.6 Arbiter.scala 128:19:freechips.rocketchip.system.DefaultRV32Config.fir@191768.6 Arbiter.scala 128:19:freechips.rocketchip.system.DefaultRV32Config.fir@191776.6]
  assign metaArb_io_out_bits_addr = metaArb_io_in_0_valid ? metaArb_io_in_0_bits_addr : metaArb__GEN_34; // @[Arbiter.scala 124:15:freechips.rocketchip.system.DefaultRV32Config.fir@191720.4 Arbiter.scala 128:19:freechips.rocketchip.system.DefaultRV32Config.fir@191727.6 Arbiter.scala 128:19:freechips.rocketchip.system.DefaultRV32Config.fir@191735.6 Arbiter.scala 128:19:freechips.rocketchip.system.DefaultRV32Config.fir@191743.6 Arbiter.scala 128:19:freechips.rocketchip.system.DefaultRV32Config.fir@191751.6 Arbiter.scala 128:19:freechips.rocketchip.system.DefaultRV32Config.fir@191759.6 Arbiter.scala 128:19:freechips.rocketchip.system.DefaultRV32Config.fir@191767.6 Arbiter.scala 128:19:freechips.rocketchip.system.DefaultRV32Config.fir@191775.6]
  assign metaArb_io_out_bits_idx = metaArb_io_in_0_valid ? metaArb_io_in_0_bits_idx : metaArb__GEN_33; // @[Arbiter.scala 124:15:freechips.rocketchip.system.DefaultRV32Config.fir@191719.4 Arbiter.scala 128:19:freechips.rocketchip.system.DefaultRV32Config.fir@191726.6 Arbiter.scala 128:19:freechips.rocketchip.system.DefaultRV32Config.fir@191734.6 Arbiter.scala 128:19:freechips.rocketchip.system.DefaultRV32Config.fir@191742.6 Arbiter.scala 128:19:freechips.rocketchip.system.DefaultRV32Config.fir@191750.6 Arbiter.scala 128:19:freechips.rocketchip.system.DefaultRV32Config.fir@191758.6 Arbiter.scala 128:19:freechips.rocketchip.system.DefaultRV32Config.fir@191766.6 Arbiter.scala 128:19:freechips.rocketchip.system.DefaultRV32Config.fir@191774.6]
  assign metaArb_io_out_bits_way_en = metaArb_io_in_0_valid ? 4'hf : metaArb__GEN_32; // @[Arbiter.scala 124:15:freechips.rocketchip.system.DefaultRV32Config.fir@191718.4 Arbiter.scala 128:19:freechips.rocketchip.system.DefaultRV32Config.fir@191725.6 Arbiter.scala 128:19:freechips.rocketchip.system.DefaultRV32Config.fir@191733.6 Arbiter.scala 128:19:freechips.rocketchip.system.DefaultRV32Config.fir@191741.6 Arbiter.scala 128:19:freechips.rocketchip.system.DefaultRV32Config.fir@191749.6 Arbiter.scala 128:19:freechips.rocketchip.system.DefaultRV32Config.fir@191757.6 Arbiter.scala 128:19:freechips.rocketchip.system.DefaultRV32Config.fir@191765.6 Arbiter.scala 128:19:freechips.rocketchip.system.DefaultRV32Config.fir@191773.6]
  assign metaArb_io_out_bits_data = metaArb_io_in_0_valid ? metaArb_io_in_0_bits_data : metaArb__GEN_31; // @[Arbiter.scala 124:15:freechips.rocketchip.system.DefaultRV32Config.fir@191717.4 Arbiter.scala 128:19:freechips.rocketchip.system.DefaultRV32Config.fir@191724.6 Arbiter.scala 128:19:freechips.rocketchip.system.DefaultRV32Config.fir@191732.6 Arbiter.scala 128:19:freechips.rocketchip.system.DefaultRV32Config.fir@191740.6 Arbiter.scala 128:19:freechips.rocketchip.system.DefaultRV32Config.fir@191748.6 Arbiter.scala 128:19:freechips.rocketchip.system.DefaultRV32Config.fir@191756.6 Arbiter.scala 128:19:freechips.rocketchip.system.DefaultRV32Config.fir@191764.6 Arbiter.scala 128:19:freechips.rocketchip.system.DefaultRV32Config.fir@191772.6]
  assign dataArb__GEN_4 = dataArb_io_in_2_valid ? dataArb_io_in_2_bits_wdata : dataArb_io_in_3_bits_wdata; // @[Arbiter.scala 126:27:freechips.rocketchip.system.DefaultRV32Config.fir@191975.4]
  assign dataArb__GEN_6 = dataArb_io_in_2_valid ? dataArb_io_in_2_bits_addr : dataArb_io_in_3_bits_addr; // @[Arbiter.scala 126:27:freechips.rocketchip.system.DefaultRV32Config.fir@191975.4]
  assign dataArb__GEN_8 = dataArb_io_in_1_valid ? dataArb_io_in_1_bits_way_en : 4'hf; // @[Arbiter.scala 126:27:freechips.rocketchip.system.DefaultRV32Config.fir@191984.4]
  assign dataArb__GEN_11 = dataArb_io_in_1_valid ? dataArb_io_in_1_bits_wdata : dataArb__GEN_4; // @[Arbiter.scala 126:27:freechips.rocketchip.system.DefaultRV32Config.fir@191984.4]
  assign dataArb__GEN_12 = dataArb_io_in_1_valid & dataArb_io_in_1_bits_write; // @[Arbiter.scala 126:27:freechips.rocketchip.system.DefaultRV32Config.fir@191984.4]
  assign dataArb__GEN_13 = dataArb_io_in_1_valid ? dataArb_io_in_1_bits_addr : dataArb__GEN_6; // @[Arbiter.scala 126:27:freechips.rocketchip.system.DefaultRV32Config.fir@191984.4]
  assign dataArb__T = dataArb_io_in_0_valid | dataArb_io_in_1_valid; // @[Arbiter.scala 31:68:freechips.rocketchip.system.DefaultRV32Config.fir@192002.4]
  assign dataArb__T_1 = dataArb__T | dataArb_io_in_2_valid; // @[Arbiter.scala 31:68:freechips.rocketchip.system.DefaultRV32Config.fir@192003.4]
  assign dataArb_grant_3 = ~dataArb__T_1; // @[Arbiter.scala 31:78:freechips.rocketchip.system.DefaultRV32Config.fir@192006.4]
  assign dataArb__T_6 = ~dataArb_grant_3; // @[Arbiter.scala 135:19:freechips.rocketchip.system.DefaultRV32Config.fir@192015.4]
  assign dataArb_io_in_1_ready = ~dataArb_io_in_0_valid; // @[Arbiter.scala 134:14:freechips.rocketchip.system.DefaultRV32Config.fir@192010.4]
  assign dataArb_io_in_2_ready = ~dataArb__T; // @[Arbiter.scala 134:14:freechips.rocketchip.system.DefaultRV32Config.fir@192012.4]
  assign dataArb_io_in_3_ready = ~dataArb__T_1; // @[Arbiter.scala 134:14:freechips.rocketchip.system.DefaultRV32Config.fir@192014.4]
  assign dataArb_io_out_valid = dataArb__T_6 | dataArb_io_in_3_valid; // @[Arbiter.scala 135:16:freechips.rocketchip.system.DefaultRV32Config.fir@192017.4]
  assign dataArb_io_out_bits_addr = dataArb_io_in_0_valid ? dataArb_io_in_0_bits_addr : dataArb__GEN_13; // @[Arbiter.scala 124:15:freechips.rocketchip.system.DefaultRV32Config.fir@191974.4 Arbiter.scala 128:19:freechips.rocketchip.system.DefaultRV32Config.fir@191982.6 Arbiter.scala 128:19:freechips.rocketchip.system.DefaultRV32Config.fir@191991.6 Arbiter.scala 128:19:freechips.rocketchip.system.DefaultRV32Config.fir@192000.6]
  assign dataArb_io_out_bits_write = dataArb_io_in_0_valid ? dataArb_io_in_0_bits_write : dataArb__GEN_12; // @[Arbiter.scala 124:15:freechips.rocketchip.system.DefaultRV32Config.fir@191973.4 Arbiter.scala 128:19:freechips.rocketchip.system.DefaultRV32Config.fir@191981.6 Arbiter.scala 128:19:freechips.rocketchip.system.DefaultRV32Config.fir@191990.6 Arbiter.scala 128:19:freechips.rocketchip.system.DefaultRV32Config.fir@191999.6]
  assign dataArb_io_out_bits_wdata = dataArb_io_in_0_valid ? dataArb_io_in_0_bits_wdata : dataArb__GEN_11; // @[Arbiter.scala 124:15:freechips.rocketchip.system.DefaultRV32Config.fir@191972.4 Arbiter.scala 128:19:freechips.rocketchip.system.DefaultRV32Config.fir@191980.6 Arbiter.scala 128:19:freechips.rocketchip.system.DefaultRV32Config.fir@191989.6 Arbiter.scala 128:19:freechips.rocketchip.system.DefaultRV32Config.fir@191998.6]
  assign dataArb_io_out_bits_eccMask = dataArb_io_in_0_valid ? dataArb_io_in_0_bits_eccMask : 4'hf; // @[Arbiter.scala 124:15:freechips.rocketchip.system.DefaultRV32Config.fir@191970.4 Arbiter.scala 128:19:freechips.rocketchip.system.DefaultRV32Config.fir@191978.6 Arbiter.scala 128:19:freechips.rocketchip.system.DefaultRV32Config.fir@191987.6 Arbiter.scala 128:19:freechips.rocketchip.system.DefaultRV32Config.fir@191996.6]
  assign dataArb_io_out_bits_way_en = dataArb_io_in_0_valid ? dataArb_io_in_0_bits_way_en : dataArb__GEN_8; // @[Arbiter.scala 124:15:freechips.rocketchip.system.DefaultRV32Config.fir@191969.4 Arbiter.scala 128:19:freechips.rocketchip.system.DefaultRV32Config.fir@191977.6 Arbiter.scala 128:19:freechips.rocketchip.system.DefaultRV32Config.fir@191986.6 Arbiter.scala 128:19:freechips.rocketchip.system.DefaultRV32Config.fir@191995.6]
  assign _T_7 = {MaxPeriodFibonacciLFSR_io_out_7,MaxPeriodFibonacciLFSR_io_out_6,MaxPeriodFibonacciLFSR_io_out_5,MaxPeriodFibonacciLFSR_io_out_4,MaxPeriodFibonacciLFSR_io_out_3,MaxPeriodFibonacciLFSR_io_out_2,MaxPeriodFibonacciLFSR_io_out_1,MaxPeriodFibonacciLFSR_io_out_0}; // @[PRNG.scala 86:17:freechips.rocketchip.system.DefaultRV32Config.fir@192146.4]
  assign _T_15 = {MaxPeriodFibonacciLFSR_io_out_15,MaxPeriodFibonacciLFSR_io_out_14,MaxPeriodFibonacciLFSR_io_out_13,MaxPeriodFibonacciLFSR_io_out_12,MaxPeriodFibonacciLFSR_io_out_11,MaxPeriodFibonacciLFSR_io_out_10,MaxPeriodFibonacciLFSR_io_out_9,MaxPeriodFibonacciLFSR_io_out_8,_T_7}; // @[PRNG.scala 86:17:freechips.rocketchip.system.DefaultRV32Config.fir@192154.4]
  assign _T_16 = io_cpu_req_ready & io_cpu_req_valid; // @[Decoupled.scala 40:37:freechips.rocketchip.system.DefaultRV32Config.fir@192188.4]
  assign _T_2338 = blockProbeAfterGrantCount > 3'h0; // @[DCache.scala 709:65:freechips.rocketchip.system.DefaultRV32Config.fir@195310.4]
  assign lrscValid = lrscCount > 7'h3; // @[DCache.scala 424:29:freechips.rocketchip.system.DefaultRV32Config.fir@193433.4]
  assign block_probe_for_core_progress = _T_2338 | lrscValid; // @[DCache.scala 709:69:freechips.rocketchip.system.DefaultRV32Config.fir@195311.4]
  assign _T_365 = s1_probe | s2_probe; // @[DCache.scala 286:34:freechips.rocketchip.system.DefaultRV32Config.fir@192768.4]
  assign _T_366 = release_state != 3'h0; // @[DCache.scala 286:63:freechips.rocketchip.system.DefaultRV32Config.fir@192769.4]
  assign releaseInFlight = _T_365 | _T_366; // @[DCache.scala 286:46:freechips.rocketchip.system.DefaultRV32Config.fir@192770.4]
  assign _T_2339 = auto_out_b_bits_address ^ release_ack_addr; // @[DCache.scala 710:88:freechips.rocketchip.system.DefaultRV32Config.fir@195312.4]
  assign _T_2341 = _T_2339[11:6] == 6'h0; // @[DCache.scala 710:124:freechips.rocketchip.system.DefaultRV32Config.fir@195314.4]
  assign block_probe_for_pending_release_ack = release_ack_wait & _T_2341; // @[DCache.scala 710:62:freechips.rocketchip.system.DefaultRV32Config.fir@195315.4]
  assign _T_2342 = releaseInFlight | block_probe_for_pending_release_ack; // @[DCache.scala 711:50:freechips.rocketchip.system.DefaultRV32Config.fir@195316.4]
  assign block_probe_for_ordering = _T_2342 | grantInProgress; // @[DCache.scala 711:89:freechips.rocketchip.system.DefaultRV32Config.fir@195317.4]
  assign _T_2346 = block_probe_for_core_progress | block_probe_for_ordering; // @[DCache.scala 713:79:freechips.rocketchip.system.DefaultRV32Config.fir@195322.4]
  assign _T_2347 = _T_2346 | s1_valid; // @[DCache.scala 713:107:freechips.rocketchip.system.DefaultRV32Config.fir@195323.4]
  assign _T_2348 = _T_2347 | s2_valid; // @[DCache.scala 713:119:freechips.rocketchip.system.DefaultRV32Config.fir@195324.4]
  assign _T_2349 = ~_T_2348; // @[DCache.scala 713:47:freechips.rocketchip.system.DefaultRV32Config.fir@195325.4]
  assign tl_out__b_ready = metaArb_io_in_6_ready & _T_2349; // @[DCache.scala 713:44:freechips.rocketchip.system.DefaultRV32Config.fir@195326.4]
  assign _T_17 = tl_out__b_ready & auto_out_b_valid; // @[Decoupled.scala 40:37:freechips.rocketchip.system.DefaultRV32Config.fir@192191.4]
  assign _T_19 = ~io_cpu_s1_kill; // @[DCache.scala 163:37:freechips.rocketchip.system.DefaultRV32Config.fir@192209.4]
  assign s1_valid_masked = s1_valid & _T_19; // @[DCache.scala 163:34:freechips.rocketchip.system.DefaultRV32Config.fir@192210.4]
  assign _T_640 = {probe_bits_param,s2_probe_state_state}; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@193206.4]
  assign _T_697 = 4'h3 == _T_640; // @[Misc.scala 55:20:freechips.rocketchip.system.DefaultRV32Config.fir@193263.4]
  assign _T_693 = 4'h2 == _T_640; // @[Misc.scala 55:20:freechips.rocketchip.system.DefaultRV32Config.fir@193259.4]
  assign _T_689 = 4'h1 == _T_640; // @[Misc.scala 55:20:freechips.rocketchip.system.DefaultRV32Config.fir@193255.4]
  assign _T_685 = 4'h0 == _T_640; // @[Misc.scala 55:20:freechips.rocketchip.system.DefaultRV32Config.fir@193251.4]
  assign _T_681 = 4'h7 == _T_640; // @[Misc.scala 55:20:freechips.rocketchip.system.DefaultRV32Config.fir@193247.4]
  assign _T_677 = 4'h6 == _T_640; // @[Misc.scala 55:20:freechips.rocketchip.system.DefaultRV32Config.fir@193243.4]
  assign _T_673 = 4'h5 == _T_640; // @[Misc.scala 55:20:freechips.rocketchip.system.DefaultRV32Config.fir@193239.4]
  assign _T_669 = 4'h4 == _T_640; // @[Misc.scala 55:20:freechips.rocketchip.system.DefaultRV32Config.fir@193235.4]
  assign _T_665 = 4'hb == _T_640; // @[Misc.scala 55:20:freechips.rocketchip.system.DefaultRV32Config.fir@193231.4]
  assign _T_661 = 4'ha == _T_640; // @[Misc.scala 55:20:freechips.rocketchip.system.DefaultRV32Config.fir@193227.4]
  assign _T_657 = 4'h9 == _T_640; // @[Misc.scala 55:20:freechips.rocketchip.system.DefaultRV32Config.fir@193223.4]
  assign _T_653 = 4'h8 == _T_640; // @[Misc.scala 55:20:freechips.rocketchip.system.DefaultRV32Config.fir@193219.4]
  assign _T_670 = _T_669 ? 1'h0 : _T_665; // @[Misc.scala 37:9:freechips.rocketchip.system.DefaultRV32Config.fir@193236.4]
  assign _T_674 = _T_673 ? 1'h0 : _T_670; // @[Misc.scala 37:9:freechips.rocketchip.system.DefaultRV32Config.fir@193240.4]
  assign _T_678 = _T_677 ? 1'h0 : _T_674; // @[Misc.scala 37:9:freechips.rocketchip.system.DefaultRV32Config.fir@193244.4]
  assign _T_682 = _T_681 | _T_678; // @[Misc.scala 37:9:freechips.rocketchip.system.DefaultRV32Config.fir@193248.4]
  assign _T_686 = _T_685 ? 1'h0 : _T_682; // @[Misc.scala 37:9:freechips.rocketchip.system.DefaultRV32Config.fir@193252.4]
  assign _T_690 = _T_689 ? 1'h0 : _T_686; // @[Misc.scala 37:9:freechips.rocketchip.system.DefaultRV32Config.fir@193256.4]
  assign _T_694 = _T_693 ? 1'h0 : _T_690; // @[Misc.scala 37:9:freechips.rocketchip.system.DefaultRV32Config.fir@193260.4]
  assign s2_prb_ack_data = _T_697 | _T_694; // @[Misc.scala 37:9:freechips.rocketchip.system.DefaultRV32Config.fir@193264.4]
  assign _T_2399 = s2_probe_state_state > 2'h0; // @[Metadata.scala 50:45:freechips.rocketchip.system.DefaultRV32Config.fir@195454.10]
  assign _T_2365 = _T_2362 == 10'h1; // @[Edges.scala 233:25:freechips.rocketchip.system.DefaultRV32Config.fir@195348.4]
  assign _T_2410 = release_state == 3'h1; // @[package.scala 15:47:freechips.rocketchip.system.DefaultRV32Config.fir@195507.4]
  assign _T_2411 = release_state == 3'h6; // @[package.scala 15:47:freechips.rocketchip.system.DefaultRV32Config.fir@195508.4]
  assign _T_2412 = _T_2410 | _T_2411; // @[package.scala 64:59:freechips.rocketchip.system.DefaultRV32Config.fir@195509.4]
  assign _T_2409 = release_state == 3'h2; // @[DCache.scala 779:25:freechips.rocketchip.system.DefaultRV32Config.fir@195500.4]
  assign _T_2408 = release_state == 3'h3; // @[DCache.scala 774:25:freechips.rocketchip.system.DefaultRV32Config.fir@195492.4]
  assign _GEN_310 = _T_2409 ? 3'h5 : 3'h4; // @[DCache.scala 779:48:freechips.rocketchip.system.DefaultRV32Config.fir@195501.4]
  assign tl_out__c_bits_opcode = _T_2412 ? 3'h7 : _GEN_310; // @[DCache.scala 783:81:freechips.rocketchip.system.DefaultRV32Config.fir@195510.4]
  assign tl_out__c_bits_size = _T_2412 ? 4'h6 : probe_bits_size; // @[DCache.scala 783:81:freechips.rocketchip.system.DefaultRV32Config.fir@195510.4]
  assign _T_2356 = 27'hfff << tl_out__c_bits_size; // @[package.scala 207:77:freechips.rocketchip.system.DefaultRV32Config.fir@195338.4]
  assign _T_2358 = ~_T_2356[11:0]; // @[package.scala 207:46:freechips.rocketchip.system.DefaultRV32Config.fir@195340.4]
  assign _T_2361 = tl_out__c_bits_opcode[0] ? _T_2358[11:2] : 10'h0; // @[Edges.scala 222:14:freechips.rocketchip.system.DefaultRV32Config.fir@195343.4]
  assign _T_2366 = _T_2361 == 10'h0; // @[Edges.scala 233:47:freechips.rocketchip.system.DefaultRV32Config.fir@195349.4]
  assign c_last = _T_2365 | _T_2366; // @[Edges.scala 233:37:freechips.rocketchip.system.DefaultRV32Config.fir@195350.4]
  assign _T_2407 = release_state == 3'h5; // @[DCache.scala 770:25:freechips.rocketchip.system.DefaultRV32Config.fir@195485.4]
  assign c_first = _T_2362 == 10'h0; // @[Edges.scala 232:25:freechips.rocketchip.system.DefaultRV32Config.fir@195347.4]
  assign _T_2381 = c_first & release_ack_wait; // @[DCache.scala 732:56:freechips.rocketchip.system.DefaultRV32Config.fir@195405.4]
  assign _T_2382 = ~_T_2381; // @[DCache.scala 732:46:freechips.rocketchip.system.DefaultRV32Config.fir@195406.4]
  assign _T_2383 = s2_release_data_valid & _T_2382; // @[DCache.scala 732:43:freechips.rocketchip.system.DefaultRV32Config.fir@195407.4]
  assign _GEN_259 = s2_prb_ack_data ? _T_2383 : 1'h1; // @[DCache.scala 748:36:freechips.rocketchip.system.DefaultRV32Config.fir@195450.8]
  assign _GEN_269 = pma_checker__T_2026 ? _T_2383 : _GEN_259; // @[DCache.scala 746:28:freechips.rocketchip.system.DefaultRV32Config.fir@195446.6]
  assign _GEN_280 = s2_probe ? _GEN_269 : _T_2383; // @[DCache.scala 744:21:freechips.rocketchip.system.DefaultRV32Config.fir@195442.4]
  assign _GEN_297 = _T_2407 | _GEN_280; // @[DCache.scala 770:47:freechips.rocketchip.system.DefaultRV32Config.fir@195486.4]
  assign tl_out__c_valid = _T_2408 | _GEN_297; // @[DCache.scala 774:48:freechips.rocketchip.system.DefaultRV32Config.fir@195493.4]
  assign _T_2354 = auto_out_c_ready & tl_out__c_valid; // @[Decoupled.scala 40:37:freechips.rocketchip.system.DefaultRV32Config.fir@195336.4]
  assign releaseDone = c_last & _T_2354; // @[Edges.scala 234:22:freechips.rocketchip.system.DefaultRV32Config.fir@195351.4]
  assign _T_2401 = ~releaseDone; // @[DCache.scala 756:22:freechips.rocketchip.system.DefaultRV32Config.fir@195463.12]
  assign _GEN_257 = _T_2399 | _T_2401; // @[DCache.scala 750:45:freechips.rocketchip.system.DefaultRV32Config.fir@195455.10]
  assign _GEN_267 = s2_prb_ack_data | _GEN_257; // @[DCache.scala 748:36:freechips.rocketchip.system.DefaultRV32Config.fir@195450.8]
  assign probeNack = pma_checker__T_2026 | _GEN_267; // @[DCache.scala 746:28:freechips.rocketchip.system.DefaultRV32Config.fir@195446.6]
  assign _T_30 = s1_req_cmd == 5'h0; // @[Consts.scala 82:31:freechips.rocketchip.system.DefaultRV32Config.fir@192264.4]
  assign _T_31 = s1_req_cmd == 5'h6; // @[Consts.scala 82:48:freechips.rocketchip.system.DefaultRV32Config.fir@192265.4]
  assign _T_32 = _T_30 | _T_31; // @[Consts.scala 82:41:freechips.rocketchip.system.DefaultRV32Config.fir@192266.4]
  assign _T_33 = s1_req_cmd == 5'h7; // @[Consts.scala 82:65:freechips.rocketchip.system.DefaultRV32Config.fir@192267.4]
  assign _T_34 = _T_32 | _T_33; // @[Consts.scala 82:58:freechips.rocketchip.system.DefaultRV32Config.fir@192268.4]
  assign _T_35 = s1_req_cmd == 5'h4; // @[package.scala 15:47:freechips.rocketchip.system.DefaultRV32Config.fir@192269.4]
  assign _T_36 = s1_req_cmd == 5'h9; // @[package.scala 15:47:freechips.rocketchip.system.DefaultRV32Config.fir@192270.4]
  assign _T_39 = _T_35 | _T_36; // @[package.scala 64:59:freechips.rocketchip.system.DefaultRV32Config.fir@192273.4]
  assign _T_37 = s1_req_cmd == 5'ha; // @[package.scala 15:47:freechips.rocketchip.system.DefaultRV32Config.fir@192271.4]
  assign _T_40 = _T_39 | _T_37; // @[package.scala 64:59:freechips.rocketchip.system.DefaultRV32Config.fir@192274.4]
  assign _T_38 = s1_req_cmd == 5'hb; // @[package.scala 15:47:freechips.rocketchip.system.DefaultRV32Config.fir@192272.4]
  assign _T_41 = _T_40 | _T_38; // @[package.scala 64:59:freechips.rocketchip.system.DefaultRV32Config.fir@192275.4]
  assign _T_42 = s1_req_cmd == 5'h8; // @[package.scala 15:47:freechips.rocketchip.system.DefaultRV32Config.fir@192276.4]
  assign _T_43 = s1_req_cmd == 5'hc; // @[package.scala 15:47:freechips.rocketchip.system.DefaultRV32Config.fir@192277.4]
  assign _T_47 = _T_42 | _T_43; // @[package.scala 64:59:freechips.rocketchip.system.DefaultRV32Config.fir@192281.4]
  assign _T_44 = s1_req_cmd == 5'hd; // @[package.scala 15:47:freechips.rocketchip.system.DefaultRV32Config.fir@192278.4]
  assign _T_48 = _T_47 | _T_44; // @[package.scala 64:59:freechips.rocketchip.system.DefaultRV32Config.fir@192282.4]
  assign _T_45 = s1_req_cmd == 5'he; // @[package.scala 15:47:freechips.rocketchip.system.DefaultRV32Config.fir@192279.4]
  assign _T_49 = _T_48 | _T_45; // @[package.scala 64:59:freechips.rocketchip.system.DefaultRV32Config.fir@192283.4]
  assign _T_46 = s1_req_cmd == 5'hf; // @[package.scala 15:47:freechips.rocketchip.system.DefaultRV32Config.fir@192280.4]
  assign _T_50 = _T_49 | _T_46; // @[package.scala 64:59:freechips.rocketchip.system.DefaultRV32Config.fir@192284.4]
  assign _T_51 = _T_41 | _T_50; // @[Consts.scala 80:44:freechips.rocketchip.system.DefaultRV32Config.fir@192285.4]
  assign s1_read = _T_34 | _T_51; // @[Consts.scala 82:75:freechips.rocketchip.system.DefaultRV32Config.fir@192286.4]
  assign _T_402 = s2_req_cmd == 5'h1; // @[Consts.scala 83:32:freechips.rocketchip.system.DefaultRV32Config.fir@192828.4]
  assign _T_403 = s2_req_cmd == 5'h11; // @[Consts.scala 83:49:freechips.rocketchip.system.DefaultRV32Config.fir@192829.4]
  assign _T_404 = _T_402 | _T_403; // @[Consts.scala 83:42:freechips.rocketchip.system.DefaultRV32Config.fir@192830.4]
  assign _T_405 = s2_req_cmd == 5'h7; // @[Consts.scala 83:66:freechips.rocketchip.system.DefaultRV32Config.fir@192831.4]
  assign _T_406 = _T_404 | _T_405; // @[Consts.scala 83:59:freechips.rocketchip.system.DefaultRV32Config.fir@192832.4]
  assign _T_407 = s2_req_cmd == 5'h4; // @[package.scala 15:47:freechips.rocketchip.system.DefaultRV32Config.fir@192833.4]
  assign _T_408 = s2_req_cmd == 5'h9; // @[package.scala 15:47:freechips.rocketchip.system.DefaultRV32Config.fir@192834.4]
  assign _T_411 = _T_407 | _T_408; // @[package.scala 64:59:freechips.rocketchip.system.DefaultRV32Config.fir@192837.4]
  assign _T_409 = s2_req_cmd == 5'ha; // @[package.scala 15:47:freechips.rocketchip.system.DefaultRV32Config.fir@192835.4]
  assign _T_412 = _T_411 | _T_409; // @[package.scala 64:59:freechips.rocketchip.system.DefaultRV32Config.fir@192838.4]
  assign _T_410 = s2_req_cmd == 5'hb; // @[package.scala 15:47:freechips.rocketchip.system.DefaultRV32Config.fir@192836.4]
  assign _T_413 = _T_412 | _T_410; // @[package.scala 64:59:freechips.rocketchip.system.DefaultRV32Config.fir@192839.4]
  assign _T_414 = s2_req_cmd == 5'h8; // @[package.scala 15:47:freechips.rocketchip.system.DefaultRV32Config.fir@192840.4]
  assign _T_415 = s2_req_cmd == 5'hc; // @[package.scala 15:47:freechips.rocketchip.system.DefaultRV32Config.fir@192841.4]
  assign _T_419 = _T_414 | _T_415; // @[package.scala 64:59:freechips.rocketchip.system.DefaultRV32Config.fir@192845.4]
  assign _T_416 = s2_req_cmd == 5'hd; // @[package.scala 15:47:freechips.rocketchip.system.DefaultRV32Config.fir@192842.4]
  assign _T_420 = _T_419 | _T_416; // @[package.scala 64:59:freechips.rocketchip.system.DefaultRV32Config.fir@192846.4]
  assign _T_417 = s2_req_cmd == 5'he; // @[package.scala 15:47:freechips.rocketchip.system.DefaultRV32Config.fir@192843.4]
  assign _T_421 = _T_420 | _T_417; // @[package.scala 64:59:freechips.rocketchip.system.DefaultRV32Config.fir@192847.4]
  assign _T_418 = s2_req_cmd == 5'hf; // @[package.scala 15:47:freechips.rocketchip.system.DefaultRV32Config.fir@192844.4]
  assign _T_422 = _T_421 | _T_418; // @[package.scala 64:59:freechips.rocketchip.system.DefaultRV32Config.fir@192848.4]
  assign _T_423 = _T_413 | _T_422; // @[Consts.scala 80:44:freechips.rocketchip.system.DefaultRV32Config.fir@192849.4]
  assign s2_write = _T_406 | _T_423; // @[Consts.scala 83:76:freechips.rocketchip.system.DefaultRV32Config.fir@192850.4]
  assign _T_977 = s2_valid & s2_write; // @[DCache.scala 456:39:freechips.rocketchip.system.DefaultRV32Config.fir@193647.4]
  assign pstore1_valid_likely = _T_977 | pstore1_held; // @[DCache.scala 456:51:freechips.rocketchip.system.DefaultRV32Config.fir@193648.4]
  assign _T_1094 = pstore1_addr[11:2] == s1_req_addr[11:2]; // @[DCache.scala 508:31:freechips.rocketchip.system.DefaultRV32Config.fir@193812.4]
  assign _T_52 = s1_req_cmd == 5'h1; // @[Consts.scala 83:32:freechips.rocketchip.system.DefaultRV32Config.fir@192287.4]
  assign _T_53 = s1_req_cmd == 5'h11; // @[Consts.scala 83:49:freechips.rocketchip.system.DefaultRV32Config.fir@192288.4]
  assign _T_54 = _T_52 | _T_53; // @[Consts.scala 83:42:freechips.rocketchip.system.DefaultRV32Config.fir@192289.4]
  assign _T_56 = _T_54 | _T_33; // @[Consts.scala 83:59:freechips.rocketchip.system.DefaultRV32Config.fir@192291.4]
  assign s1_write = _T_56 | _T_51; // @[Consts.scala 83:76:freechips.rocketchip.system.DefaultRV32Config.fir@192309.4]
  assign _T_1102 = |pstore1_mask[3]; // @[DCache.scala 1076:66:freechips.rocketchip.system.DefaultRV32Config.fir@193820.4]
  assign _T_1101 = |pstore1_mask[2]; // @[DCache.scala 1076:66:freechips.rocketchip.system.DefaultRV32Config.fir@193819.4]
  assign _T_1100 = |pstore1_mask[1]; // @[DCache.scala 1076:66:freechips.rocketchip.system.DefaultRV32Config.fir@193818.4]
  assign _T_1099 = |pstore1_mask[0]; // @[DCache.scala 1076:66:freechips.rocketchip.system.DefaultRV32Config.fir@193817.4]
  assign _T_1105 = {_T_1102,_T_1101,_T_1100,_T_1099}; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@193823.4]
  assign _T_1112 = {_T_1105[3],_T_1105[2],_T_1105[1],_T_1105[0]}; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@193830.4]
  assign _T_332 = s1_req_size >= 2'h1; // @[AMOALU.scala 17:57:freechips.rocketchip.system.DefaultRV32Config.fir@192724.4]
  assign _T_334 = s1_req_addr[0] | _T_332; // @[AMOALU.scala 17:46:freechips.rocketchip.system.DefaultRV32Config.fir@192726.4]
  assign _T_336 = s1_req_addr[0] ? 1'h0 : 1'h1; // @[AMOALU.scala 18:22:freechips.rocketchip.system.DefaultRV32Config.fir@192728.4]
  assign _T_337 = {_T_334,_T_336}; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@192729.4]
  assign _T_339 = s1_req_addr[1] ? _T_337 : 2'h0; // @[AMOALU.scala 17:22:freechips.rocketchip.system.DefaultRV32Config.fir@192731.4]
  assign _T_340 = s1_req_size >= 2'h2; // @[AMOALU.scala 17:57:freechips.rocketchip.system.DefaultRV32Config.fir@192732.4]
  assign _T_341 = _T_340 ? 2'h3 : 2'h0; // @[AMOALU.scala 17:51:freechips.rocketchip.system.DefaultRV32Config.fir@192733.4]
  assign _T_342 = _T_339 | _T_341; // @[AMOALU.scala 17:46:freechips.rocketchip.system.DefaultRV32Config.fir@192734.4]
  assign _T_344 = s1_req_addr[1] ? 2'h0 : _T_337; // @[AMOALU.scala 18:22:freechips.rocketchip.system.DefaultRV32Config.fir@192736.4]
  assign s1_mask_xwr = {_T_342,_T_344}; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@192737.4]
  assign _T_1120 = |s1_mask_xwr[3]; // @[DCache.scala 1076:66:freechips.rocketchip.system.DefaultRV32Config.fir@193838.4]
  assign _T_1119 = |s1_mask_xwr[2]; // @[DCache.scala 1076:66:freechips.rocketchip.system.DefaultRV32Config.fir@193837.4]
  assign _T_1118 = |s1_mask_xwr[1]; // @[DCache.scala 1076:66:freechips.rocketchip.system.DefaultRV32Config.fir@193836.4]
  assign _T_1117 = |s1_mask_xwr[0]; // @[DCache.scala 1076:66:freechips.rocketchip.system.DefaultRV32Config.fir@193835.4]
  assign _T_1123 = {_T_1120,_T_1119,_T_1118,_T_1117}; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@193841.4]
  assign _T_1130 = {_T_1123[3],_T_1123[2],_T_1123[1],_T_1123[0]}; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@193848.4]
  assign _T_1131 = _T_1112 & _T_1130; // @[DCache.scala 509:38:freechips.rocketchip.system.DefaultRV32Config.fir@193849.4]
  assign _T_1132 = |_T_1131; // @[DCache.scala 509:66:freechips.rocketchip.system.DefaultRV32Config.fir@193850.4]
  assign _T_1133 = pstore1_mask & s1_mask_xwr; // @[DCache.scala 509:77:freechips.rocketchip.system.DefaultRV32Config.fir@193851.4]
  assign _T_1134 = |_T_1133; // @[DCache.scala 509:92:freechips.rocketchip.system.DefaultRV32Config.fir@193852.4]
  assign _T_1135 = s1_write ? _T_1132 : _T_1134; // @[DCache.scala 509:8:freechips.rocketchip.system.DefaultRV32Config.fir@193853.4]
  assign _T_1136 = _T_1094 & _T_1135; // @[DCache.scala 508:68:freechips.rocketchip.system.DefaultRV32Config.fir@193854.4]
  assign _T_1137 = pstore1_valid_likely & _T_1136; // @[DCache.scala 511:27:freechips.rocketchip.system.DefaultRV32Config.fir@193855.4]
  assign _T_1140 = pstore2_addr[11:2] == s1_req_addr[11:2]; // @[DCache.scala 508:31:freechips.rocketchip.system.DefaultRV32Config.fir@193858.4]
  assign _T_1148 = |mask[3]; // @[DCache.scala 1076:66:freechips.rocketchip.system.DefaultRV32Config.fir@193866.4]
  assign _T_1147 = |mask[2]; // @[DCache.scala 1076:66:freechips.rocketchip.system.DefaultRV32Config.fir@193865.4]
  assign _T_1146 = |mask[1]; // @[DCache.scala 1076:66:freechips.rocketchip.system.DefaultRV32Config.fir@193864.4]
  assign _T_1145 = |mask[0]; // @[DCache.scala 1076:66:freechips.rocketchip.system.DefaultRV32Config.fir@193863.4]
  assign _T_1151 = {_T_1148,_T_1147,_T_1146,_T_1145}; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@193869.4]
  assign _T_1158 = {_T_1151[3],_T_1151[2],_T_1151[1],_T_1151[0]}; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@193876.4]
  assign _T_1177 = _T_1158 & _T_1130; // @[DCache.scala 509:38:freechips.rocketchip.system.DefaultRV32Config.fir@193895.4]
  assign _T_1178 = |_T_1177; // @[DCache.scala 509:66:freechips.rocketchip.system.DefaultRV32Config.fir@193896.4]
  assign _T_1179 = mask & s1_mask_xwr; // @[DCache.scala 509:77:freechips.rocketchip.system.DefaultRV32Config.fir@193897.4]
  assign _T_1180 = |_T_1179; // @[DCache.scala 509:92:freechips.rocketchip.system.DefaultRV32Config.fir@193898.4]
  assign _T_1181 = s1_write ? _T_1178 : _T_1180; // @[DCache.scala 509:8:freechips.rocketchip.system.DefaultRV32Config.fir@193899.4]
  assign _T_1182 = _T_1140 & _T_1181; // @[DCache.scala 508:68:freechips.rocketchip.system.DefaultRV32Config.fir@193900.4]
  assign _T_1183 = pstore2_valid & _T_1182; // @[DCache.scala 512:21:freechips.rocketchip.system.DefaultRV32Config.fir@193901.4]
  assign s1_hazard = _T_1137 | _T_1183; // @[DCache.scala 511:69:freechips.rocketchip.system.DefaultRV32Config.fir@193902.4]
  assign s1_raw_hazard = s1_read & s1_hazard; // @[DCache.scala 513:31:freechips.rocketchip.system.DefaultRV32Config.fir@193903.4]
  assign _T_1184 = s1_valid & s1_raw_hazard; // @[DCache.scala 518:18:freechips.rocketchip.system.DefaultRV32Config.fir@193905.4]
  assign _T_362 = {io_cpu_s2_xcpt_ma_ld,io_cpu_s2_xcpt_ma_st,io_cpu_s2_xcpt_pf_ld,io_cpu_s2_xcpt_pf_st,io_cpu_s2_xcpt_ae_ld,io_cpu_s2_xcpt_ae_st}; // @[DCache.scala 284:54:freechips.rocketchip.system.DefaultRV32Config.fir@192762.4]
  assign _T_363 = |_T_362; // @[DCache.scala 284:61:freechips.rocketchip.system.DefaultRV32Config.fir@192763.4]
  assign _T_364 = ~_T_363; // @[DCache.scala 284:38:freechips.rocketchip.system.DefaultRV32Config.fir@192764.4]
  assign s2_valid_no_xcpt = s2_valid & _T_364; // @[DCache.scala 284:35:freechips.rocketchip.system.DefaultRV32Config.fir@192765.4]
  assign s2_valid_masked = s2_valid_no_xcpt & s2_not_nacked_in_s1; // @[DCache.scala 289:42:freechips.rocketchip.system.DefaultRV32Config.fir@192775.4]
  assign _T_603 = ~pma_checker__T_2026; // @[DCache.scala 349:74:freechips.rocketchip.system.DefaultRV32Config.fir@193144.4]
  assign _T_604 = s2_valid_masked & _T_603; // @[DCache.scala 349:71:freechips.rocketchip.system.DefaultRV32Config.fir@193145.4]
  assign _T_523 = s2_req_cmd == 5'h3; // @[Consts.scala 84:54:freechips.rocketchip.system.DefaultRV32Config.fir@193055.4]
  assign _T_524 = s2_write | _T_523; // @[Consts.scala 84:47:freechips.rocketchip.system.DefaultRV32Config.fir@193056.4]
  assign _T_525 = s2_req_cmd == 5'h6; // @[Consts.scala 84:71:freechips.rocketchip.system.DefaultRV32Config.fir@193057.4]
  assign _T_526 = _T_524 | _T_525; // @[Consts.scala 84:64:freechips.rocketchip.system.DefaultRV32Config.fir@193058.4]
  assign _T_528 = {s2_write,_T_526,s2_hit_state_state}; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@193060.4]
  assign _T_586 = 4'h3 == _T_528; // @[Misc.scala 48:20:freechips.rocketchip.system.DefaultRV32Config.fir@193118.4]
  assign _T_583 = 4'h2 == _T_528; // @[Misc.scala 48:20:freechips.rocketchip.system.DefaultRV32Config.fir@193115.4]
  assign _T_580 = 4'h1 == _T_528; // @[Misc.scala 48:20:freechips.rocketchip.system.DefaultRV32Config.fir@193112.4]
  assign _T_577 = 4'h7 == _T_528; // @[Misc.scala 48:20:freechips.rocketchip.system.DefaultRV32Config.fir@193109.4]
  assign _T_574 = 4'h6 == _T_528; // @[Misc.scala 48:20:freechips.rocketchip.system.DefaultRV32Config.fir@193106.4]
  assign _T_571 = 4'hf == _T_528; // @[Misc.scala 48:20:freechips.rocketchip.system.DefaultRV32Config.fir@193103.4]
  assign _T_568 = 4'he == _T_528; // @[Misc.scala 48:20:freechips.rocketchip.system.DefaultRV32Config.fir@193100.4]
  assign _T_565 = 4'h0 == _T_528; // @[Misc.scala 48:20:freechips.rocketchip.system.DefaultRV32Config.fir@193097.4]
  assign _T_562 = 4'h5 == _T_528; // @[Misc.scala 48:20:freechips.rocketchip.system.DefaultRV32Config.fir@193094.4]
  assign _T_559 = 4'h4 == _T_528; // @[Misc.scala 48:20:freechips.rocketchip.system.DefaultRV32Config.fir@193091.4]
  assign _T_556 = 4'hd == _T_528; // @[Misc.scala 48:20:freechips.rocketchip.system.DefaultRV32Config.fir@193088.4]
  assign _T_553 = 4'hc == _T_528; // @[Misc.scala 48:20:freechips.rocketchip.system.DefaultRV32Config.fir@193085.4]
  assign _T_572 = _T_571 | _T_568; // @[Misc.scala 34:9:freechips.rocketchip.system.DefaultRV32Config.fir@193104.4]
  assign _T_575 = _T_574 | _T_572; // @[Misc.scala 34:9:freechips.rocketchip.system.DefaultRV32Config.fir@193107.4]
  assign _T_578 = _T_577 | _T_575; // @[Misc.scala 34:9:freechips.rocketchip.system.DefaultRV32Config.fir@193110.4]
  assign _T_581 = _T_580 | _T_578; // @[Misc.scala 34:9:freechips.rocketchip.system.DefaultRV32Config.fir@193113.4]
  assign _T_584 = _T_583 | _T_581; // @[Misc.scala 34:9:freechips.rocketchip.system.DefaultRV32Config.fir@193116.4]
  assign s2_hit = _T_586 | _T_584; // @[Misc.scala 34:9:freechips.rocketchip.system.DefaultRV32Config.fir@193119.4]
  assign s2_valid_hit_maybe_flush_pre_data_ecc_and_waw = _T_604 & s2_hit; // @[DCache.scala 349:89:freechips.rocketchip.system.DefaultRV32Config.fir@193146.4]
  assign _T_380 = s2_req_cmd == 5'h0; // @[Consts.scala 82:31:freechips.rocketchip.system.DefaultRV32Config.fir@192805.4]
  assign _T_382 = _T_380 | _T_525; // @[Consts.scala 82:41:freechips.rocketchip.system.DefaultRV32Config.fir@192807.4]
  assign _T_384 = _T_382 | _T_405; // @[Consts.scala 82:58:freechips.rocketchip.system.DefaultRV32Config.fir@192809.4]
  assign s2_read = _T_384 | _T_423; // @[Consts.scala 82:75:freechips.rocketchip.system.DefaultRV32Config.fir@192827.4]
  assign s2_readwrite = s2_read | s2_write; // @[DCache.scala 306:30:freechips.rocketchip.system.DefaultRV32Config.fir@192851.4]
  assign s2_valid_hit_pre_data_ecc_and_waw = s2_valid_hit_maybe_flush_pre_data_ecc_and_waw & s2_readwrite; // @[DCache.scala 370:89:freechips.rocketchip.system.DefaultRV32Config.fir@193147.4]
  assign _T_555 = _T_553 ? 2'h1 : 2'h0; // @[Misc.scala 34:36:freechips.rocketchip.system.DefaultRV32Config.fir@193087.4]
  assign _T_558 = _T_556 ? 2'h2 : _T_555; // @[Misc.scala 34:36:freechips.rocketchip.system.DefaultRV32Config.fir@193090.4]
  assign _T_561 = _T_559 ? 2'h1 : _T_558; // @[Misc.scala 34:36:freechips.rocketchip.system.DefaultRV32Config.fir@193093.4]
  assign _T_564 = _T_562 ? 2'h2 : _T_561; // @[Misc.scala 34:36:freechips.rocketchip.system.DefaultRV32Config.fir@193096.4]
  assign _T_567 = _T_565 ? 2'h0 : _T_564; // @[Misc.scala 34:36:freechips.rocketchip.system.DefaultRV32Config.fir@193099.4]
  assign _T_570 = _T_568 ? 2'h3 : _T_567; // @[Misc.scala 34:36:freechips.rocketchip.system.DefaultRV32Config.fir@193102.4]
  assign _T_573 = _T_571 ? 2'h3 : _T_570; // @[Misc.scala 34:36:freechips.rocketchip.system.DefaultRV32Config.fir@193105.4]
  assign _T_576 = _T_574 ? 2'h2 : _T_573; // @[Misc.scala 34:36:freechips.rocketchip.system.DefaultRV32Config.fir@193108.4]
  assign _T_579 = _T_577 ? 2'h3 : _T_576; // @[Misc.scala 34:36:freechips.rocketchip.system.DefaultRV32Config.fir@193111.4]
  assign _T_582 = _T_580 ? 2'h1 : _T_579; // @[Misc.scala 34:36:freechips.rocketchip.system.DefaultRV32Config.fir@193114.4]
  assign _T_585 = _T_583 ? 2'h2 : _T_582; // @[Misc.scala 34:36:freechips.rocketchip.system.DefaultRV32Config.fir@193117.4]
  assign s2_grow_param = _T_586 ? 2'h3 : _T_585; // @[Misc.scala 34:36:freechips.rocketchip.system.DefaultRV32Config.fir@193120.4]
  assign _T_764 = s2_hit_state_state == s2_grow_param; // @[Metadata.scala 46:46:freechips.rocketchip.system.DefaultRV32Config.fir@193340.4]
  assign s2_update_meta = ~_T_764; // @[Metadata.scala 47:40:freechips.rocketchip.system.DefaultRV32Config.fir@193341.4]
  assign _T_783 = s2_valid_hit_pre_data_ecc_and_waw & s2_update_meta; // @[DCache.scala 397:62:freechips.rocketchip.system.DefaultRV32Config.fir@193363.4]
  assign _T_784 = io_cpu_s2_nack | _T_783; // @[DCache.scala 397:24:freechips.rocketchip.system.DefaultRV32Config.fir@193364.4]
  assign s1_readwrite = s1_read | s1_write; // @[DCache.scala 185:30:freechips.rocketchip.system.DefaultRV32Config.fir@192310.4]
  assign _T_74 = s1_req_cmd == 5'h5; // @[DCache.scala 187:34:freechips.rocketchip.system.DefaultRV32Config.fir@192312.4]
  assign s1_flush_line = _T_74 & s1_req_size[0]; // @[DCache.scala 187:50:freechips.rocketchip.system.DefaultRV32Config.fir@192314.4]
  assign _T_227 = s1_readwrite | s1_flush_line; // @[DCache.scala 229:38:freechips.rocketchip.system.DefaultRV32Config.fir@192517.4]
  assign _T_228 = s1_req_cmd == 5'h17; // @[DCache.scala 229:69:freechips.rocketchip.system.DefaultRV32Config.fir@192518.4]
  assign s1_cmd_uses_tlb = _T_227 | _T_228; // @[DCache.scala 229:55:freechips.rocketchip.system.DefaultRV32Config.fir@192519.4]
  assign _T_242 = s1_valid & s1_cmd_uses_tlb; // @[DCache.scala 235:39:freechips.rocketchip.system.DefaultRV32Config.fir@192540.4]
  assign _T_243 = _T_242 & tlb_io_resp_miss; // @[DCache.scala 235:58:freechips.rocketchip.system.DefaultRV32Config.fir@192541.4]
  assign _GEN_118 = _T_784 | _T_243; // @[DCache.scala 397:82:freechips.rocketchip.system.DefaultRV32Config.fir@193365.4]
  assign _GEN_138 = _T_1184 | _GEN_118; // @[DCache.scala 518:36:freechips.rocketchip.system.DefaultRV32Config.fir@193906.4]
  assign _GEN_278 = probeNack | _GEN_138; // @[DCache.scala 759:24:freechips.rocketchip.system.DefaultRV32Config.fir@195468.6]
  assign s1_nack = s2_probe ? _GEN_278 : _GEN_138; // @[DCache.scala 744:21:freechips.rocketchip.system.DefaultRV32Config.fir@195442.4]
  assign _T_20 = ~s1_nack; // @[DCache.scala 164:41:freechips.rocketchip.system.DefaultRV32Config.fir@192211.4]
  assign s1_valid_not_nacked = s1_valid & _T_20; // @[DCache.scala 164:38:freechips.rocketchip.system.DefaultRV32Config.fir@192212.4]
  assign _T_22 = ~metaArb_io_out_bits_write; // @[DCache.scala 167:43:freechips.rocketchip.system.DefaultRV32Config.fir@192218.4]
  assign s0_clk_en = metaArb_io_out_valid & _T_22; // @[DCache.scala 167:40:freechips.rocketchip.system.DefaultRV32Config.fir@192219.4]
  assign s0_req_addr = {metaArb_io_out_bits_addr[31:6],io_cpu_req_bits_addr[5:0]}; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@192225.4]
  assign _T_26 = ~metaArb_io_in_7_ready; // @[DCache.scala 171:9:freechips.rocketchip.system.DefaultRV32Config.fir@192227.4]
  assign s0_req_phys = _T_26 | io_cpu_req_bits_phys; // @[DCache.scala 171:34:freechips.rocketchip.system.DefaultRV32Config.fir@192228.4]
  assign s1_sfence = s1_req_cmd == 5'h14; // @[DCache.scala 186:30:freechips.rocketchip.system.DefaultRV32Config.fir@192311.4]
  assign inWriteback = _T_2410 | _T_2409; // @[package.scala 64:59:freechips.rocketchip.system.DefaultRV32Config.fir@192329.4]
  assign _T_78 = release_state == 3'h0; // @[DCache.scala 203:38:freechips.rocketchip.system.DefaultRV32Config.fir@192332.4]
  assign _T_79 = ~cached_grant_wait; // @[DCache.scala 203:54:freechips.rocketchip.system.DefaultRV32Config.fir@192333.4]
  assign _T_80 = _T_78 & _T_79; // @[DCache.scala 203:51:freechips.rocketchip.system.DefaultRV32Config.fir@192334.4]
  assign _T_82 = _T_80 & _T_20; // @[DCache.scala 203:73:freechips.rocketchip.system.DefaultRV32Config.fir@192336.4]
  assign _T_84 = io_cpu_req_bits_cmd == 5'h0; // @[Consts.scala 82:31:freechips.rocketchip.system.DefaultRV32Config.fir@192346.4]
  assign _T_85 = io_cpu_req_bits_cmd == 5'h6; // @[Consts.scala 82:48:freechips.rocketchip.system.DefaultRV32Config.fir@192347.4]
  assign _T_86 = _T_84 | _T_85; // @[Consts.scala 82:41:freechips.rocketchip.system.DefaultRV32Config.fir@192348.4]
  assign _T_87 = io_cpu_req_bits_cmd == 5'h7; // @[Consts.scala 82:65:freechips.rocketchip.system.DefaultRV32Config.fir@192349.4]
  assign _T_88 = _T_86 | _T_87; // @[Consts.scala 82:58:freechips.rocketchip.system.DefaultRV32Config.fir@192350.4]
  assign _T_89 = io_cpu_req_bits_cmd == 5'h4; // @[package.scala 15:47:freechips.rocketchip.system.DefaultRV32Config.fir@192351.4]
  assign _T_90 = io_cpu_req_bits_cmd == 5'h9; // @[package.scala 15:47:freechips.rocketchip.system.DefaultRV32Config.fir@192352.4]
  assign _T_91 = io_cpu_req_bits_cmd == 5'ha; // @[package.scala 15:47:freechips.rocketchip.system.DefaultRV32Config.fir@192353.4]
  assign _T_92 = io_cpu_req_bits_cmd == 5'hb; // @[package.scala 15:47:freechips.rocketchip.system.DefaultRV32Config.fir@192354.4]
  assign _T_93 = _T_89 | _T_90; // @[package.scala 64:59:freechips.rocketchip.system.DefaultRV32Config.fir@192355.4]
  assign _T_94 = _T_93 | _T_91; // @[package.scala 64:59:freechips.rocketchip.system.DefaultRV32Config.fir@192356.4]
  assign _T_95 = _T_94 | _T_92; // @[package.scala 64:59:freechips.rocketchip.system.DefaultRV32Config.fir@192357.4]
  assign _T_96 = io_cpu_req_bits_cmd == 5'h8; // @[package.scala 15:47:freechips.rocketchip.system.DefaultRV32Config.fir@192358.4]
  assign _T_97 = io_cpu_req_bits_cmd == 5'hc; // @[package.scala 15:47:freechips.rocketchip.system.DefaultRV32Config.fir@192359.4]
  assign _T_98 = io_cpu_req_bits_cmd == 5'hd; // @[package.scala 15:47:freechips.rocketchip.system.DefaultRV32Config.fir@192360.4]
  assign _T_99 = io_cpu_req_bits_cmd == 5'he; // @[package.scala 15:47:freechips.rocketchip.system.DefaultRV32Config.fir@192361.4]
  assign _T_100 = io_cpu_req_bits_cmd == 5'hf; // @[package.scala 15:47:freechips.rocketchip.system.DefaultRV32Config.fir@192362.4]
  assign _T_101 = _T_96 | _T_97; // @[package.scala 64:59:freechips.rocketchip.system.DefaultRV32Config.fir@192363.4]
  assign _T_102 = _T_101 | _T_98; // @[package.scala 64:59:freechips.rocketchip.system.DefaultRV32Config.fir@192364.4]
  assign _T_103 = _T_102 | _T_99; // @[package.scala 64:59:freechips.rocketchip.system.DefaultRV32Config.fir@192365.4]
  assign _T_104 = _T_103 | _T_100; // @[package.scala 64:59:freechips.rocketchip.system.DefaultRV32Config.fir@192366.4]
  assign _T_105 = _T_95 | _T_104; // @[Consts.scala 80:44:freechips.rocketchip.system.DefaultRV32Config.fir@192367.4]
  assign s0_read = _T_88 | _T_105; // @[Consts.scala 82:75:freechips.rocketchip.system.DefaultRV32Config.fir@192368.4]
  assign _T_106 = io_cpu_req_bits_cmd == 5'h1; // @[package.scala 15:47:freechips.rocketchip.system.DefaultRV32Config.fir@192369.4]
  assign _T_107 = io_cpu_req_bits_cmd == 5'h3; // @[package.scala 15:47:freechips.rocketchip.system.DefaultRV32Config.fir@192370.4]
  assign _T_108 = _T_106 | _T_107; // @[package.scala 64:59:freechips.rocketchip.system.DefaultRV32Config.fir@192371.4]
  assign res = ~_T_108; // @[DCache.scala 1080:15:freechips.rocketchip.system.DefaultRV32Config.fir@192372.4]
  assign _T_135 = io_cpu_req_bits_cmd == 5'h11; // @[Consts.scala 83:49:freechips.rocketchip.system.DefaultRV32Config.fir@192399.4]
  assign _T_136 = _T_106 | _T_135; // @[Consts.scala 83:42:freechips.rocketchip.system.DefaultRV32Config.fir@192400.4]
  assign _T_138 = _T_136 | _T_87; // @[Consts.scala 83:59:freechips.rocketchip.system.DefaultRV32Config.fir@192402.4]
  assign _T_156 = _T_138 | _T_105; // @[Consts.scala 83:76:freechips.rocketchip.system.DefaultRV32Config.fir@192420.4]
  assign _T_160 = _T_156 & _T_135; // @[DCache.scala 1086:23:freechips.rocketchip.system.DefaultRV32Config.fir@192424.4]
  assign _T_161 = s0_read | _T_160; // @[DCache.scala 1085:21:freechips.rocketchip.system.DefaultRV32Config.fir@192425.4]
  assign _T_162 = ~_T_161; // @[DCache.scala 1081:12:freechips.rocketchip.system.DefaultRV32Config.fir@192426.4]
  assign _T_163 = _T_162 | res; // @[DCache.scala 1081:28:freechips.rocketchip.system.DefaultRV32Config.fir@192427.4]
  assign _T_165 = _T_163 | reset; // @[DCache.scala 1081:11:freechips.rocketchip.system.DefaultRV32Config.fir@192429.4]
  assign _T_166 = ~_T_165; // @[DCache.scala 1081:11:freechips.rocketchip.system.DefaultRV32Config.fir@192430.4]
  assign _T_167 = io_cpu_req_valid & res; // @[DCache.scala 212:46:freechips.rocketchip.system.DefaultRV32Config.fir@192435.4]
  assign _T_170 = ~dataArb_io_in_3_ready; // @[DCache.scala 218:9:freechips.rocketchip.system.DefaultRV32Config.fir@192444.4]
  assign _T_171 = _T_170 & s0_read; // @[DCache.scala 218:33:freechips.rocketchip.system.DefaultRV32Config.fir@192445.4]
  assign _GEN_28 = _T_171 ? 1'h0 : _T_82; // @[DCache.scala 218:45:freechips.rocketchip.system.DefaultRV32Config.fir@192446.4]
  assign _T_223 = io_cpu_req_valid & _T_161; // @[DCache.scala 219:75:freechips.rocketchip.system.DefaultRV32Config.fir@192500.4]
  assign _T_224 = dataArb_io_in_3_ready & _T_223; // @[DCache.scala 219:54:freechips.rocketchip.system.DefaultRV32Config.fir@192501.4]
  assign _GEN_30 = _T_26 ? 1'h0 : _GEN_28; // @[DCache.scala 226:34:freechips.rocketchip.system.DefaultRV32Config.fir@192514.4]
  assign _T_235 = ~tlb_io_req_ready; // @[DCache.scala 234:9:freechips.rocketchip.system.DefaultRV32Config.fir@192530.4]
  assign _T_236 = ~tlb_io_ptw_resp_valid; // @[DCache.scala 234:30:freechips.rocketchip.system.DefaultRV32Config.fir@192531.4]
  assign _T_237 = _T_235 & _T_236; // @[DCache.scala 234:27:freechips.rocketchip.system.DefaultRV32Config.fir@192532.4]
  assign _T_238 = ~io_cpu_req_bits_phys; // @[DCache.scala 234:56:freechips.rocketchip.system.DefaultRV32Config.fir@192533.4]
  assign _T_239 = _T_237 & _T_238; // @[DCache.scala 234:53:freechips.rocketchip.system.DefaultRV32Config.fir@192534.4]
  assign _GEN_31 = _T_239 ? 1'h0 : _GEN_30; // @[DCache.scala 234:79:freechips.rocketchip.system.DefaultRV32Config.fir@192535.4]
  assign s1_paddr = {tlb_io_resp_paddr[31:12],s1_req_addr[11:0]}; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@192570.4]
  assign s1_victim_way = _T_15[1:0]; // @[package.scala 138:13:freechips.rocketchip.system.DefaultRV32Config.fir@192571.4]
  assign _T_258 = metaArb_io_out_valid & metaArb_io_out_bits_write; // @[DCache.scala 262:27:freechips.rocketchip.system.DefaultRV32Config.fir@192575.4]
  assign _T_266 = tag_array_RW0_rdata_0; // @[:freechips.rocketchip.system.DefaultRV32Config.fir@192614.4 :freechips.rocketchip.system.DefaultRV32Config.fir@192616.4]
  assign s1_meta_uncorrected_0_tag = _T_266[19:0]; // @[DCache.scala 267:80:freechips.rocketchip.system.DefaultRV32Config.fir@192617.4]
  assign s1_meta_uncorrected_0_coh_state = _T_266[21:20]; // @[DCache.scala 267:80:freechips.rocketchip.system.DefaultRV32Config.fir@192619.4]
  assign _T_269 = tag_array_RW0_rdata_1; // @[:freechips.rocketchip.system.DefaultRV32Config.fir@192623.4 :freechips.rocketchip.system.DefaultRV32Config.fir@192625.4]
  assign s1_meta_uncorrected_1_tag = _T_269[19:0]; // @[DCache.scala 267:80:freechips.rocketchip.system.DefaultRV32Config.fir@192626.4]
  assign s1_meta_uncorrected_1_coh_state = _T_269[21:20]; // @[DCache.scala 267:80:freechips.rocketchip.system.DefaultRV32Config.fir@192628.4]
  assign _T_272 = tag_array_RW0_rdata_2; // @[:freechips.rocketchip.system.DefaultRV32Config.fir@192632.4 :freechips.rocketchip.system.DefaultRV32Config.fir@192634.4]
  assign s1_meta_uncorrected_2_tag = _T_272[19:0]; // @[DCache.scala 267:80:freechips.rocketchip.system.DefaultRV32Config.fir@192635.4]
  assign s1_meta_uncorrected_2_coh_state = _T_272[21:20]; // @[DCache.scala 267:80:freechips.rocketchip.system.DefaultRV32Config.fir@192637.4]
  assign _T_275 = tag_array_RW0_rdata_3; // @[:freechips.rocketchip.system.DefaultRV32Config.fir@192641.4 :freechips.rocketchip.system.DefaultRV32Config.fir@192643.4]
  assign s1_meta_uncorrected_3_tag = _T_275[19:0]; // @[DCache.scala 267:80:freechips.rocketchip.system.DefaultRV32Config.fir@192644.4]
  assign s1_meta_uncorrected_3_coh_state = _T_275[21:20]; // @[DCache.scala 267:80:freechips.rocketchip.system.DefaultRV32Config.fir@192646.4]
  assign s1_tag = s1_paddr[31:12]; // @[DCache.scala 268:29:freechips.rocketchip.system.DefaultRV32Config.fir@192648.4]
  assign _T_278 = s1_meta_uncorrected_0_coh_state > 2'h0; // @[Metadata.scala 50:45:freechips.rocketchip.system.DefaultRV32Config.fir@192649.4]
  assign _T_279 = s1_meta_uncorrected_0_tag == s1_tag; // @[DCache.scala 269:83:freechips.rocketchip.system.DefaultRV32Config.fir@192650.4]
  assign _T_280 = _T_278 & _T_279; // @[DCache.scala 269:74:freechips.rocketchip.system.DefaultRV32Config.fir@192651.4]
  assign _T_281 = s1_meta_uncorrected_1_coh_state > 2'h0; // @[Metadata.scala 50:45:freechips.rocketchip.system.DefaultRV32Config.fir@192652.4]
  assign _T_282 = s1_meta_uncorrected_1_tag == s1_tag; // @[DCache.scala 269:83:freechips.rocketchip.system.DefaultRV32Config.fir@192653.4]
  assign _T_283 = _T_281 & _T_282; // @[DCache.scala 269:74:freechips.rocketchip.system.DefaultRV32Config.fir@192654.4]
  assign _T_284 = s1_meta_uncorrected_2_coh_state > 2'h0; // @[Metadata.scala 50:45:freechips.rocketchip.system.DefaultRV32Config.fir@192655.4]
  assign _T_285 = s1_meta_uncorrected_2_tag == s1_tag; // @[DCache.scala 269:83:freechips.rocketchip.system.DefaultRV32Config.fir@192656.4]
  assign _T_286 = _T_284 & _T_285; // @[DCache.scala 269:74:freechips.rocketchip.system.DefaultRV32Config.fir@192657.4]
  assign _T_287 = s1_meta_uncorrected_3_coh_state > 2'h0; // @[Metadata.scala 50:45:freechips.rocketchip.system.DefaultRV32Config.fir@192658.4]
  assign _T_288 = s1_meta_uncorrected_3_tag == s1_tag; // @[DCache.scala 269:83:freechips.rocketchip.system.DefaultRV32Config.fir@192659.4]
  assign _T_289 = _T_287 & _T_288; // @[DCache.scala 269:74:freechips.rocketchip.system.DefaultRV32Config.fir@192660.4]
  assign s1_meta_hit_way = {_T_289,_T_286,_T_283,_T_280}; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@192663.4]
  assign _T_296 = _T_279 ? s1_meta_uncorrected_0_coh_state : 2'h0; // @[DCache.scala 271:41:freechips.rocketchip.system.DefaultRV32Config.fir@192670.4]
  assign _T_300 = _T_282 ? s1_meta_uncorrected_1_coh_state : 2'h0; // @[DCache.scala 271:41:freechips.rocketchip.system.DefaultRV32Config.fir@192674.4]
  assign _T_304 = _T_285 ? s1_meta_uncorrected_2_coh_state : 2'h0; // @[DCache.scala 271:41:freechips.rocketchip.system.DefaultRV32Config.fir@192678.4]
  assign _T_308 = _T_288 ? s1_meta_uncorrected_3_coh_state : 2'h0; // @[DCache.scala 271:41:freechips.rocketchip.system.DefaultRV32Config.fir@192682.4]
  assign _T_309 = _T_296 | _T_300; // @[DCache.scala 272:19:freechips.rocketchip.system.DefaultRV32Config.fir@192683.4]
  assign _T_310 = _T_309 | _T_304; // @[DCache.scala 272:19:freechips.rocketchip.system.DefaultRV32Config.fir@192684.4]
  assign s1_meta_hit_state_state = _T_310 | _T_308; // @[DCache.scala 272:19:freechips.rocketchip.system.DefaultRV32Config.fir@192685.4]
  assign _T_316 = s1_victim_way == 2'h1; // @[package.scala 32:86:freechips.rocketchip.system.DefaultRV32Config.fir@192695.4]
  assign _T_318 = s1_victim_way == 2'h2; // @[package.scala 32:86:freechips.rocketchip.system.DefaultRV32Config.fir@192697.4]
  assign _T_320 = s1_victim_way == 2'h3; // @[package.scala 32:86:freechips.rocketchip.system.DefaultRV32Config.fir@192699.4]
  assign s2_hit_valid = s2_hit_state_state > 2'h0; // @[Metadata.scala 50:45:freechips.rocketchip.system.DefaultRV32Config.fir@193008.4]
  assign _T_633 = 4'h1 << _T_632; // @[OneHot.scala 58:35:freechips.rocketchip.system.DefaultRV32Config.fir@193190.4]
  assign s2_victim_way = s2_hit_valid ? s2_hit_way : _T_633; // @[DCache.scala 383:26:freechips.rocketchip.system.DefaultRV32Config.fir@193191.4]
  assign releaseWay = _T_2412 ? s2_victim_way : s2_probe_way; // @[DCache.scala 783:81:freechips.rocketchip.system.DefaultRV32Config.fir@195510.4]
  assign _T_321 = inWriteback ? releaseWay : s1_meta_hit_way; // @[DCache.scala 275:61:freechips.rocketchip.system.DefaultRV32Config.fir@192701.4]
  assign _T_326 = {auto_out_d_bits_data[15:8],auto_out_d_bits_data[7:0]}; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@192709.4]
  assign _T_327 = {auto_out_d_bits_data[31:24],auto_out_d_bits_data[23:16]}; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@192710.4]
  assign _T_328 = {auto_out_d_bits_data[31:24],auto_out_d_bits_data[23:16],auto_out_d_bits_data[15:8],auto_out_d_bits_data[7:0]}; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@192711.4]
  assign _T_347 = s1_valid_masked & _T_53; // @[DCache.scala 281:28:freechips.rocketchip.system.DefaultRV32Config.fir@192741.4]
  assign _T_348 = ~_T_347; // @[DCache.scala 281:10:freechips.rocketchip.system.DefaultRV32Config.fir@192742.4]
  assign _T_349 = ~io_cpu_s1_data_mask; // @[DCache.scala 281:71:freechips.rocketchip.system.DefaultRV32Config.fir@192743.4]
  assign _T_350 = s1_mask_xwr | _T_349; // @[DCache.scala 281:69:freechips.rocketchip.system.DefaultRV32Config.fir@192744.4]
  assign _T_351 = &_T_350; // @[DCache.scala 281:93:freechips.rocketchip.system.DefaultRV32Config.fir@192745.4]
  assign _T_352 = _T_348 | _T_351; // @[DCache.scala 281:53:freechips.rocketchip.system.DefaultRV32Config.fir@192746.4]
  assign _T_354 = _T_352 | reset; // @[DCache.scala 281:9:freechips.rocketchip.system.DefaultRV32Config.fir@192748.4]
  assign _T_355 = ~_T_354; // @[DCache.scala 281:9:freechips.rocketchip.system.DefaultRV32Config.fir@192749.4]
  assign _T_356 = ~s1_sfence; // @[DCache.scala 283:46:freechips.rocketchip.system.DefaultRV32Config.fir@192754.4]
  assign _T_357 = s1_valid_masked & _T_356; // @[DCache.scala 283:43:freechips.rocketchip.system.DefaultRV32Config.fir@192755.4]
  assign _T_369 = s2_req_cmd == 5'h5; // @[DCache.scala 292:37:freechips.rocketchip.system.DefaultRV32Config.fir@192779.4]
  assign s2_cmd_flush_line = _T_369 & s2_req_size[0]; // @[DCache.scala 293:54:freechips.rocketchip.system.DefaultRV32Config.fir@192785.4]
  assign s2_vaddr = {_T_377[31:12],s2_req_addr[11:0]}; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@192804.4]
  assign s1_meta_clk_en = s1_valid_not_nacked | s1_probe; // @[DCache.scala 309:62:freechips.rocketchip.system.DefaultRV32Config.fir@192855.4]
  assign s2_meta_corrected_3_tag = _T_449[19:0]; // @[DCache.scala 313:99:freechips.rocketchip.system.DefaultRV32Config.fir@192943.4]
  assign s2_meta_corrected_3_coh_state = _T_449[21:20]; // @[DCache.scala 313:99:freechips.rocketchip.system.DefaultRV32Config.fir@192945.4]
  assign _T_455 = s1_valid | inWriteback; // @[DCache.scala 318:23:freechips.rocketchip.system.DefaultRV32Config.fir@192951.4]
  assign en = _T_455 | io_cpu_replay_next; // @[DCache.scala 318:38:freechips.rocketchip.system.DefaultRV32Config.fir@192952.4]
  assign _T_456 = ~s1_did_read; // @[DCache.scala 319:64:freechips.rocketchip.system.DefaultRV32Config.fir@192953.4]
  assign _T_457 = _T_456 ? 1'h0 : 1'h1; // @[DCache.scala 319:63:freechips.rocketchip.system.DefaultRV32Config.fir@192954.4]
  assign word_en = inWriteback | _T_457; // @[DCache.scala 319:22:freechips.rocketchip.system.DefaultRV32Config.fir@192955.4]
  assign s1_all_data_ways_0 = data_io_resp_0; // @[DCache.scala 277:29:freechips.rocketchip.system.DefaultRV32Config.fir@192714.4 DCache.scala 277:29:freechips.rocketchip.system.DefaultRV32Config.fir@192716.4]
  assign s1_all_data_ways_1 = data_io_resp_1; // @[DCache.scala 277:29:freechips.rocketchip.system.DefaultRV32Config.fir@192714.4 DCache.scala 277:29:freechips.rocketchip.system.DefaultRV32Config.fir@192717.4]
  assign s1_all_data_ways_2 = data_io_resp_2; // @[DCache.scala 277:29:freechips.rocketchip.system.DefaultRV32Config.fir@192714.4 DCache.scala 277:29:freechips.rocketchip.system.DefaultRV32Config.fir@192718.4]
  assign s1_all_data_ways_3 = data_io_resp_3; // @[DCache.scala 277:29:freechips.rocketchip.system.DefaultRV32Config.fir@192714.4 DCache.scala 277:29:freechips.rocketchip.system.DefaultRV32Config.fir@192719.4]
  assign _T_458 = ~io_cpu_replay_next; // @[DCache.scala 329:28:freechips.rocketchip.system.DefaultRV32Config.fir@192961.4]
  assign s1_word_en = _T_458 ? word_en : 1'h1; // @[DCache.scala 329:27:freechips.rocketchip.system.DefaultRV32Config.fir@192962.4]
  assign grantIsUncachedData = auto_out_d_bits_opcode == 3'h1; // @[package.scala 15:47:freechips.rocketchip.system.DefaultRV32Config.fir@195063.4]
  assign _T_2333 = blockUncachedGrant | s1_valid; // @[DCache.scala 695:54:freechips.rocketchip.system.DefaultRV32Config.fir@195296.4]
  assign _T_2334 = grantIsUncachedData & _T_2333; // @[DCache.scala 695:31:freechips.rocketchip.system.DefaultRV32Config.fir@195297.4]
  assign grantIsRefill = auto_out_d_bits_opcode == 3'h5; // @[DCache.scala 609:29:freechips.rocketchip.system.DefaultRV32Config.fir@195081.4]
  assign _T_2247 = ~dataArb_io_in_1_ready; // @[DCache.scala 665:26:freechips.rocketchip.system.DefaultRV32Config.fir@195187.4]
  assign _T_2248 = grantIsRefill & _T_2247; // @[DCache.scala 665:23:freechips.rocketchip.system.DefaultRV32Config.fir@195188.4]
  assign _T_2201 = auto_out_d_bits_opcode == 3'h4; // @[package.scala 15:47:freechips.rocketchip.system.DefaultRV32Config.fir@195077.4]
  assign grantIsCached = _T_2201 | grantIsRefill; // @[package.scala 64:59:freechips.rocketchip.system.DefaultRV32Config.fir@195079.4]
  assign d_first = _T_2177 == 10'h0; // @[Edges.scala 232:25:freechips.rocketchip.system.DefaultRV32Config.fir@195046.4]
  assign _T_2209 = ~d_first; // @[DCache.scala 614:41:freechips.rocketchip.system.DefaultRV32Config.fir@195094.4]
  assign _T_2210 = _T_2209 | auto_out_e_ready; // @[DCache.scala 614:50:freechips.rocketchip.system.DefaultRV32Config.fir@195095.4]
  assign canAcceptCachedGrant = ~_T_2412; // @[DCache.scala 613:30:freechips.rocketchip.system.DefaultRV32Config.fir@195093.4]
  assign _T_2211 = _T_2210 & canAcceptCachedGrant; // @[DCache.scala 614:69:freechips.rocketchip.system.DefaultRV32Config.fir@195096.4]
  assign _T_2212 = grantIsCached ? _T_2211 : 1'h1; // @[DCache.scala 614:24:freechips.rocketchip.system.DefaultRV32Config.fir@195097.4]
  assign _GEN_228 = _T_2248 ? 1'h0 : _T_2212; // @[DCache.scala 665:51:freechips.rocketchip.system.DefaultRV32Config.fir@195189.4]
  assign tl_out__d_ready = _T_2334 ? 1'h0 : _GEN_228; // @[DCache.scala 695:68:freechips.rocketchip.system.DefaultRV32Config.fir@195298.4]
  assign _T_2217 = tl_out__d_ready & auto_out_d_valid; // @[Decoupled.scala 40:37:freechips.rocketchip.system.DefaultRV32Config.fir@195105.4]
  assign _T_2186 = auto_out_d_bits_opcode == 3'h0; // @[package.scala 15:47:freechips.rocketchip.system.DefaultRV32Config.fir@195059.4]
  assign _T_2188 = grantIsUncachedData | _T_2186; // @[package.scala 64:59:freechips.rocketchip.system.DefaultRV32Config.fir@195061.4]
  assign _T_2187 = auto_out_d_bits_opcode == 3'h2; // @[package.scala 15:47:freechips.rocketchip.system.DefaultRV32Config.fir@195060.4]
  assign grantIsUncached = _T_2188 | _T_2187; // @[package.scala 64:59:freechips.rocketchip.system.DefaultRV32Config.fir@195062.4]
  assign _GEN_184 = grantIsUncachedData ? 5'h10 : {{1'd0}, _T_321}; // @[DCache.scala 634:34:freechips.rocketchip.system.DefaultRV32Config.fir@195137.10]
  assign _GEN_193 = grantIsUncached ? _GEN_184 : {{1'd0}, _T_321}; // @[DCache.scala 627:35:freechips.rocketchip.system.DefaultRV32Config.fir@195124.8]
  assign _GEN_206 = grantIsCached ? {{1'd0}, _T_321} : _GEN_193; // @[DCache.scala 618:26:freechips.rocketchip.system.DefaultRV32Config.fir@195107.6]
  assign s1_data_way = _T_2217 ? _GEN_206 : {{1'd0}, _T_321}; // @[DCache.scala 617:26:freechips.rocketchip.system.DefaultRV32Config.fir@195106.4]
  assign _T_460 = s1_word_en ? s1_data_way : 5'h0; // @[DCache.scala 331:28:freechips.rocketchip.system.DefaultRV32Config.fir@192964.4]
  assign _T_466 = _T_460[0] ? s1_all_data_ways_0 : 32'h0; // @[Mux.scala 27:72:freechips.rocketchip.system.DefaultRV32Config.fir@192970.4]
  assign _T_467 = _T_460[1] ? s1_all_data_ways_1 : 32'h0; // @[Mux.scala 27:72:freechips.rocketchip.system.DefaultRV32Config.fir@192971.4]
  assign _T_468 = _T_460[2] ? s1_all_data_ways_2 : 32'h0; // @[Mux.scala 27:72:freechips.rocketchip.system.DefaultRV32Config.fir@192972.4]
  assign _T_469 = _T_460[3] ? s1_all_data_ways_3 : 32'h0; // @[Mux.scala 27:72:freechips.rocketchip.system.DefaultRV32Config.fir@192973.4]
  assign _T_470 = _T_460[4] ? _T_328 : 32'h0; // @[Mux.scala 27:72:freechips.rocketchip.system.DefaultRV32Config.fir@192974.4]
  assign _T_471 = _T_466 | _T_467; // @[Mux.scala 27:72:freechips.rocketchip.system.DefaultRV32Config.fir@192975.4]
  assign _T_472 = _T_471 | _T_468; // @[Mux.scala 27:72:freechips.rocketchip.system.DefaultRV32Config.fir@192976.4]
  assign _T_473 = _T_472 | _T_469; // @[Mux.scala 27:72:freechips.rocketchip.system.DefaultRV32Config.fir@192977.4]
  assign _T_474 = _T_473 | _T_470; // @[Mux.scala 27:72:freechips.rocketchip.system.DefaultRV32Config.fir@192978.4]
  assign _T_599 = {s2_data[15:8],s2_data[7:0]}; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@193138.4]
  assign _T_600 = {s2_data[31:24],s2_data[23:16]}; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@193139.4]
  assign s2_data_corrected = {s2_data[31:24],s2_data[23:16],s2_data[15:8],s2_data[7:0]}; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@193140.4]
  assign s2_valid_flush_line = s2_valid_hit_maybe_flush_pre_data_ecc_and_waw & s2_cmd_flush_line; // @[DCache.scala 371:75:freechips.rocketchip.system.DefaultRV32Config.fir@193150.4]
  assign _T_610 = s2_valid_masked & s2_readwrite; // @[DCache.scala 375:39:freechips.rocketchip.system.DefaultRV32Config.fir@193157.4]
  assign _T_612 = _T_610 & _T_603; // @[DCache.scala 375:55:freechips.rocketchip.system.DefaultRV32Config.fir@193159.4]
  assign _T_613 = ~s2_hit; // @[DCache.scala 375:76:freechips.rocketchip.system.DefaultRV32Config.fir@193160.4]
  assign s2_valid_miss = _T_612 & _T_613; // @[DCache.scala 375:73:freechips.rocketchip.system.DefaultRV32Config.fir@193161.4]
  assign s2_uncached = ~s2_pma_cacheable; // @[DCache.scala 376:21:freechips.rocketchip.system.DefaultRV32Config.fir@193162.4]
  assign _T_619 = ~s2_uncached; // @[DCache.scala 377:47:freechips.rocketchip.system.DefaultRV32Config.fir@193168.4]
  assign _T_620 = s2_valid_miss & _T_619; // @[DCache.scala 377:44:freechips.rocketchip.system.DefaultRV32Config.fir@193169.4]
  assign _T_621 = |uncachedInFlight_0; // @[DCache.scala 377:88:freechips.rocketchip.system.DefaultRV32Config.fir@193170.4]
  assign _T_622 = ~_T_621; // @[DCache.scala 377:63:freechips.rocketchip.system.DefaultRV32Config.fir@193171.4]
  assign s2_valid_cached_miss = _T_620 & _T_622; // @[DCache.scala 377:60:freechips.rocketchip.system.DefaultRV32Config.fir@193172.4]
  assign s2_want_victimize = s2_valid_cached_miss | s2_valid_flush_line; // @[DCache.scala 379:79:freechips.rocketchip.system.DefaultRV32Config.fir@193173.4]
  assign _T_628 = s2_valid_miss & s2_uncached; // @[DCache.scala 382:49:freechips.rocketchip.system.DefaultRV32Config.fir@193181.4]
  assign _T_629 = &uncachedInFlight_0; // @[DCache.scala 382:92:freechips.rocketchip.system.DefaultRV32Config.fir@193182.4]
  assign _T_630 = ~_T_629; // @[DCache.scala 382:67:freechips.rocketchip.system.DefaultRV32Config.fir@193183.4]
  assign s2_valid_uncached_pending = _T_628 & _T_630; // @[DCache.scala 382:64:freechips.rocketchip.system.DefaultRV32Config.fir@193184.4]
  assign s2_victim_tag = s2_valid_flush_line ? s2_req_addr[31:12] : _T_637; // @[DCache.scala 384:26:freechips.rocketchip.system.DefaultRV32Config.fir@193199.4]
  assign s2_victim_state_state = s2_hit_valid ? s2_hit_state_state : _T_639_state; // @[DCache.scala 385:28:freechips.rocketchip.system.DefaultRV32Config.fir@193205.4]
  assign _T_655 = _T_653 ? 3'h5 : 3'h0; // @[Misc.scala 37:36:freechips.rocketchip.system.DefaultRV32Config.fir@193221.4]
  assign _T_659 = _T_657 ? 3'h2 : _T_655; // @[Misc.scala 37:36:freechips.rocketchip.system.DefaultRV32Config.fir@193225.4]
  assign _T_663 = _T_661 ? 3'h1 : _T_659; // @[Misc.scala 37:36:freechips.rocketchip.system.DefaultRV32Config.fir@193229.4]
  assign _T_667 = _T_665 ? 3'h1 : _T_663; // @[Misc.scala 37:36:freechips.rocketchip.system.DefaultRV32Config.fir@193233.4]
  assign _T_671 = _T_669 ? 3'h5 : _T_667; // @[Misc.scala 37:36:freechips.rocketchip.system.DefaultRV32Config.fir@193237.4]
  assign _T_675 = _T_673 ? 3'h4 : _T_671; // @[Misc.scala 37:36:freechips.rocketchip.system.DefaultRV32Config.fir@193241.4]
  assign _T_676 = _T_673 ? 2'h1 : 2'h0; // @[Misc.scala 37:63:freechips.rocketchip.system.DefaultRV32Config.fir@193242.4]
  assign _T_679 = _T_677 ? 3'h0 : _T_675; // @[Misc.scala 37:36:freechips.rocketchip.system.DefaultRV32Config.fir@193245.4]
  assign _T_680 = _T_677 ? 2'h1 : _T_676; // @[Misc.scala 37:63:freechips.rocketchip.system.DefaultRV32Config.fir@193246.4]
  assign _T_683 = _T_681 ? 3'h0 : _T_679; // @[Misc.scala 37:36:freechips.rocketchip.system.DefaultRV32Config.fir@193249.4]
  assign _T_684 = _T_681 ? 2'h1 : _T_680; // @[Misc.scala 37:63:freechips.rocketchip.system.DefaultRV32Config.fir@193250.4]
  assign _T_687 = _T_685 ? 3'h5 : _T_683; // @[Misc.scala 37:36:freechips.rocketchip.system.DefaultRV32Config.fir@193253.4]
  assign _T_688 = _T_685 ? 2'h0 : _T_684; // @[Misc.scala 37:63:freechips.rocketchip.system.DefaultRV32Config.fir@193254.4]
  assign _T_691 = _T_689 ? 3'h4 : _T_687; // @[Misc.scala 37:36:freechips.rocketchip.system.DefaultRV32Config.fir@193257.4]
  assign _T_692 = _T_689 ? 2'h1 : _T_688; // @[Misc.scala 37:63:freechips.rocketchip.system.DefaultRV32Config.fir@193258.4]
  assign _T_695 = _T_693 ? 3'h3 : _T_691; // @[Misc.scala 37:36:freechips.rocketchip.system.DefaultRV32Config.fir@193261.4]
  assign _T_696 = _T_693 ? 2'h2 : _T_692; // @[Misc.scala 37:63:freechips.rocketchip.system.DefaultRV32Config.fir@193262.4]
  assign s2_report_param = _T_697 ? 3'h3 : _T_695; // @[Misc.scala 37:36:freechips.rocketchip.system.DefaultRV32Config.fir@193265.4]
  assign probeNewCoh_state = _T_697 ? 2'h2 : _T_696; // @[Misc.scala 37:63:freechips.rocketchip.system.DefaultRV32Config.fir@193266.4]
  assign _T_705 = {2'h2,s2_victim_state_state}; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@193276.4]
  assign _T_718 = 4'h8 == _T_705; // @[Misc.scala 55:20:freechips.rocketchip.system.DefaultRV32Config.fir@193289.4]
  assign _T_720 = _T_718 ? 3'h5 : 3'h0; // @[Misc.scala 37:36:freechips.rocketchip.system.DefaultRV32Config.fir@193291.4]
  assign _T_722 = 4'h9 == _T_705; // @[Misc.scala 55:20:freechips.rocketchip.system.DefaultRV32Config.fir@193293.4]
  assign _T_724 = _T_722 ? 3'h2 : _T_720; // @[Misc.scala 37:36:freechips.rocketchip.system.DefaultRV32Config.fir@193295.4]
  assign _T_726 = 4'ha == _T_705; // @[Misc.scala 55:20:freechips.rocketchip.system.DefaultRV32Config.fir@193297.4]
  assign _T_728 = _T_726 ? 3'h1 : _T_724; // @[Misc.scala 37:36:freechips.rocketchip.system.DefaultRV32Config.fir@193299.4]
  assign _T_730 = 4'hb == _T_705; // @[Misc.scala 55:20:freechips.rocketchip.system.DefaultRV32Config.fir@193301.4]
  assign _T_732 = _T_730 ? 3'h1 : _T_728; // @[Misc.scala 37:36:freechips.rocketchip.system.DefaultRV32Config.fir@193303.4]
  assign _T_734 = 4'h4 == _T_705; // @[Misc.scala 55:20:freechips.rocketchip.system.DefaultRV32Config.fir@193305.4]
  assign _T_735 = _T_734 ? 1'h0 : _T_730; // @[Misc.scala 37:9:freechips.rocketchip.system.DefaultRV32Config.fir@193306.4]
  assign _T_736 = _T_734 ? 3'h5 : _T_732; // @[Misc.scala 37:36:freechips.rocketchip.system.DefaultRV32Config.fir@193307.4]
  assign _T_738 = 4'h5 == _T_705; // @[Misc.scala 55:20:freechips.rocketchip.system.DefaultRV32Config.fir@193309.4]
  assign _T_739 = _T_738 ? 1'h0 : _T_735; // @[Misc.scala 37:9:freechips.rocketchip.system.DefaultRV32Config.fir@193310.4]
  assign _T_740 = _T_738 ? 3'h4 : _T_736; // @[Misc.scala 37:36:freechips.rocketchip.system.DefaultRV32Config.fir@193311.4]
  assign _T_741 = _T_738 ? 2'h1 : 2'h0; // @[Misc.scala 37:63:freechips.rocketchip.system.DefaultRV32Config.fir@193312.4]
  assign _T_742 = 4'h6 == _T_705; // @[Misc.scala 55:20:freechips.rocketchip.system.DefaultRV32Config.fir@193313.4]
  assign _T_743 = _T_742 ? 1'h0 : _T_739; // @[Misc.scala 37:9:freechips.rocketchip.system.DefaultRV32Config.fir@193314.4]
  assign _T_744 = _T_742 ? 3'h0 : _T_740; // @[Misc.scala 37:36:freechips.rocketchip.system.DefaultRV32Config.fir@193315.4]
  assign _T_745 = _T_742 ? 2'h1 : _T_741; // @[Misc.scala 37:63:freechips.rocketchip.system.DefaultRV32Config.fir@193316.4]
  assign _T_746 = 4'h7 == _T_705; // @[Misc.scala 55:20:freechips.rocketchip.system.DefaultRV32Config.fir@193317.4]
  assign _T_747 = _T_746 | _T_743; // @[Misc.scala 37:9:freechips.rocketchip.system.DefaultRV32Config.fir@193318.4]
  assign _T_748 = _T_746 ? 3'h0 : _T_744; // @[Misc.scala 37:36:freechips.rocketchip.system.DefaultRV32Config.fir@193319.4]
  assign _T_749 = _T_746 ? 2'h1 : _T_745; // @[Misc.scala 37:63:freechips.rocketchip.system.DefaultRV32Config.fir@193320.4]
  assign _T_750 = 4'h0 == _T_705; // @[Misc.scala 55:20:freechips.rocketchip.system.DefaultRV32Config.fir@193321.4]
  assign _T_751 = _T_750 ? 1'h0 : _T_747; // @[Misc.scala 37:9:freechips.rocketchip.system.DefaultRV32Config.fir@193322.4]
  assign _T_752 = _T_750 ? 3'h5 : _T_748; // @[Misc.scala 37:36:freechips.rocketchip.system.DefaultRV32Config.fir@193323.4]
  assign _T_753 = _T_750 ? 2'h0 : _T_749; // @[Misc.scala 37:63:freechips.rocketchip.system.DefaultRV32Config.fir@193324.4]
  assign _T_754 = 4'h1 == _T_705; // @[Misc.scala 55:20:freechips.rocketchip.system.DefaultRV32Config.fir@193325.4]
  assign _T_755 = _T_754 ? 1'h0 : _T_751; // @[Misc.scala 37:9:freechips.rocketchip.system.DefaultRV32Config.fir@193326.4]
  assign _T_756 = _T_754 ? 3'h4 : _T_752; // @[Misc.scala 37:36:freechips.rocketchip.system.DefaultRV32Config.fir@193327.4]
  assign _T_757 = _T_754 ? 2'h1 : _T_753; // @[Misc.scala 37:63:freechips.rocketchip.system.DefaultRV32Config.fir@193328.4]
  assign _T_758 = 4'h2 == _T_705; // @[Misc.scala 55:20:freechips.rocketchip.system.DefaultRV32Config.fir@193329.4]
  assign _T_759 = _T_758 ? 1'h0 : _T_755; // @[Misc.scala 37:9:freechips.rocketchip.system.DefaultRV32Config.fir@193330.4]
  assign _T_760 = _T_758 ? 3'h3 : _T_756; // @[Misc.scala 37:36:freechips.rocketchip.system.DefaultRV32Config.fir@193331.4]
  assign _T_761 = _T_758 ? 2'h2 : _T_757; // @[Misc.scala 37:63:freechips.rocketchip.system.DefaultRV32Config.fir@193332.4]
  assign _T_762 = 4'h3 == _T_705; // @[Misc.scala 55:20:freechips.rocketchip.system.DefaultRV32Config.fir@193333.4]
  assign s2_victim_dirty = _T_762 | _T_759; // @[Misc.scala 37:9:freechips.rocketchip.system.DefaultRV32Config.fir@193334.4]
  assign s2_shrink_param = _T_762 ? 3'h3 : _T_760; // @[Misc.scala 37:36:freechips.rocketchip.system.DefaultRV32Config.fir@193335.4]
  assign voluntaryNewCoh_state = _T_762 ? 2'h2 : _T_761; // @[Misc.scala 37:63:freechips.rocketchip.system.DefaultRV32Config.fir@193336.4]
  assign s2_dont_nack_uncached = s2_valid_uncached_pending & auto_out_a_ready; // @[DCache.scala 391:57:freechips.rocketchip.system.DefaultRV32Config.fir@193342.4]
  assign _T_775 = s2_req_cmd == 5'h17; // @[DCache.scala 395:17:freechips.rocketchip.system.DefaultRV32Config.fir@193353.4]
  assign s2_dont_nack_misc = _T_604 & _T_775; // @[DCache.scala 392:61:freechips.rocketchip.system.DefaultRV32Config.fir@193355.4]
  assign _T_777 = ~s2_dont_nack_uncached; // @[DCache.scala 396:41:freechips.rocketchip.system.DefaultRV32Config.fir@193356.4]
  assign _T_778 = s2_valid_no_xcpt & _T_777; // @[DCache.scala 396:38:freechips.rocketchip.system.DefaultRV32Config.fir@193357.4]
  assign _T_779 = ~s2_dont_nack_misc; // @[DCache.scala 396:67:freechips.rocketchip.system.DefaultRV32Config.fir@193358.4]
  assign _T_780 = _T_778 & _T_779; // @[DCache.scala 396:64:freechips.rocketchip.system.DefaultRV32Config.fir@193359.4]
  assign _T_781 = ~s2_valid_hit_pre_data_ecc_and_waw; // @[DCache.scala 396:89:freechips.rocketchip.system.DefaultRV32Config.fir@193360.4]
  assign _T_792 = s2_valid_masked | s2_probe; // @[DCache.scala 401:93:freechips.rocketchip.system.DefaultRV32Config.fir@193376.4]
  assign _T_808 = {metaArb_io_in_1_bits_idx, 6'h0}; // @[DCache.scala 405:98:freechips.rocketchip.system.DefaultRV32Config.fir@193396.4]
  assign new_meta_coh_state = pma_checker__T_2026 ? 2'h0 : s2_meta_corrected_3_coh_state; // @[DCache.scala 408:40:freechips.rocketchip.system.DefaultRV32Config.fir@193402.4]
  assign _T_823 = lrscCount > 7'h0; // @[DCache.scala 425:34:freechips.rocketchip.system.DefaultRV32Config.fir@193434.4]
  assign _T_824 = ~lrscValid; // @[DCache.scala 425:41:freechips.rocketchip.system.DefaultRV32Config.fir@193435.4]
  assign lrscBackingOff = _T_823 & _T_824; // @[DCache.scala 425:38:freechips.rocketchip.system.DefaultRV32Config.fir@193436.4]
  assign lrscAddrMatch = lrscAddr == s2_req_addr[31:6]; // @[DCache.scala 427:32:freechips.rocketchip.system.DefaultRV32Config.fir@193439.4]
  assign _T_826 = lrscValid & lrscAddrMatch; // @[DCache.scala 428:41:freechips.rocketchip.system.DefaultRV32Config.fir@193440.4]
  assign _T_827 = ~_T_826; // @[DCache.scala 428:29:freechips.rocketchip.system.DefaultRV32Config.fir@193441.4]
  assign s2_sc_fail = _T_405 & _T_827; // @[DCache.scala 428:26:freechips.rocketchip.system.DefaultRV32Config.fir@193442.4]
  assign _T_828 = s2_valid_hit_pre_data_ecc_and_waw & _T_525; // @[DCache.scala 429:23:freechips.rocketchip.system.DefaultRV32Config.fir@193443.4]
  assign _T_830 = _T_828 & _T_79; // @[DCache.scala 429:32:freechips.rocketchip.system.DefaultRV32Config.fir@193445.4]
  assign _T_831 = _T_830 | s2_valid_cached_miss; // @[DCache.scala 429:54:freechips.rocketchip.system.DefaultRV32Config.fir@193446.4]
  assign _T_838 = lrscCount - 7'h1; // @[DCache.scala 433:49:freechips.rocketchip.system.DefaultRV32Config.fir@193458.6]
  assign _T_839 = s2_valid_masked & lrscValid; // @[DCache.scala 434:29:freechips.rocketchip.system.DefaultRV32Config.fir@193461.4]
  assign _T_847 = s1_valid_not_nacked & s1_write; // @[DCache.scala 443:63:freechips.rocketchip.system.DefaultRV32Config.fir@193478.4]
  assign _T_901 = s1_write & _T_53; // @[DCache.scala 1086:23:freechips.rocketchip.system.DefaultRV32Config.fir@193555.4]
  assign _T_902 = s1_read | _T_901; // @[DCache.scala 1085:21:freechips.rocketchip.system.DefaultRV32Config.fir@193556.4]
  assign _T_906 = s2_valid_hit_pre_data_ecc_and_waw & s2_write; // @[DCache.scala 441:46:freechips.rocketchip.system.DefaultRV32Config.fir@193565.4]
  assign _T_907 = ~s2_sc_fail; // @[DCache.scala 441:61:freechips.rocketchip.system.DefaultRV32Config.fir@193566.4]
  assign _T_908 = _T_906 & _T_907; // @[DCache.scala 441:58:freechips.rocketchip.system.DefaultRV32Config.fir@193567.4]
  assign pstore_drain_opportunistic = ~_T_167; // @[DCache.scala 453:36:freechips.rocketchip.system.DefaultRV32Config.fir@193639.4]
  assign pstore_drain_on_miss = releaseInFlight | _T_976; // @[DCache.scala 454:46:freechips.rocketchip.system.DefaultRV32Config.fir@193645.4]
  assign pstore1_valid = _T_908 | pstore1_held; // @[DCache.scala 458:38:freechips.rocketchip.system.DefaultRV32Config.fir@193654.4]
  assign _T_984 = pstore1_valid_likely & pstore2_valid; // @[DCache.scala 460:54:freechips.rocketchip.system.DefaultRV32Config.fir@193657.4]
  assign _T_985 = s1_valid & s1_write; // @[DCache.scala 460:85:freechips.rocketchip.system.DefaultRV32Config.fir@193658.4]
  assign _T_986 = _T_985 | pstore1_rmw; // @[DCache.scala 460:98:freechips.rocketchip.system.DefaultRV32Config.fir@193659.4]
  assign pstore_drain_structural = _T_984 & _T_986; // @[DCache.scala 460:71:freechips.rocketchip.system.DefaultRV32Config.fir@193660.4]
  assign _T_990 = _T_906 | pstore1_held; // @[DCache.scala 457:96:freechips.rocketchip.system.DefaultRV32Config.fir@193664.4]
  assign _T_991 = _T_990 == pstore1_valid; // @[DCache.scala 461:63:freechips.rocketchip.system.DefaultRV32Config.fir@193665.4]
  assign _T_992 = pstore1_rmw | _T_991; // @[DCache.scala 461:22:freechips.rocketchip.system.DefaultRV32Config.fir@193666.4]
  assign _T_994 = _T_992 | reset; // @[DCache.scala 461:9:freechips.rocketchip.system.DefaultRV32Config.fir@193668.4]
  assign _T_995 = ~_T_994; // @[DCache.scala 461:9:freechips.rocketchip.system.DefaultRV32Config.fir@193669.4]
  assign _T_1004 = ~pstore1_rmw; // @[DCache.scala 469:44:freechips.rocketchip.system.DefaultRV32Config.fir@193683.4]
  assign _T_1005 = _T_990 & _T_1004; // @[DCache.scala 469:41:freechips.rocketchip.system.DefaultRV32Config.fir@193684.4]
  assign _T_1006 = _T_1005 | pstore2_valid; // @[DCache.scala 469:58:freechips.rocketchip.system.DefaultRV32Config.fir@193685.4]
  assign _T_1007 = pstore_drain_opportunistic | pstore_drain_on_miss; // @[DCache.scala 469:107:freechips.rocketchip.system.DefaultRV32Config.fir@193686.4]
  assign _T_1008 = _T_1006 & _T_1007; // @[DCache.scala 469:76:freechips.rocketchip.system.DefaultRV32Config.fir@193687.4]
  assign pstore_drain = pstore_drain_structural | _T_1008; // @[DCache.scala 468:48:freechips.rocketchip.system.DefaultRV32Config.fir@193688.4]
  assign _T_1018 = pstore1_valid & pstore2_valid; // @[DCache.scala 472:71:freechips.rocketchip.system.DefaultRV32Config.fir@193698.4]
  assign _T_1019 = ~pstore_drain; // @[DCache.scala 472:91:freechips.rocketchip.system.DefaultRV32Config.fir@193699.4]
  assign _T_1022 = pstore2_valid == pstore_drain; // @[DCache.scala 473:79:freechips.rocketchip.system.DefaultRV32Config.fir@193703.4]
  assign advance_pstore1 = pstore1_valid & _T_1022; // @[DCache.scala 473:61:freechips.rocketchip.system.DefaultRV32Config.fir@193704.4]
  assign _T_1024 = pstore2_valid & _T_1019; // @[DCache.scala 474:34:freechips.rocketchip.system.DefaultRV32Config.fir@193706.4]
  assign pstore1_storegen_data = amoalu_io_out; // @[:freechips.rocketchip.system.DefaultRV32Config.fir@193503.4 :freechips.rocketchip.system.DefaultRV32Config.fir@193505.4 DCache.scala 888:27:freechips.rocketchip.system.DefaultRV32Config.fir@195717.4]
  assign pstore2_storegen_data = {_T_1047,_T_1042,_T_1037,_T_1032}; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@193753.4]
  assign _T_1052 = ~pstore1_mask; // @[DCache.scala 485:37:freechips.rocketchip.system.DefaultRV32Config.fir@193759.6]
  assign _T_1054 = ~_T_1052; // @[DCache.scala 485:15:freechips.rocketchip.system.DefaultRV32Config.fir@193761.6]
  assign _T_1068 = pstore2_valid ? pstore2_addr : pstore1_addr; // @[DCache.scala 500:36:freechips.rocketchip.system.DefaultRV32Config.fir@193781.4]
  assign _T_1070 = pstore2_valid ? pstore2_storegen_data : pstore1_data; // @[DCache.scala 502:63:freechips.rocketchip.system.DefaultRV32Config.fir@193785.4]
  assign _T_1075 = {_T_1070[15:8],_T_1070[7:0]}; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@193790.4]
  assign _T_1076 = {_T_1070[31:24],_T_1070[23:16]}; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@193791.4]
  assign _T_1080 = pstore2_valid ? mask : pstore1_mask; // @[DCache.scala 504:47:freechips.rocketchip.system.DefaultRV32Config.fir@193797.4]
  assign _T_1085 = |_T_1080[0]; // @[DCache.scala 1076:66:freechips.rocketchip.system.DefaultRV32Config.fir@193802.4]
  assign _T_1086 = |_T_1080[1]; // @[DCache.scala 1076:66:freechips.rocketchip.system.DefaultRV32Config.fir@193803.4]
  assign _T_1087 = |_T_1080[2]; // @[DCache.scala 1076:66:freechips.rocketchip.system.DefaultRV32Config.fir@193804.4]
  assign _T_1088 = |_T_1080[3]; // @[DCache.scala 1076:66:freechips.rocketchip.system.DefaultRV32Config.fir@193805.4]
  assign _T_1089 = {_T_1086,_T_1085}; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@193806.4]
  assign _T_1090 = {_T_1088,_T_1087}; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@193807.4]
  assign _T_1190 = ~uncachedInFlight_0; // @[DCache.scala 524:34:freechips.rocketchip.system.DefaultRV32Config.fir@193916.4]
  assign _T_1191 = {_T_1190, 1'h0}; // @[DCache.scala 524:59:freechips.rocketchip.system.DefaultRV32Config.fir@193917.4]
  assign a_source = _T_1191[0] ? 1'h0 : 1'h1; // @[Mux.scala 47:69:freechips.rocketchip.system.DefaultRV32Config.fir@193920.4]
  assign acquire_address = {s2_req_addr[31:6], 6'h0}; // @[DCache.scala 525:49:freechips.rocketchip.system.DefaultRV32Config.fir@193922.4]
  assign a_mask = {{15'd0}, pstore1_mask}; // @[DCache.scala 529:29:freechips.rocketchip.system.DefaultRV32Config.fir@193924.4]
  assign _T_1250 = 2'h1 << s2_req_size[0]; // @[OneHot.scala 65:12:freechips.rocketchip.system.DefaultRV32Config.fir@193986.4]
  assign _T_1252 = _T_1250 | 2'h1; // @[Misc.scala 201:81:freechips.rocketchip.system.DefaultRV32Config.fir@193988.4]
  assign _T_1253 = s2_req_size >= 2'h2; // @[Misc.scala 205:21:freechips.rocketchip.system.DefaultRV32Config.fir@193989.4]
  assign _T_1256 = ~s2_req_addr[1]; // @[Misc.scala 210:20:freechips.rocketchip.system.DefaultRV32Config.fir@193992.4]
  assign _T_1258 = _T_1252[1] & _T_1256; // @[Misc.scala 214:38:freechips.rocketchip.system.DefaultRV32Config.fir@193994.4]
  assign _T_1259 = _T_1253 | _T_1258; // @[Misc.scala 214:29:freechips.rocketchip.system.DefaultRV32Config.fir@193995.4]
  assign _T_1261 = _T_1252[1] & s2_req_addr[1]; // @[Misc.scala 214:38:freechips.rocketchip.system.DefaultRV32Config.fir@193997.4]
  assign _T_1262 = _T_1253 | _T_1261; // @[Misc.scala 214:29:freechips.rocketchip.system.DefaultRV32Config.fir@193998.4]
  assign _T_1265 = ~s2_req_addr[0]; // @[Misc.scala 210:20:freechips.rocketchip.system.DefaultRV32Config.fir@194001.4]
  assign _T_1266 = _T_1256 & _T_1265; // @[Misc.scala 213:27:freechips.rocketchip.system.DefaultRV32Config.fir@194002.4]
  assign _T_1267 = _T_1252[0] & _T_1266; // @[Misc.scala 214:38:freechips.rocketchip.system.DefaultRV32Config.fir@194003.4]
  assign _T_1268 = _T_1259 | _T_1267; // @[Misc.scala 214:29:freechips.rocketchip.system.DefaultRV32Config.fir@194004.4]
  assign _T_1269 = _T_1256 & s2_req_addr[0]; // @[Misc.scala 213:27:freechips.rocketchip.system.DefaultRV32Config.fir@194005.4]
  assign _T_1270 = _T_1252[0] & _T_1269; // @[Misc.scala 214:38:freechips.rocketchip.system.DefaultRV32Config.fir@194006.4]
  assign _T_1271 = _T_1259 | _T_1270; // @[Misc.scala 214:29:freechips.rocketchip.system.DefaultRV32Config.fir@194007.4]
  assign _T_1272 = s2_req_addr[1] & _T_1265; // @[Misc.scala 213:27:freechips.rocketchip.system.DefaultRV32Config.fir@194008.4]
  assign _T_1273 = _T_1252[0] & _T_1272; // @[Misc.scala 214:38:freechips.rocketchip.system.DefaultRV32Config.fir@194009.4]
  assign _T_1274 = _T_1262 | _T_1273; // @[Misc.scala 214:29:freechips.rocketchip.system.DefaultRV32Config.fir@194010.4]
  assign _T_1275 = s2_req_addr[1] & s2_req_addr[0]; // @[Misc.scala 213:27:freechips.rocketchip.system.DefaultRV32Config.fir@194011.4]
  assign _T_1276 = _T_1252[0] & _T_1275; // @[Misc.scala 214:38:freechips.rocketchip.system.DefaultRV32Config.fir@194012.4]
  assign _T_1277 = _T_1262 | _T_1276; // @[Misc.scala 214:29:freechips.rocketchip.system.DefaultRV32Config.fir@194013.4]
  assign get_mask = {_T_1277,_T_1274,_T_1271,_T_1268}; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@194016.4]
  assign _T_2072 = 5'h4 == s2_req_cmd; // @[Mux.scala 80:60:freechips.rocketchip.system.DefaultRV32Config.fir@194913.4]
  assign _T_2073_opcode = _T_2072 ? 3'h3 : 3'h0; // @[Mux.scala 80:57:freechips.rocketchip.system.DefaultRV32Config.fir@194914.4]
  assign _T_1470_size = {{2'd0}, s2_req_size}; // @[Edges.scala 515:17:freechips.rocketchip.system.DefaultRV32Config.fir@194230.4 Edges.scala 518:15:freechips.rocketchip.system.DefaultRV32Config.fir@194234.4]
  assign _T_2073_size = _T_2072 ? _T_1470_size : 4'h0; // @[Mux.scala 80:57:freechips.rocketchip.system.DefaultRV32Config.fir@194914.4]
  assign _T_2073_source = _T_2072 & a_source; // @[Mux.scala 80:57:freechips.rocketchip.system.DefaultRV32Config.fir@194914.4]
  assign _T_2073_address = _T_2072 ? s2_req_addr : 32'h0; // @[Mux.scala 80:57:freechips.rocketchip.system.DefaultRV32Config.fir@194914.4]
  assign _T_2073_mask = _T_2072 ? get_mask : 4'h0; // @[Mux.scala 80:57:freechips.rocketchip.system.DefaultRV32Config.fir@194914.4]
  assign _T_2073_data = _T_2072 ? pstore1_data : 32'h0; // @[Mux.scala 80:57:freechips.rocketchip.system.DefaultRV32Config.fir@194914.4]
  assign _T_2074 = 5'h9 == s2_req_cmd; // @[Mux.scala 80:60:freechips.rocketchip.system.DefaultRV32Config.fir@194915.4]
  assign _T_2075_opcode = _T_2074 ? 3'h3 : _T_2073_opcode; // @[Mux.scala 80:57:freechips.rocketchip.system.DefaultRV32Config.fir@194916.4]
  assign _T_2075_param = _T_2074 ? 3'h0 : _T_2073_opcode; // @[Mux.scala 80:57:freechips.rocketchip.system.DefaultRV32Config.fir@194916.4]
  assign _T_2075_size = _T_2074 ? _T_1470_size : _T_2073_size; // @[Mux.scala 80:57:freechips.rocketchip.system.DefaultRV32Config.fir@194916.4]
  assign _T_2075_source = _T_2074 ? a_source : _T_2073_source; // @[Mux.scala 80:57:freechips.rocketchip.system.DefaultRV32Config.fir@194916.4]
  assign _T_2075_address = _T_2074 ? s2_req_addr : _T_2073_address; // @[Mux.scala 80:57:freechips.rocketchip.system.DefaultRV32Config.fir@194916.4]
  assign _T_2075_mask = _T_2074 ? get_mask : _T_2073_mask; // @[Mux.scala 80:57:freechips.rocketchip.system.DefaultRV32Config.fir@194916.4]
  assign _T_2075_data = _T_2074 ? pstore1_data : _T_2073_data; // @[Mux.scala 80:57:freechips.rocketchip.system.DefaultRV32Config.fir@194916.4]
  assign _T_2076 = 5'ha == s2_req_cmd; // @[Mux.scala 80:60:freechips.rocketchip.system.DefaultRV32Config.fir@194917.4]
  assign _T_2077_opcode = _T_2076 ? 3'h3 : _T_2075_opcode; // @[Mux.scala 80:57:freechips.rocketchip.system.DefaultRV32Config.fir@194918.4]
  assign _T_2077_param = _T_2076 ? 3'h1 : _T_2075_param; // @[Mux.scala 80:57:freechips.rocketchip.system.DefaultRV32Config.fir@194918.4]
  assign _T_2077_size = _T_2076 ? _T_1470_size : _T_2075_size; // @[Mux.scala 80:57:freechips.rocketchip.system.DefaultRV32Config.fir@194918.4]
  assign _T_2077_source = _T_2076 ? a_source : _T_2075_source; // @[Mux.scala 80:57:freechips.rocketchip.system.DefaultRV32Config.fir@194918.4]
  assign _T_2077_address = _T_2076 ? s2_req_addr : _T_2075_address; // @[Mux.scala 80:57:freechips.rocketchip.system.DefaultRV32Config.fir@194918.4]
  assign _T_2077_mask = _T_2076 ? get_mask : _T_2075_mask; // @[Mux.scala 80:57:freechips.rocketchip.system.DefaultRV32Config.fir@194918.4]
  assign _T_2077_data = _T_2076 ? pstore1_data : _T_2075_data; // @[Mux.scala 80:57:freechips.rocketchip.system.DefaultRV32Config.fir@194918.4]
  assign _T_2078 = 5'hb == s2_req_cmd; // @[Mux.scala 80:60:freechips.rocketchip.system.DefaultRV32Config.fir@194919.4]
  assign _T_2079_opcode = _T_2078 ? 3'h3 : _T_2077_opcode; // @[Mux.scala 80:57:freechips.rocketchip.system.DefaultRV32Config.fir@194920.4]
  assign _T_2079_param = _T_2078 ? 3'h2 : _T_2077_param; // @[Mux.scala 80:57:freechips.rocketchip.system.DefaultRV32Config.fir@194920.4]
  assign _T_2079_size = _T_2078 ? _T_1470_size : _T_2077_size; // @[Mux.scala 80:57:freechips.rocketchip.system.DefaultRV32Config.fir@194920.4]
  assign _T_2079_source = _T_2078 ? a_source : _T_2077_source; // @[Mux.scala 80:57:freechips.rocketchip.system.DefaultRV32Config.fir@194920.4]
  assign _T_2079_address = _T_2078 ? s2_req_addr : _T_2077_address; // @[Mux.scala 80:57:freechips.rocketchip.system.DefaultRV32Config.fir@194920.4]
  assign _T_2079_mask = _T_2078 ? get_mask : _T_2077_mask; // @[Mux.scala 80:57:freechips.rocketchip.system.DefaultRV32Config.fir@194920.4]
  assign _T_2079_data = _T_2078 ? pstore1_data : _T_2077_data; // @[Mux.scala 80:57:freechips.rocketchip.system.DefaultRV32Config.fir@194920.4]
  assign _T_2080 = 5'h8 == s2_req_cmd; // @[Mux.scala 80:60:freechips.rocketchip.system.DefaultRV32Config.fir@194921.4]
  assign _T_2081_opcode = _T_2080 ? 3'h2 : _T_2079_opcode; // @[Mux.scala 80:57:freechips.rocketchip.system.DefaultRV32Config.fir@194922.4]
  assign _T_2081_param = _T_2080 ? 3'h4 : _T_2079_param; // @[Mux.scala 80:57:freechips.rocketchip.system.DefaultRV32Config.fir@194922.4]
  assign _T_2081_size = _T_2080 ? _T_1470_size : _T_2079_size; // @[Mux.scala 80:57:freechips.rocketchip.system.DefaultRV32Config.fir@194922.4]
  assign _T_2081_source = _T_2080 ? a_source : _T_2079_source; // @[Mux.scala 80:57:freechips.rocketchip.system.DefaultRV32Config.fir@194922.4]
  assign _T_2081_address = _T_2080 ? s2_req_addr : _T_2079_address; // @[Mux.scala 80:57:freechips.rocketchip.system.DefaultRV32Config.fir@194922.4]
  assign _T_2081_mask = _T_2080 ? get_mask : _T_2079_mask; // @[Mux.scala 80:57:freechips.rocketchip.system.DefaultRV32Config.fir@194922.4]
  assign _T_2081_data = _T_2080 ? pstore1_data : _T_2079_data; // @[Mux.scala 80:57:freechips.rocketchip.system.DefaultRV32Config.fir@194922.4]
  assign _T_2082 = 5'hc == s2_req_cmd; // @[Mux.scala 80:60:freechips.rocketchip.system.DefaultRV32Config.fir@194923.4]
  assign _T_2083_opcode = _T_2082 ? 3'h2 : _T_2081_opcode; // @[Mux.scala 80:57:freechips.rocketchip.system.DefaultRV32Config.fir@194924.4]
  assign _T_2083_param = _T_2082 ? 3'h0 : _T_2081_param; // @[Mux.scala 80:57:freechips.rocketchip.system.DefaultRV32Config.fir@194924.4]
  assign _T_2083_size = _T_2082 ? _T_1470_size : _T_2081_size; // @[Mux.scala 80:57:freechips.rocketchip.system.DefaultRV32Config.fir@194924.4]
  assign _T_2083_source = _T_2082 ? a_source : _T_2081_source; // @[Mux.scala 80:57:freechips.rocketchip.system.DefaultRV32Config.fir@194924.4]
  assign _T_2083_address = _T_2082 ? s2_req_addr : _T_2081_address; // @[Mux.scala 80:57:freechips.rocketchip.system.DefaultRV32Config.fir@194924.4]
  assign _T_2083_mask = _T_2082 ? get_mask : _T_2081_mask; // @[Mux.scala 80:57:freechips.rocketchip.system.DefaultRV32Config.fir@194924.4]
  assign _T_2083_data = _T_2082 ? pstore1_data : _T_2081_data; // @[Mux.scala 80:57:freechips.rocketchip.system.DefaultRV32Config.fir@194924.4]
  assign _T_2084 = 5'hd == s2_req_cmd; // @[Mux.scala 80:60:freechips.rocketchip.system.DefaultRV32Config.fir@194925.4]
  assign _T_2085_opcode = _T_2084 ? 3'h2 : _T_2083_opcode; // @[Mux.scala 80:57:freechips.rocketchip.system.DefaultRV32Config.fir@194926.4]
  assign _T_2085_param = _T_2084 ? 3'h1 : _T_2083_param; // @[Mux.scala 80:57:freechips.rocketchip.system.DefaultRV32Config.fir@194926.4]
  assign _T_2085_size = _T_2084 ? _T_1470_size : _T_2083_size; // @[Mux.scala 80:57:freechips.rocketchip.system.DefaultRV32Config.fir@194926.4]
  assign _T_2085_source = _T_2084 ? a_source : _T_2083_source; // @[Mux.scala 80:57:freechips.rocketchip.system.DefaultRV32Config.fir@194926.4]
  assign _T_2085_address = _T_2084 ? s2_req_addr : _T_2083_address; // @[Mux.scala 80:57:freechips.rocketchip.system.DefaultRV32Config.fir@194926.4]
  assign _T_2085_mask = _T_2084 ? get_mask : _T_2083_mask; // @[Mux.scala 80:57:freechips.rocketchip.system.DefaultRV32Config.fir@194926.4]
  assign _T_2085_data = _T_2084 ? pstore1_data : _T_2083_data; // @[Mux.scala 80:57:freechips.rocketchip.system.DefaultRV32Config.fir@194926.4]
  assign _T_2086 = 5'he == s2_req_cmd; // @[Mux.scala 80:60:freechips.rocketchip.system.DefaultRV32Config.fir@194927.4]
  assign _T_2087_opcode = _T_2086 ? 3'h2 : _T_2085_opcode; // @[Mux.scala 80:57:freechips.rocketchip.system.DefaultRV32Config.fir@194928.4]
  assign _T_2087_param = _T_2086 ? 3'h2 : _T_2085_param; // @[Mux.scala 80:57:freechips.rocketchip.system.DefaultRV32Config.fir@194928.4]
  assign _T_2087_size = _T_2086 ? _T_1470_size : _T_2085_size; // @[Mux.scala 80:57:freechips.rocketchip.system.DefaultRV32Config.fir@194928.4]
  assign _T_2087_source = _T_2086 ? a_source : _T_2085_source; // @[Mux.scala 80:57:freechips.rocketchip.system.DefaultRV32Config.fir@194928.4]
  assign _T_2087_address = _T_2086 ? s2_req_addr : _T_2085_address; // @[Mux.scala 80:57:freechips.rocketchip.system.DefaultRV32Config.fir@194928.4]
  assign _T_2087_mask = _T_2086 ? get_mask : _T_2085_mask; // @[Mux.scala 80:57:freechips.rocketchip.system.DefaultRV32Config.fir@194928.4]
  assign _T_2087_data = _T_2086 ? pstore1_data : _T_2085_data; // @[Mux.scala 80:57:freechips.rocketchip.system.DefaultRV32Config.fir@194928.4]
  assign _T_2088 = 5'hf == s2_req_cmd; // @[Mux.scala 80:60:freechips.rocketchip.system.DefaultRV32Config.fir@194929.4]
  assign atomics_opcode = _T_2088 ? 3'h2 : _T_2087_opcode; // @[Mux.scala 80:57:freechips.rocketchip.system.DefaultRV32Config.fir@194930.4]
  assign atomics_param = _T_2088 ? 3'h3 : _T_2087_param; // @[Mux.scala 80:57:freechips.rocketchip.system.DefaultRV32Config.fir@194930.4]
  assign atomics_size = _T_2088 ? _T_1470_size : _T_2087_size; // @[Mux.scala 80:57:freechips.rocketchip.system.DefaultRV32Config.fir@194930.4]
  assign atomics_source = _T_2088 ? a_source : _T_2087_source; // @[Mux.scala 80:57:freechips.rocketchip.system.DefaultRV32Config.fir@194930.4]
  assign atomics_address = _T_2088 ? s2_req_addr : _T_2087_address; // @[Mux.scala 80:57:freechips.rocketchip.system.DefaultRV32Config.fir@194930.4]
  assign atomics_mask = _T_2088 ? get_mask : _T_2087_mask; // @[Mux.scala 80:57:freechips.rocketchip.system.DefaultRV32Config.fir@194930.4]
  assign atomics_data = _T_2088 ? pstore1_data : _T_2087_data; // @[Mux.scala 80:57:freechips.rocketchip.system.DefaultRV32Config.fir@194930.4]
  assign _T_2090 = ~release_ack_wait; // @[DCache.scala 551:30:freechips.rocketchip.system.DefaultRV32Config.fir@194932.4]
  assign _T_2091 = s2_valid_cached_miss & _T_2090; // @[DCache.scala 551:27:freechips.rocketchip.system.DefaultRV32Config.fir@194933.4]
  assign _T_2093 = ~s2_victim_dirty; // @[DCache.scala 551:117:freechips.rocketchip.system.DefaultRV32Config.fir@194935.4]
  assign _T_2095 = _T_2091 & _T_2093; // @[DCache.scala 551:48:freechips.rocketchip.system.DefaultRV32Config.fir@194937.4]
  assign tl_out_a_valid = s2_valid_uncached_pending | _T_2095; // @[DCache.scala 550:67:freechips.rocketchip.system.DefaultRV32Config.fir@194938.4]
  assign _T_2154 = ~s2_write; // @[DCache.scala 553:9:freechips.rocketchip.system.DefaultRV32Config.fir@195006.4]
  assign _T_2156 = ~s2_read; // @[DCache.scala 555:9:freechips.rocketchip.system.DefaultRV32Config.fir@195008.4]
  assign _T_2157_opcode = _T_2156 ? 3'h0 : atomics_opcode; // @[DCache.scala 555:8:freechips.rocketchip.system.DefaultRV32Config.fir@195009.4]
  assign _T_2157_param = _T_2156 ? 3'h0 : atomics_param; // @[DCache.scala 555:8:freechips.rocketchip.system.DefaultRV32Config.fir@195009.4]
  assign _T_2157_size = _T_2156 ? _T_1470_size : atomics_size; // @[DCache.scala 555:8:freechips.rocketchip.system.DefaultRV32Config.fir@195009.4]
  assign _T_2157_source = _T_2156 ? a_source : atomics_source; // @[DCache.scala 555:8:freechips.rocketchip.system.DefaultRV32Config.fir@195009.4]
  assign _T_2157_address = _T_2156 ? s2_req_addr : atomics_address; // @[DCache.scala 555:8:freechips.rocketchip.system.DefaultRV32Config.fir@195009.4]
  assign _T_2157_mask = _T_2156 ? get_mask : atomics_mask; // @[DCache.scala 555:8:freechips.rocketchip.system.DefaultRV32Config.fir@195009.4]
  assign _T_2157_data = _T_2156 ? pstore1_data : atomics_data; // @[DCache.scala 555:8:freechips.rocketchip.system.DefaultRV32Config.fir@195009.4]
  assign _T_2158_opcode = _T_403 ? 3'h1 : _T_2157_opcode; // @[DCache.scala 554:8:freechips.rocketchip.system.DefaultRV32Config.fir@195010.4]
  assign _T_2158_param = _T_403 ? 3'h0 : _T_2157_param; // @[DCache.scala 554:8:freechips.rocketchip.system.DefaultRV32Config.fir@195010.4]
  assign _T_2158_size = _T_403 ? _T_1470_size : _T_2157_size; // @[DCache.scala 554:8:freechips.rocketchip.system.DefaultRV32Config.fir@195010.4]
  assign _T_2158_source = _T_403 ? a_source : _T_2157_source; // @[DCache.scala 554:8:freechips.rocketchip.system.DefaultRV32Config.fir@195010.4]
  assign _T_2158_address = _T_403 ? s2_req_addr : _T_2157_address; // @[DCache.scala 554:8:freechips.rocketchip.system.DefaultRV32Config.fir@195010.4]
  assign putpartial_mask = a_mask[3:0]; // @[Edges.scala 485:17:freechips.rocketchip.system.DefaultRV32Config.fir@194181.4 Edges.scala 491:15:freechips.rocketchip.system.DefaultRV32Config.fir@194188.4]
  assign _T_2158_mask = _T_403 ? putpartial_mask : _T_2157_mask; // @[DCache.scala 554:8:freechips.rocketchip.system.DefaultRV32Config.fir@195010.4]
  assign _T_2158_data = _T_403 ? pstore1_data : _T_2157_data; // @[DCache.scala 554:8:freechips.rocketchip.system.DefaultRV32Config.fir@195010.4]
  assign _T_2159_opcode = _T_2154 ? 3'h4 : _T_2158_opcode; // @[DCache.scala 553:8:freechips.rocketchip.system.DefaultRV32Config.fir@195011.4]
  assign _T_2159_param = _T_2154 ? 3'h0 : _T_2158_param; // @[DCache.scala 553:8:freechips.rocketchip.system.DefaultRV32Config.fir@195011.4]
  assign _T_2159_size = _T_2154 ? _T_1470_size : _T_2158_size; // @[DCache.scala 553:8:freechips.rocketchip.system.DefaultRV32Config.fir@195011.4]
  assign _T_2159_source = _T_2154 ? a_source : _T_2158_source; // @[DCache.scala 553:8:freechips.rocketchip.system.DefaultRV32Config.fir@195011.4]
  assign _T_2159_address = _T_2154 ? s2_req_addr : _T_2158_address; // @[DCache.scala 553:8:freechips.rocketchip.system.DefaultRV32Config.fir@195011.4]
  assign _T_2159_mask = _T_2154 ? get_mask : _T_2158_mask; // @[DCache.scala 553:8:freechips.rocketchip.system.DefaultRV32Config.fir@195011.4]
  assign _T_2159_data = _T_2154 ? 32'h0 : _T_2158_data; // @[DCache.scala 553:8:freechips.rocketchip.system.DefaultRV32Config.fir@195011.4]
  assign _T_2120_param = {{1'd0}, s2_grow_param}; // @[Edges.scala 347:17:freechips.rocketchip.system.DefaultRV32Config.fir@194963.4 Edges.scala 349:15:freechips.rocketchip.system.DefaultRV32Config.fir@194966.4]
  assign _T_2162 = 2'h1 << a_source; // @[OneHot.scala 65:12:freechips.rocketchip.system.DefaultRV32Config.fir@195015.4]
  assign a_sel = _T_2162[1]; // @[DCache.scala 574:66:freechips.rocketchip.system.DefaultRV32Config.fir@195017.4]
  assign _T_2164 = auto_out_a_ready & tl_out_a_valid; // @[Decoupled.scala 40:37:freechips.rocketchip.system.DefaultRV32Config.fir@195018.4]
  assign _GEN_139 = a_sel | uncachedInFlight_0; // @[DCache.scala 578:18:freechips.rocketchip.system.DefaultRV32Config.fir@195022.8]
  assign _T_2171 = 27'hfff << auto_out_d_bits_size; // @[package.scala 207:77:freechips.rocketchip.system.DefaultRV32Config.fir@195037.4]
  assign _T_2173 = ~_T_2171[11:0]; // @[package.scala 207:46:freechips.rocketchip.system.DefaultRV32Config.fir@195039.4]
  assign _T_2176 = auto_out_d_bits_opcode[0] ? _T_2173[11:2] : 10'h0; // @[Edges.scala 222:14:freechips.rocketchip.system.DefaultRV32Config.fir@195042.4]
  assign _T_2179 = _T_2177 - 10'h1; // @[Edges.scala 231:28:freechips.rocketchip.system.DefaultRV32Config.fir@195045.4]
  assign _T_2180 = _T_2177 == 10'h1; // @[Edges.scala 233:25:freechips.rocketchip.system.DefaultRV32Config.fir@195047.4]
  assign _T_2181 = _T_2176 == 10'h0; // @[Edges.scala 233:47:freechips.rocketchip.system.DefaultRV32Config.fir@195048.4]
  assign d_last = _T_2180 | _T_2181; // @[Edges.scala 233:37:freechips.rocketchip.system.DefaultRV32Config.fir@195049.4]
  assign d_done = d_last & _T_2217; // @[Edges.scala 234:22:freechips.rocketchip.system.DefaultRV32Config.fir@195050.4]
  assign _T_2182 = ~_T_2179; // @[Edges.scala 235:27:freechips.rocketchip.system.DefaultRV32Config.fir@195051.4]
  assign _T_2183 = _T_2176 & _T_2182; // @[Edges.scala 235:25:freechips.rocketchip.system.DefaultRV32Config.fir@195052.4]
  assign d_address_inc = {_T_2183, 2'h0}; // @[Edges.scala 270:29:freechips.rocketchip.system.DefaultRV32Config.fir@195057.4]
  assign _T_2192 = ~grantIsUncached; // @[DCache.scala 606:129:freechips.rocketchip.system.DefaultRV32Config.fir@195067.4]
  assign grantIsVoluntary = auto_out_d_bits_opcode == 3'h6; // @[DCache.scala 608:32:freechips.rocketchip.system.DefaultRV32Config.fir@195080.4]
  assign _T_2205 = blockProbeAfterGrantCount - 3'h1; // @[DCache.scala 612:97:freechips.rocketchip.system.DefaultRV32Config.fir@195087.6]
  assign _T_2214 = 2'h1 << auto_out_d_bits_source; // @[OneHot.scala 65:12:freechips.rocketchip.system.DefaultRV32Config.fir@195100.4]
  assign uncachedRespIdxOH = _T_2214[1]; // @[DCache.scala 615:90:freechips.rocketchip.system.DefaultRV32Config.fir@195102.4]
  assign _T_2219 = cached_grant_wait | reset; // @[DCache.scala 620:13:freechips.rocketchip.system.DefaultRV32Config.fir@195110.8]
  assign _T_2220 = ~_T_2219; // @[DCache.scala 620:13:freechips.rocketchip.system.DefaultRV32Config.fir@195111.8]
  assign _T_2222 = uncachedRespIdxOH & d_last; // @[DCache.scala 629:17:freechips.rocketchip.system.DefaultRV32Config.fir@195126.10]
  assign _T_2224 = uncachedInFlight_0 | reset; // @[DCache.scala 630:17:freechips.rocketchip.system.DefaultRV32Config.fir@195129.12]
  assign _T_2225 = ~_T_2224; // @[DCache.scala 630:17:freechips.rocketchip.system.DefaultRV32Config.fir@195130.12]
  assign dontCareBits = {s1_paddr[31:2], 2'h0}; // @[DCache.scala 644:55:freechips.rocketchip.system.DefaultRV32Config.fir@195145.12]
  assign _GEN_376 = {{30'd0}, uncachedReqs_0_addr[1:0]}; // @[DCache.scala 645:26:freechips.rocketchip.system.DefaultRV32Config.fir@195147.12]
  assign _T_2229 = dontCareBits | _GEN_376; // @[DCache.scala 645:26:freechips.rocketchip.system.DefaultRV32Config.fir@195147.12]
  assign _T_2231 = release_ack_wait | reset; // @[DCache.scala 651:13:freechips.rocketchip.system.DefaultRV32Config.fir@195155.12]
  assign _T_2232 = ~_T_2231; // @[DCache.scala 651:13:freechips.rocketchip.system.DefaultRV32Config.fir@195156.12]
  assign _GEN_191 = grantIsVoluntary ? 1'h0 : release_ack_wait; // @[DCache.scala 650:36:freechips.rocketchip.system.DefaultRV32Config.fir@195153.10]
  assign _GEN_200 = grantIsUncached ? release_ack_wait : _GEN_191; // @[DCache.scala 627:35:freechips.rocketchip.system.DefaultRV32Config.fir@195124.8]
  assign _GEN_204 = grantIsCached & d_last; // @[DCache.scala 618:26:freechips.rocketchip.system.DefaultRV32Config.fir@195107.6]
  assign _GEN_213 = grantIsCached ? release_ack_wait : _GEN_200; // @[DCache.scala 618:26:freechips.rocketchip.system.DefaultRV32Config.fir@195107.6]
  assign _GEN_226 = _T_2217 ? _GEN_213 : release_ack_wait; // @[DCache.scala 617:26:freechips.rocketchip.system.DefaultRV32Config.fir@195106.4]
  assign _T_2233 = auto_out_d_valid & d_first; // @[DCache.scala 657:36:freechips.rocketchip.system.DefaultRV32Config.fir@195164.4]
  assign _T_2234 = _T_2233 & grantIsCached; // @[DCache.scala 657:47:freechips.rocketchip.system.DefaultRV32Config.fir@195165.4]
  assign _T_2235 = _T_2234 & canAcceptCachedGrant; // @[DCache.scala 657:64:freechips.rocketchip.system.DefaultRV32Config.fir@195166.4]
  assign tl_out__e_valid = _T_2248 ? 1'h0 : _T_2235; // @[DCache.scala 665:51:freechips.rocketchip.system.DefaultRV32Config.fir@195189.4]
  assign _T_2237 = auto_out_e_ready & tl_out__e_valid; // @[Decoupled.scala 40:37:freechips.rocketchip.system.DefaultRV32Config.fir@195172.4]
  assign _T_2239 = _T_2217 & d_first; // @[DCache.scala 659:47:freechips.rocketchip.system.DefaultRV32Config.fir@195174.4]
  assign _T_2240 = _T_2239 & grantIsCached; // @[DCache.scala 659:58:freechips.rocketchip.system.DefaultRV32Config.fir@195175.4]
  assign _T_2241 = _T_2237 == _T_2240; // @[DCache.scala 659:26:freechips.rocketchip.system.DefaultRV32Config.fir@195176.4]
  assign _T_2243 = _T_2241 | reset; // @[DCache.scala 659:9:freechips.rocketchip.system.DefaultRV32Config.fir@195178.4]
  assign _T_2244 = ~_T_2243; // @[DCache.scala 659:9:freechips.rocketchip.system.DefaultRV32Config.fir@195179.4]
  assign _T_2245 = auto_out_d_valid & grantIsRefill; // @[DCache.scala 664:44:freechips.rocketchip.system.DefaultRV32Config.fir@195184.4]
  assign _T_2246 = _T_2245 & canAcceptCachedGrant; // @[DCache.scala 664:61:freechips.rocketchip.system.DefaultRV32Config.fir@195185.4]
  assign _T_2250 = {s2_vaddr[31:6], 6'h0}; // @[DCache.scala 671:57:freechips.rocketchip.system.DefaultRV32Config.fir@195195.4]
  assign _GEN_377 = {{20'd0}, d_address_inc}; // @[DCache.scala 671:67:freechips.rocketchip.system.DefaultRV32Config.fir@195196.4]
  assign _T_2251 = _T_2250 | _GEN_377; // @[DCache.scala 671:67:freechips.rocketchip.system.DefaultRV32Config.fir@195196.4]
  assign _T_2254 = grantIsCached & d_done; // @[DCache.scala 684:43:freechips.rocketchip.system.DefaultRV32Config.fir@195204.4]
  assign _T_2255 = ~auto_out_d_bits_denied; // @[DCache.scala 684:56:freechips.rocketchip.system.DefaultRV32Config.fir@195205.4]
  assign _T_2313 = {s2_write,_T_526,auto_out_d_bits_param}; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@195268.4]
  assign _T_2322 = 4'h1 == _T_2313; // @[Mux.scala 80:60:freechips.rocketchip.system.DefaultRV32Config.fir@195277.4]
  assign _T_2323 = _T_2322 ? 2'h1 : 2'h0; // @[Mux.scala 80:57:freechips.rocketchip.system.DefaultRV32Config.fir@195278.4]
  assign _T_2324 = 4'h0 == _T_2313; // @[Mux.scala 80:60:freechips.rocketchip.system.DefaultRV32Config.fir@195279.4]
  assign _T_2325 = _T_2324 ? 2'h2 : _T_2323; // @[Mux.scala 80:57:freechips.rocketchip.system.DefaultRV32Config.fir@195280.4]
  assign _T_2326 = 4'h4 == _T_2313; // @[Mux.scala 80:60:freechips.rocketchip.system.DefaultRV32Config.fir@195281.4]
  assign _T_2327 = _T_2326 ? 2'h2 : _T_2325; // @[Mux.scala 80:57:freechips.rocketchip.system.DefaultRV32Config.fir@195282.4]
  assign _T_2328 = 4'hc == _T_2313; // @[Mux.scala 80:60:freechips.rocketchip.system.DefaultRV32Config.fir@195283.4]
  assign _T_2329 = _T_2328 ? 2'h3 : _T_2327; // @[Mux.scala 80:57:freechips.rocketchip.system.DefaultRV32Config.fir@195284.4]
  assign _GEN_229 = auto_out_d_valid ? 1'h0 : _GEN_31; // @[DCache.scala 698:29:freechips.rocketchip.system.DefaultRV32Config.fir@195300.6]
  assign _GEN_230 = auto_out_d_valid | _T_2246; // @[DCache.scala 698:29:freechips.rocketchip.system.DefaultRV32Config.fir@195300.6]
  assign _GEN_231 = auto_out_d_valid ? 1'h0 : 1'h1; // @[DCache.scala 698:29:freechips.rocketchip.system.DefaultRV32Config.fir@195300.6]
  assign _T_2343 = ~block_probe_for_core_progress; // @[DCache.scala 712:48:freechips.rocketchip.system.DefaultRV32Config.fir@195318.4]
  assign _T_2344 = _T_2343 | lrscBackingOff; // @[DCache.scala 712:79:freechips.rocketchip.system.DefaultRV32Config.fir@195319.4]
  assign _T_2345 = auto_out_b_valid & _T_2344; // @[DCache.scala 712:44:freechips.rocketchip.system.DefaultRV32Config.fir@195320.4]
  assign _T_2353 = {1'h0,auto_out_b_bits_address}; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@195332.4]
  assign _T_2364 = _T_2362 - 10'h1; // @[Edges.scala 231:28:freechips.rocketchip.system.DefaultRV32Config.fir@195346.4]
  assign _T_2367 = ~_T_2364; // @[Edges.scala 235:27:freechips.rocketchip.system.DefaultRV32Config.fir@195352.4]
  assign c_count = _T_2361 & _T_2367; // @[Edges.scala 235:25:freechips.rocketchip.system.DefaultRV32Config.fir@195353.4]
  assign _T_2373 = ~_T_2354; // @[DCache.scala 725:47:freechips.rocketchip.system.DefaultRV32Config.fir@195368.4]
  assign releaseRejected = s2_release_data_valid & _T_2373; // @[DCache.scala 725:44:freechips.rocketchip.system.DefaultRV32Config.fir@195369.4]
  assign _T_2370 = ~releaseRejected; // @[DCache.scala 724:67:freechips.rocketchip.system.DefaultRV32Config.fir@195363.4]
  assign _T_2375 = {1'h0,c_count}; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@195371.4]
  assign _T_2376 = {1'h0,s2_release_data_valid}; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@195372.4]
  assign _GEN_378 = {{1'd0}, s1_release_data_valid}; // @[DCache.scala 726:101:freechips.rocketchip.system.DefaultRV32Config.fir@195373.4]
  assign _T_2378 = _GEN_378 + _T_2376; // @[DCache.scala 726:101:freechips.rocketchip.system.DefaultRV32Config.fir@195374.4]
  assign _T_2379 = releaseRejected ? 2'h0 : _T_2378; // @[DCache.scala 726:52:freechips.rocketchip.system.DefaultRV32Config.fir@195375.4]
  assign _GEN_379 = {{9'd0}, _T_2379}; // @[DCache.scala 726:47:freechips.rocketchip.system.DefaultRV32Config.fir@195376.4]
  assign releaseDataBeat = _T_2375 + _GEN_379; // @[DCache.scala 726:47:freechips.rocketchip.system.DefaultRV32Config.fir@195377.4]
  assign _T_2385 = s2_valid_flush_line | io_cpu_s2_nack; // @[DCache.scala 739:52:freechips.rocketchip.system.DefaultRV32Config.fir@195416.6]
  assign _T_2387 = _T_2385 | reset; // @[DCache.scala 739:13:freechips.rocketchip.system.DefaultRV32Config.fir@195418.6]
  assign _T_2388 = ~_T_2387; // @[DCache.scala 739:13:freechips.rocketchip.system.DefaultRV32Config.fir@195419.6]
  assign discard_line = s2_valid_flush_line & s2_req_size[1]; // @[DCache.scala 740:46:freechips.rocketchip.system.DefaultRV32Config.fir@195425.6]
  assign _T_2393 = ~discard_line; // @[DCache.scala 741:47:freechips.rocketchip.system.DefaultRV32Config.fir@195429.6]
  assign _T_2394 = s2_victim_dirty & _T_2393; // @[DCache.scala 741:44:freechips.rocketchip.system.DefaultRV32Config.fir@195430.6]
  assign _T_2395 = _T_2394 ? 3'h1 : 3'h6; // @[DCache.scala 741:27:freechips.rocketchip.system.DefaultRV32Config.fir@195431.6]
  assign _T_2397 = {s2_victim_tag,s2_req_addr[11:6]}; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@195434.6]
  assign res_2_address = {_T_2397, 6'h0}; // @[DCache.scala 742:96:freechips.rocketchip.system.DefaultRV32Config.fir@195435.6]
  assign _GEN_239 = s2_want_victimize ? _T_2395 : release_state; // @[DCache.scala 738:25:freechips.rocketchip.system.DefaultRV32Config.fir@195414.4]
  assign _T_2400 = releaseDone ? 3'h7 : 3'h3; // @[DCache.scala 753:29:freechips.rocketchip.system.DefaultRV32Config.fir@195458.12]
  assign _T_2402 = releaseDone ? 3'h0 : 3'h5; // @[DCache.scala 757:29:freechips.rocketchip.system.DefaultRV32Config.fir@195465.12]
  assign _GEN_250 = _T_2399 ? s2_report_param : 3'h5; // @[DCache.scala 750:45:freechips.rocketchip.system.DefaultRV32Config.fir@195455.10]
  assign _GEN_256 = _T_2399 ? _T_2400 : _T_2402; // @[DCache.scala 750:45:freechips.rocketchip.system.DefaultRV32Config.fir@195455.10]
  assign _GEN_258 = s2_prb_ack_data ? 3'h2 : _GEN_256; // @[DCache.scala 748:36:freechips.rocketchip.system.DefaultRV32Config.fir@195450.8]
  assign _GEN_261 = s2_prb_ack_data ? 3'h5 : _GEN_250; // @[DCache.scala 748:36:freechips.rocketchip.system.DefaultRV32Config.fir@195450.8]
  assign _GEN_268 = pma_checker__T_2026 ? 3'h4 : _GEN_258; // @[DCache.scala 746:28:freechips.rocketchip.system.DefaultRV32Config.fir@195446.6]
  assign _GEN_271 = pma_checker__T_2026 ? 3'h5 : _GEN_261; // @[DCache.scala 746:28:freechips.rocketchip.system.DefaultRV32Config.fir@195446.6]
  assign _GEN_279 = s2_probe ? _GEN_268 : _GEN_239; // @[DCache.scala 744:21:freechips.rocketchip.system.DefaultRV32Config.fir@195442.4]
  assign _GEN_282 = s2_probe ? _GEN_271 : 3'h5; // @[DCache.scala 744:21:freechips.rocketchip.system.DefaultRV32Config.fir@195442.4]
  assign _T_2403 = release_state == 3'h4; // @[DCache.scala 761:25:freechips.rocketchip.system.DefaultRV32Config.fir@195472.4]
  assign _T_2406 = {1'h0,probe_bits_address}; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@195478.6]
  assign _GEN_289 = metaArb_io_in_6_ready ? 3'h0 : _GEN_279; // @[DCache.scala 765:37:freechips.rocketchip.system.DefaultRV32Config.fir@195480.6]
  assign _GEN_290 = metaArb_io_in_6_ready | _T_17; // @[DCache.scala 765:37:freechips.rocketchip.system.DefaultRV32Config.fir@195480.6]
  assign _GEN_293 = _T_2403 ? _T_2406 : _T_2353; // @[DCache.scala 761:44:freechips.rocketchip.system.DefaultRV32Config.fir@195473.4]
  assign _GEN_294 = _T_2403 ? _GEN_289 : _GEN_279; // @[DCache.scala 761:44:freechips.rocketchip.system.DefaultRV32Config.fir@195473.4]
  assign _GEN_296 = releaseDone ? 3'h0 : _GEN_294; // @[DCache.scala 772:26:freechips.rocketchip.system.DefaultRV32Config.fir@195488.6]
  assign _GEN_298 = _T_2407 ? _GEN_296 : _GEN_294; // @[DCache.scala 770:47:freechips.rocketchip.system.DefaultRV32Config.fir@195486.4]
  assign _GEN_302 = _T_2408 ? s2_report_param : _GEN_282; // @[DCache.scala 774:48:freechips.rocketchip.system.DefaultRV32Config.fir@195493.4]
  assign _GEN_311 = _T_2409 ? s2_report_param : _GEN_302; // @[DCache.scala 779:48:freechips.rocketchip.system.DefaultRV32Config.fir@195501.4]
  assign _T_2434 = _T_2354 & c_first; // @[DCache.scala 792:29:freechips.rocketchip.system.DefaultRV32Config.fir@195546.6]
  assign _GEN_319 = _T_2434 | _GEN_226; // @[DCache.scala 792:41:freechips.rocketchip.system.DefaultRV32Config.fir@195547.6]
  assign newCoh_state = _T_2412 ? voluntaryNewCoh_state : probeNewCoh_state; // @[DCache.scala 783:81:freechips.rocketchip.system.DefaultRV32Config.fir@195510.4]
  assign _T_2436 = releaseDataBeat < 11'h10; // @[DCache.scala 803:60:freechips.rocketchip.system.DefaultRV32Config.fir@195557.4]
  assign _T_2439 = {probe_bits_address[11:6], 6'h0}; // @[DCache.scala 806:55:freechips.rocketchip.system.DefaultRV32Config.fir@195563.4]
  assign _T_2441 = {releaseDataBeat[3:0], 2'h0}; // @[DCache.scala 806:117:freechips.rocketchip.system.DefaultRV32Config.fir@195565.4]
  assign _GEN_381 = {{6'd0}, _T_2441}; // @[DCache.scala 806:72:freechips.rocketchip.system.DefaultRV32Config.fir@195566.4]
  assign _T_2446 = release_state == 3'h7; // @[package.scala 15:47:freechips.rocketchip.system.DefaultRV32Config.fir@195573.4]
  assign _T_2455 = metaArb_io_in_4_ready & metaArb_io_in_4_valid; // @[Decoupled.scala 40:37:freechips.rocketchip.system.DefaultRV32Config.fir@195591.4]
  assign _T_2462 = s1_valid | s2_valid; // @[DCache.scala 829:57:freechips.rocketchip.system.DefaultRV32Config.fir@195606.4]
  assign _T_2463 = _T_2462 | cached_grant_wait; // @[DCache.scala 829:94:freechips.rocketchip.system.DefaultRV32Config.fir@195607.4]
  assign _T_2465 = _T_2463 | _T_621; // @[DCache.scala 829:115:freechips.rocketchip.system.DefaultRV32Config.fir@195609.4]
  assign _T_2483 = _T_781 | reset; // @[DCache.scala 851:11:freechips.rocketchip.system.DefaultRV32Config.fir@195656.6]
  assign _T_2484 = ~_T_2483; // @[DCache.scala 851:11:freechips.rocketchip.system.DefaultRV32Config.fir@195657.6]
  assign _T_2491 = s2_req_addr[1] ? s2_data_corrected[31:16] : s2_data_corrected[15:0]; // @[AMOALU.scala 39:24:freechips.rocketchip.system.DefaultRV32Config.fir@195674.4]
  assign _T_2494 = s2_req_size == 2'h1; // @[AMOALU.scala 42:26:freechips.rocketchip.system.DefaultRV32Config.fir@195677.4]
  assign _T_2497 = s2_req_signed & _T_2491[15]; // @[AMOALU.scala 42:76:freechips.rocketchip.system.DefaultRV32Config.fir@195680.4]
  assign _T_2499 = _T_2497 ? 16'hffff : 16'h0; // @[Bitwise.scala 72:12:freechips.rocketchip.system.DefaultRV32Config.fir@195682.4]
  assign _T_2501 = _T_2494 ? _T_2499 : s2_data_corrected[31:16]; // @[AMOALU.scala 42:20:freechips.rocketchip.system.DefaultRV32Config.fir@195684.4]
  assign _T_2502 = {_T_2501,_T_2491}; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@195685.4]
  assign _T_2506 = s2_req_addr[0] ? _T_2502[15:8] : _T_2502[7:0]; // @[AMOALU.scala 39:24:freechips.rocketchip.system.DefaultRV32Config.fir@195689.4]
  assign _T_2508 = _T_405 ? 8'h0 : _T_2506; // @[AMOALU.scala 41:23:freechips.rocketchip.system.DefaultRV32Config.fir@195691.4]
  assign _T_2509 = s2_req_size == 2'h0; // @[AMOALU.scala 42:26:freechips.rocketchip.system.DefaultRV32Config.fir@195692.4]
  assign _T_2510 = _T_2509 | _T_405; // @[AMOALU.scala 42:38:freechips.rocketchip.system.DefaultRV32Config.fir@195693.4]
  assign _T_2512 = s2_req_signed & _T_2508[7]; // @[AMOALU.scala 42:76:freechips.rocketchip.system.DefaultRV32Config.fir@195695.4]
  assign _T_2514 = _T_2512 ? 24'hffffff : 24'h0; // @[Bitwise.scala 72:12:freechips.rocketchip.system.DefaultRV32Config.fir@195697.4]
  assign _T_2516 = _T_2510 ? _T_2514 : _T_2502[31:8]; // @[AMOALU.scala 42:20:freechips.rocketchip.system.DefaultRV32Config.fir@195699.4]
  assign _T_2517 = {_T_2516,_T_2508}; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@195700.4]
  assign _GEN_382 = {{31'd0}, s2_sc_fail}; // @[DCache.scala 873:41:freechips.rocketchip.system.DefaultRV32Config.fir@195701.4]
  assign _GEN_337 = _T_2523 | resetting; // @[DCache.scala 908:27:freechips.rocketchip.system.DefaultRV32Config.fir@195722.4]
  assign flushCounterNext = flushCounter + 8'h1; // @[DCache.scala 910:39:freechips.rocketchip.system.DefaultRV32Config.fir@195726.4]
  assign flushDone = flushCounterNext[8:6] == 3'h4; // @[DCache.scala 911:57:freechips.rocketchip.system.DefaultRV32Config.fir@195728.4]
  assign _T_2542 = {metaArb_io_in_5_bits_idx, 6'h0}; // @[DCache.scala 919:98:freechips.rocketchip.system.DefaultRV32Config.fir@195751.4]
  assign _GEN_339 = resetting ? flushCounterNext : {{1'd0}, flushCounter}; // @[DCache.scala 952:20:freechips.rocketchip.system.DefaultRV32Config.fir@195771.4]
  assign _T_2606 = _T_2604 - 10'h1; // @[Edges.scala 231:28:freechips.rocketchip.system.DefaultRV32Config.fir@195839.4]
  assign _T_2607 = _T_2604 == 10'h0; // @[Edges.scala 232:25:freechips.rocketchip.system.DefaultRV32Config.fir@195840.4]
  assign _T_2608 = _T_2604 == 10'h1; // @[Edges.scala 233:25:freechips.rocketchip.system.DefaultRV32Config.fir@195841.4]
  assign _T_2610 = _T_2608 | _T_2366; // @[Edges.scala 233:37:freechips.rocketchip.system.DefaultRV32Config.fir@195843.4]
  assign _T_2725 = ~grantIsCached; // @[DCache.scala 1028:35:freechips.rocketchip.system.DefaultRV32Config.fir@195977.4]
  assign auto_out_a_valid = s2_valid_uncached_pending | _T_2095; // @[LazyModule.scala 305:12:freechips.rocketchip.system.DefaultRV32Config.fir@192106.4]
  assign auto_out_a_bits_opcode = _T_619 ? 3'h6 : _T_2159_opcode; // @[LazyModule.scala 305:12:freechips.rocketchip.system.DefaultRV32Config.fir@192106.4]
  assign auto_out_a_bits_param = _T_619 ? _T_2120_param : _T_2159_param; // @[LazyModule.scala 305:12:freechips.rocketchip.system.DefaultRV32Config.fir@192106.4]
  assign auto_out_a_bits_size = _T_619 ? 4'h6 : _T_2159_size; // @[LazyModule.scala 305:12:freechips.rocketchip.system.DefaultRV32Config.fir@192106.4]
  assign auto_out_a_bits_source = _T_619 ? 1'h0 : _T_2159_source; // @[LazyModule.scala 305:12:freechips.rocketchip.system.DefaultRV32Config.fir@192106.4]
  assign auto_out_a_bits_address = _T_619 ? acquire_address : _T_2159_address; // @[LazyModule.scala 305:12:freechips.rocketchip.system.DefaultRV32Config.fir@192106.4]
  assign auto_out_a_bits_mask = _T_619 ? 4'hf : _T_2159_mask; // @[LazyModule.scala 305:12:freechips.rocketchip.system.DefaultRV32Config.fir@192106.4]
  assign auto_out_a_bits_data = _T_619 ? 32'h0 : _T_2159_data; // @[LazyModule.scala 305:12:freechips.rocketchip.system.DefaultRV32Config.fir@192106.4]
  assign auto_out_b_ready = metaArb_io_in_6_ready & _T_2349; // @[LazyModule.scala 305:12:freechips.rocketchip.system.DefaultRV32Config.fir@192106.4]
  assign auto_out_c_valid = _T_2408 | _GEN_297; // @[LazyModule.scala 305:12:freechips.rocketchip.system.DefaultRV32Config.fir@192106.4]
  assign auto_out_c_bits_opcode = _T_2412 ? 3'h7 : _GEN_310; // @[LazyModule.scala 305:12:freechips.rocketchip.system.DefaultRV32Config.fir@192106.4]
  assign auto_out_c_bits_param = _T_2412 ? s2_shrink_param : _GEN_311; // @[LazyModule.scala 305:12:freechips.rocketchip.system.DefaultRV32Config.fir@192106.4]
  assign auto_out_c_bits_size = _T_2412 ? 4'h6 : probe_bits_size; // @[LazyModule.scala 305:12:freechips.rocketchip.system.DefaultRV32Config.fir@192106.4]
  assign auto_out_c_bits_source = probe_bits_source; // @[LazyModule.scala 305:12:freechips.rocketchip.system.DefaultRV32Config.fir@192106.4]
  assign auto_out_c_bits_address = probe_bits_address; // @[LazyModule.scala 305:12:freechips.rocketchip.system.DefaultRV32Config.fir@192106.4]
  assign auto_out_c_bits_data = {_T_600,_T_599}; // @[LazyModule.scala 305:12:freechips.rocketchip.system.DefaultRV32Config.fir@192106.4]
  assign auto_out_d_ready = _T_2334 ? 1'h0 : _GEN_228; // @[LazyModule.scala 305:12:freechips.rocketchip.system.DefaultRV32Config.fir@192106.4]
  assign auto_out_e_valid = _T_2248 ? 1'h0 : _T_2235; // @[LazyModule.scala 305:12:freechips.rocketchip.system.DefaultRV32Config.fir@192106.4]
  assign auto_out_e_bits_sink = auto_out_d_bits_sink; // @[LazyModule.scala 305:12:freechips.rocketchip.system.DefaultRV32Config.fir@192106.4]
  assign io_cpu_req_ready = _T_2334 ? _GEN_229 : _GEN_31; // @[DCache.scala 203:20:freechips.rocketchip.system.DefaultRV32Config.fir@192337.4 DCache.scala 218:64:freechips.rocketchip.system.DefaultRV32Config.fir@192447.6 DCache.scala 226:53:freechips.rocketchip.system.DefaultRV32Config.fir@192515.6 DCache.scala 234:98:freechips.rocketchip.system.DefaultRV32Config.fir@192536.6 DCache.scala 699:26:freechips.rocketchip.system.DefaultRV32Config.fir@195301.8]
  assign io_cpu_s2_nack = _T_780 & _T_781; // @[DCache.scala 396:18:freechips.rocketchip.system.DefaultRV32Config.fir@193362.4]
  assign io_cpu_resp_valid = s2_valid_hit_pre_data_ecc_and_waw | doUncachedResp; // @[DCache.scala 848:21:freechips.rocketchip.system.DefaultRV32Config.fir@195648.4]
  assign io_cpu_resp_bits_addr = doUncachedResp ? s2_uncached_resp_addr : s2_req_addr; // @[DCache.scala 819:20:freechips.rocketchip.system.DefaultRV32Config.fir@195595.4 DCache.scala 853:27:freechips.rocketchip.system.DefaultRV32Config.fir@195663.6]
  assign io_cpu_resp_bits_tag = s2_req_tag; // @[DCache.scala 819:20:freechips.rocketchip.system.DefaultRV32Config.fir@195595.4]
  assign io_cpu_resp_bits_cmd = s2_req_cmd; // @[DCache.scala 819:20:freechips.rocketchip.system.DefaultRV32Config.fir@195595.4]
  assign io_cpu_resp_bits_size = s2_req_size; // @[DCache.scala 819:20:freechips.rocketchip.system.DefaultRV32Config.fir@195595.4]
  assign io_cpu_resp_bits_signed = s2_req_signed; // @[DCache.scala 819:20:freechips.rocketchip.system.DefaultRV32Config.fir@195595.4]
  assign io_cpu_resp_bits_dprv = s2_req_dprv; // @[DCache.scala 819:20:freechips.rocketchip.system.DefaultRV32Config.fir@195595.4]
  assign io_cpu_resp_bits_data = _T_2517 | _GEN_382; // @[DCache.scala 819:20:freechips.rocketchip.system.DefaultRV32Config.fir@195595.4 DCache.scala 873:25:freechips.rocketchip.system.DefaultRV32Config.fir@195702.4]
  assign io_cpu_resp_bits_mask = 4'h0; // @[DCache.scala 819:20:freechips.rocketchip.system.DefaultRV32Config.fir@195595.4]
  assign io_cpu_resp_bits_replay = doUncachedResp; // @[DCache.scala 821:27:freechips.rocketchip.system.DefaultRV32Config.fir@195597.4 DCache.scala 852:29:freechips.rocketchip.system.DefaultRV32Config.fir@195662.6]
  assign io_cpu_resp_bits_has_data = _T_384 | _T_423; // @[DCache.scala 820:29:freechips.rocketchip.system.DefaultRV32Config.fir@195596.4]
  assign io_cpu_resp_bits_data_word_bypass = {_T_600,_T_599}; // @[DCache.scala 874:37:freechips.rocketchip.system.DefaultRV32Config.fir@195703.4]
  assign io_cpu_resp_bits_data_raw = {_T_600,_T_599}; // @[DCache.scala 875:29:freechips.rocketchip.system.DefaultRV32Config.fir@195704.4]
  assign io_cpu_resp_bits_store_data = pstore1_data; // @[DCache.scala 876:31:freechips.rocketchip.system.DefaultRV32Config.fir@195705.4]
  assign io_cpu_replay_next = _T_2217 & grantIsUncachedData; // @[DCache.scala 849:22:freechips.rocketchip.system.DefaultRV32Config.fir@195652.4]
  assign io_cpu_s2_xcpt_ma_ld = _T_2470 & s2_tlb_xcpt_ma_ld; // @[DCache.scala 832:18:freechips.rocketchip.system.DefaultRV32Config.fir@195635.4]
  assign io_cpu_s2_xcpt_ma_st = _T_2470 & s2_tlb_xcpt_ma_st; // @[DCache.scala 832:18:freechips.rocketchip.system.DefaultRV32Config.fir@195635.4]
  assign io_cpu_s2_xcpt_pf_ld = _T_2470 & s2_tlb_xcpt_pf_ld; // @[DCache.scala 832:18:freechips.rocketchip.system.DefaultRV32Config.fir@195635.4]
  assign io_cpu_s2_xcpt_pf_st = _T_2470 & s2_tlb_xcpt_pf_st; // @[DCache.scala 832:18:freechips.rocketchip.system.DefaultRV32Config.fir@195635.4]
  assign io_cpu_s2_xcpt_ae_ld = _T_2470 & s2_tlb_xcpt_ae_ld; // @[DCache.scala 832:18:freechips.rocketchip.system.DefaultRV32Config.fir@195635.4]
  assign io_cpu_s2_xcpt_ae_st = _T_2470 & s2_tlb_xcpt_ae_st; // @[DCache.scala 832:18:freechips.rocketchip.system.DefaultRV32Config.fir@195635.4]
  assign io_cpu_ordered = ~_T_2465; // @[DCache.scala 829:18:freechips.rocketchip.system.DefaultRV32Config.fir@195611.4]
  assign io_cpu_perf_release = _T_2610 & _T_2354; // @[DCache.scala 978:23:freechips.rocketchip.system.DefaultRV32Config.fir@195851.4]
  assign io_cpu_perf_grant = auto_out_d_valid & d_last; // @[DCache.scala 979:21:freechips.rocketchip.system.DefaultRV32Config.fir@195853.4]
  assign io_ptw_req_valid = tlb_io_ptw_req_valid; // @[DCache.scala 230:10:freechips.rocketchip.system.DefaultRV32Config.fir@192520.4]
  assign io_ptw_req_bits_bits_addr = tlb_io_ptw_req_bits_bits_addr; // @[DCache.scala 230:10:freechips.rocketchip.system.DefaultRV32Config.fir@192520.4]
  assign tlb_clock = gated_clock; // @[:freechips.rocketchip.system.DefaultRV32Config.fir@192111.4]
  assign tlb_reset = reset; // @[:freechips.rocketchip.system.DefaultRV32Config.fir@192112.4]
  assign tlb_io_req_valid = s1_valid_masked & s1_cmd_uses_tlb; // @[DCache.scala 232:20:freechips.rocketchip.system.DefaultRV32Config.fir@192528.4]
  assign tlb_io_req_bits_vaddr = s1_tlb_req_vaddr; // @[DCache.scala 233:19:freechips.rocketchip.system.DefaultRV32Config.fir@192529.4]
  assign tlb_io_req_bits_passthrough = s1_tlb_req_passthrough; // @[DCache.scala 233:19:freechips.rocketchip.system.DefaultRV32Config.fir@192529.4]
  assign tlb_io_req_bits_size = s1_tlb_req_size; // @[DCache.scala 233:19:freechips.rocketchip.system.DefaultRV32Config.fir@192529.4]
  assign tlb_io_req_bits_cmd = s1_tlb_req_cmd; // @[DCache.scala 233:19:freechips.rocketchip.system.DefaultRV32Config.fir@192529.4]
  assign tlb_io_sfence_valid = s1_valid_masked & s1_sfence; // @[DCache.scala 237:23:freechips.rocketchip.system.DefaultRV32Config.fir@192548.4]
  assign tlb_io_sfence_bits_rs1 = s1_req_size[0]; // @[DCache.scala 238:26:freechips.rocketchip.system.DefaultRV32Config.fir@192550.4]
  assign tlb_io_sfence_bits_rs2 = s1_req_size[1]; // @[DCache.scala 239:26:freechips.rocketchip.system.DefaultRV32Config.fir@192552.4]
  assign tlb_io_sfence_bits_addr = s1_req_addr; // @[DCache.scala 241:27:freechips.rocketchip.system.DefaultRV32Config.fir@192554.4]
  assign tlb_io_ptw_req_ready = io_ptw_req_ready; // @[DCache.scala 230:10:freechips.rocketchip.system.DefaultRV32Config.fir@192520.4]
  assign tlb_io_ptw_resp_valid = io_ptw_resp_valid; // @[DCache.scala 230:10:freechips.rocketchip.system.DefaultRV32Config.fir@192520.4]
  assign tlb_io_ptw_resp_bits_ae = io_ptw_resp_bits_ae; // @[DCache.scala 230:10:freechips.rocketchip.system.DefaultRV32Config.fir@192520.4]
  assign tlb_io_ptw_resp_bits_pte_ppn = io_ptw_resp_bits_pte_ppn; // @[DCache.scala 230:10:freechips.rocketchip.system.DefaultRV32Config.fir@192520.4]
  assign tlb_io_ptw_resp_bits_pte_d = io_ptw_resp_bits_pte_d; // @[DCache.scala 230:10:freechips.rocketchip.system.DefaultRV32Config.fir@192520.4]
  assign tlb_io_ptw_resp_bits_pte_a = io_ptw_resp_bits_pte_a; // @[DCache.scala 230:10:freechips.rocketchip.system.DefaultRV32Config.fir@192520.4]
  assign tlb_io_ptw_resp_bits_pte_g = io_ptw_resp_bits_pte_g; // @[DCache.scala 230:10:freechips.rocketchip.system.DefaultRV32Config.fir@192520.4]
  assign tlb_io_ptw_resp_bits_pte_u = io_ptw_resp_bits_pte_u; // @[DCache.scala 230:10:freechips.rocketchip.system.DefaultRV32Config.fir@192520.4]
  assign tlb_io_ptw_resp_bits_pte_x = io_ptw_resp_bits_pte_x; // @[DCache.scala 230:10:freechips.rocketchip.system.DefaultRV32Config.fir@192520.4]
  assign tlb_io_ptw_resp_bits_pte_w = io_ptw_resp_bits_pte_w; // @[DCache.scala 230:10:freechips.rocketchip.system.DefaultRV32Config.fir@192520.4]
  assign tlb_io_ptw_resp_bits_pte_r = io_ptw_resp_bits_pte_r; // @[DCache.scala 230:10:freechips.rocketchip.system.DefaultRV32Config.fir@192520.4]
  assign tlb_io_ptw_resp_bits_pte_v = io_ptw_resp_bits_pte_v; // @[DCache.scala 230:10:freechips.rocketchip.system.DefaultRV32Config.fir@192520.4]
  assign tlb_io_ptw_resp_bits_level = io_ptw_resp_bits_level; // @[DCache.scala 230:10:freechips.rocketchip.system.DefaultRV32Config.fir@192520.4]
  assign tlb_io_ptw_resp_bits_homogeneous = io_ptw_resp_bits_homogeneous; // @[DCache.scala 230:10:freechips.rocketchip.system.DefaultRV32Config.fir@192520.4]
  assign tlb_io_ptw_ptbr_mode = io_ptw_ptbr_mode; // @[DCache.scala 230:10:freechips.rocketchip.system.DefaultRV32Config.fir@192520.4]
  assign tlb_io_ptw_status_debug = io_ptw_status_debug; // @[DCache.scala 230:10:freechips.rocketchip.system.DefaultRV32Config.fir@192520.4]
  assign tlb_io_ptw_status_dprv = io_ptw_status_dprv; // @[DCache.scala 230:10:freechips.rocketchip.system.DefaultRV32Config.fir@192520.4]
  assign tlb_io_ptw_status_mxr = io_ptw_status_mxr; // @[DCache.scala 230:10:freechips.rocketchip.system.DefaultRV32Config.fir@192520.4]
  assign tlb_io_ptw_status_sum = io_ptw_status_sum; // @[DCache.scala 230:10:freechips.rocketchip.system.DefaultRV32Config.fir@192520.4]
  assign tlb_io_ptw_pmp_0_cfg_l = io_ptw_pmp_0_cfg_l; // @[DCache.scala 230:10:freechips.rocketchip.system.DefaultRV32Config.fir@192520.4]
  assign tlb_io_ptw_pmp_0_cfg_a = io_ptw_pmp_0_cfg_a; // @[DCache.scala 230:10:freechips.rocketchip.system.DefaultRV32Config.fir@192520.4]
  assign tlb_io_ptw_pmp_0_cfg_x = io_ptw_pmp_0_cfg_x; // @[DCache.scala 230:10:freechips.rocketchip.system.DefaultRV32Config.fir@192520.4]
  assign tlb_io_ptw_pmp_0_cfg_w = io_ptw_pmp_0_cfg_w; // @[DCache.scala 230:10:freechips.rocketchip.system.DefaultRV32Config.fir@192520.4]
  assign tlb_io_ptw_pmp_0_cfg_r = io_ptw_pmp_0_cfg_r; // @[DCache.scala 230:10:freechips.rocketchip.system.DefaultRV32Config.fir@192520.4]
  assign tlb_io_ptw_pmp_0_addr = io_ptw_pmp_0_addr; // @[DCache.scala 230:10:freechips.rocketchip.system.DefaultRV32Config.fir@192520.4]
  assign tlb_io_ptw_pmp_0_mask = io_ptw_pmp_0_mask; // @[DCache.scala 230:10:freechips.rocketchip.system.DefaultRV32Config.fir@192520.4]
  assign tlb_io_ptw_pmp_1_cfg_l = io_ptw_pmp_1_cfg_l; // @[DCache.scala 230:10:freechips.rocketchip.system.DefaultRV32Config.fir@192520.4]
  assign tlb_io_ptw_pmp_1_cfg_a = io_ptw_pmp_1_cfg_a; // @[DCache.scala 230:10:freechips.rocketchip.system.DefaultRV32Config.fir@192520.4]
  assign tlb_io_ptw_pmp_1_cfg_x = io_ptw_pmp_1_cfg_x; // @[DCache.scala 230:10:freechips.rocketchip.system.DefaultRV32Config.fir@192520.4]
  assign tlb_io_ptw_pmp_1_cfg_w = io_ptw_pmp_1_cfg_w; // @[DCache.scala 230:10:freechips.rocketchip.system.DefaultRV32Config.fir@192520.4]
  assign tlb_io_ptw_pmp_1_cfg_r = io_ptw_pmp_1_cfg_r; // @[DCache.scala 230:10:freechips.rocketchip.system.DefaultRV32Config.fir@192520.4]
  assign tlb_io_ptw_pmp_1_addr = io_ptw_pmp_1_addr; // @[DCache.scala 230:10:freechips.rocketchip.system.DefaultRV32Config.fir@192520.4]
  assign tlb_io_ptw_pmp_1_mask = io_ptw_pmp_1_mask; // @[DCache.scala 230:10:freechips.rocketchip.system.DefaultRV32Config.fir@192520.4]
  assign tlb_io_ptw_pmp_2_cfg_l = io_ptw_pmp_2_cfg_l; // @[DCache.scala 230:10:freechips.rocketchip.system.DefaultRV32Config.fir@192520.4]
  assign tlb_io_ptw_pmp_2_cfg_a = io_ptw_pmp_2_cfg_a; // @[DCache.scala 230:10:freechips.rocketchip.system.DefaultRV32Config.fir@192520.4]
  assign tlb_io_ptw_pmp_2_cfg_x = io_ptw_pmp_2_cfg_x; // @[DCache.scala 230:10:freechips.rocketchip.system.DefaultRV32Config.fir@192520.4]
  assign tlb_io_ptw_pmp_2_cfg_w = io_ptw_pmp_2_cfg_w; // @[DCache.scala 230:10:freechips.rocketchip.system.DefaultRV32Config.fir@192520.4]
  assign tlb_io_ptw_pmp_2_cfg_r = io_ptw_pmp_2_cfg_r; // @[DCache.scala 230:10:freechips.rocketchip.system.DefaultRV32Config.fir@192520.4]
  assign tlb_io_ptw_pmp_2_addr = io_ptw_pmp_2_addr; // @[DCache.scala 230:10:freechips.rocketchip.system.DefaultRV32Config.fir@192520.4]
  assign tlb_io_ptw_pmp_2_mask = io_ptw_pmp_2_mask; // @[DCache.scala 230:10:freechips.rocketchip.system.DefaultRV32Config.fir@192520.4]
  assign tlb_io_ptw_pmp_3_cfg_l = io_ptw_pmp_3_cfg_l; // @[DCache.scala 230:10:freechips.rocketchip.system.DefaultRV32Config.fir@192520.4]
  assign tlb_io_ptw_pmp_3_cfg_a = io_ptw_pmp_3_cfg_a; // @[DCache.scala 230:10:freechips.rocketchip.system.DefaultRV32Config.fir@192520.4]
  assign tlb_io_ptw_pmp_3_cfg_x = io_ptw_pmp_3_cfg_x; // @[DCache.scala 230:10:freechips.rocketchip.system.DefaultRV32Config.fir@192520.4]
  assign tlb_io_ptw_pmp_3_cfg_w = io_ptw_pmp_3_cfg_w; // @[DCache.scala 230:10:freechips.rocketchip.system.DefaultRV32Config.fir@192520.4]
  assign tlb_io_ptw_pmp_3_cfg_r = io_ptw_pmp_3_cfg_r; // @[DCache.scala 230:10:freechips.rocketchip.system.DefaultRV32Config.fir@192520.4]
  assign tlb_io_ptw_pmp_3_addr = io_ptw_pmp_3_addr; // @[DCache.scala 230:10:freechips.rocketchip.system.DefaultRV32Config.fir@192520.4]
  assign tlb_io_ptw_pmp_3_mask = io_ptw_pmp_3_mask; // @[DCache.scala 230:10:freechips.rocketchip.system.DefaultRV32Config.fir@192520.4]
  assign tlb_io_ptw_pmp_4_cfg_l = io_ptw_pmp_4_cfg_l; // @[DCache.scala 230:10:freechips.rocketchip.system.DefaultRV32Config.fir@192520.4]
  assign tlb_io_ptw_pmp_4_cfg_a = io_ptw_pmp_4_cfg_a; // @[DCache.scala 230:10:freechips.rocketchip.system.DefaultRV32Config.fir@192520.4]
  assign tlb_io_ptw_pmp_4_cfg_x = io_ptw_pmp_4_cfg_x; // @[DCache.scala 230:10:freechips.rocketchip.system.DefaultRV32Config.fir@192520.4]
  assign tlb_io_ptw_pmp_4_cfg_w = io_ptw_pmp_4_cfg_w; // @[DCache.scala 230:10:freechips.rocketchip.system.DefaultRV32Config.fir@192520.4]
  assign tlb_io_ptw_pmp_4_cfg_r = io_ptw_pmp_4_cfg_r; // @[DCache.scala 230:10:freechips.rocketchip.system.DefaultRV32Config.fir@192520.4]
  assign tlb_io_ptw_pmp_4_addr = io_ptw_pmp_4_addr; // @[DCache.scala 230:10:freechips.rocketchip.system.DefaultRV32Config.fir@192520.4]
  assign tlb_io_ptw_pmp_4_mask = io_ptw_pmp_4_mask; // @[DCache.scala 230:10:freechips.rocketchip.system.DefaultRV32Config.fir@192520.4]
  assign tlb_io_ptw_pmp_5_cfg_l = io_ptw_pmp_5_cfg_l; // @[DCache.scala 230:10:freechips.rocketchip.system.DefaultRV32Config.fir@192520.4]
  assign tlb_io_ptw_pmp_5_cfg_a = io_ptw_pmp_5_cfg_a; // @[DCache.scala 230:10:freechips.rocketchip.system.DefaultRV32Config.fir@192520.4]
  assign tlb_io_ptw_pmp_5_cfg_x = io_ptw_pmp_5_cfg_x; // @[DCache.scala 230:10:freechips.rocketchip.system.DefaultRV32Config.fir@192520.4]
  assign tlb_io_ptw_pmp_5_cfg_w = io_ptw_pmp_5_cfg_w; // @[DCache.scala 230:10:freechips.rocketchip.system.DefaultRV32Config.fir@192520.4]
  assign tlb_io_ptw_pmp_5_cfg_r = io_ptw_pmp_5_cfg_r; // @[DCache.scala 230:10:freechips.rocketchip.system.DefaultRV32Config.fir@192520.4]
  assign tlb_io_ptw_pmp_5_addr = io_ptw_pmp_5_addr; // @[DCache.scala 230:10:freechips.rocketchip.system.DefaultRV32Config.fir@192520.4]
  assign tlb_io_ptw_pmp_5_mask = io_ptw_pmp_5_mask; // @[DCache.scala 230:10:freechips.rocketchip.system.DefaultRV32Config.fir@192520.4]
  assign tlb_io_ptw_pmp_6_cfg_l = io_ptw_pmp_6_cfg_l; // @[DCache.scala 230:10:freechips.rocketchip.system.DefaultRV32Config.fir@192520.4]
  assign tlb_io_ptw_pmp_6_cfg_a = io_ptw_pmp_6_cfg_a; // @[DCache.scala 230:10:freechips.rocketchip.system.DefaultRV32Config.fir@192520.4]
  assign tlb_io_ptw_pmp_6_cfg_x = io_ptw_pmp_6_cfg_x; // @[DCache.scala 230:10:freechips.rocketchip.system.DefaultRV32Config.fir@192520.4]
  assign tlb_io_ptw_pmp_6_cfg_w = io_ptw_pmp_6_cfg_w; // @[DCache.scala 230:10:freechips.rocketchip.system.DefaultRV32Config.fir@192520.4]
  assign tlb_io_ptw_pmp_6_cfg_r = io_ptw_pmp_6_cfg_r; // @[DCache.scala 230:10:freechips.rocketchip.system.DefaultRV32Config.fir@192520.4]
  assign tlb_io_ptw_pmp_6_addr = io_ptw_pmp_6_addr; // @[DCache.scala 230:10:freechips.rocketchip.system.DefaultRV32Config.fir@192520.4]
  assign tlb_io_ptw_pmp_6_mask = io_ptw_pmp_6_mask; // @[DCache.scala 230:10:freechips.rocketchip.system.DefaultRV32Config.fir@192520.4]
  assign tlb_io_ptw_pmp_7_cfg_l = io_ptw_pmp_7_cfg_l; // @[DCache.scala 230:10:freechips.rocketchip.system.DefaultRV32Config.fir@192520.4]
  assign tlb_io_ptw_pmp_7_cfg_a = io_ptw_pmp_7_cfg_a; // @[DCache.scala 230:10:freechips.rocketchip.system.DefaultRV32Config.fir@192520.4]
  assign tlb_io_ptw_pmp_7_cfg_x = io_ptw_pmp_7_cfg_x; // @[DCache.scala 230:10:freechips.rocketchip.system.DefaultRV32Config.fir@192520.4]
  assign tlb_io_ptw_pmp_7_cfg_w = io_ptw_pmp_7_cfg_w; // @[DCache.scala 230:10:freechips.rocketchip.system.DefaultRV32Config.fir@192520.4]
  assign tlb_io_ptw_pmp_7_cfg_r = io_ptw_pmp_7_cfg_r; // @[DCache.scala 230:10:freechips.rocketchip.system.DefaultRV32Config.fir@192520.4]
  assign tlb_io_ptw_pmp_7_addr = io_ptw_pmp_7_addr; // @[DCache.scala 230:10:freechips.rocketchip.system.DefaultRV32Config.fir@192520.4]
  assign tlb_io_ptw_pmp_7_mask = io_ptw_pmp_7_mask; // @[DCache.scala 230:10:freechips.rocketchip.system.DefaultRV32Config.fir@192520.4]
  assign MaxPeriodFibonacciLFSR_clock = gated_clock; // @[:freechips.rocketchip.system.DefaultRV32Config.fir@192120.4]
  assign MaxPeriodFibonacciLFSR_reset = reset; // @[:freechips.rocketchip.system.DefaultRV32Config.fir@192121.4]
  assign MaxPeriodFibonacciLFSR_io_increment = _T_2217 & _GEN_204; // @[PRNG.scala 85:23:freechips.rocketchip.system.DefaultRV32Config.fir@192139.4]
  assign metaArb_io_in_0_valid = resetting; // @[DCache.scala 947:26:freechips.rocketchip.system.DefaultRV32Config.fir@195756.4]
  assign metaArb_io_in_0_bits_addr = metaArb_io_in_5_bits_addr; // @[DCache.scala 948:25:freechips.rocketchip.system.DefaultRV32Config.fir@195757.4]
  assign metaArb_io_in_0_bits_idx = metaArb_io_in_5_bits_idx; // @[DCache.scala 948:25:freechips.rocketchip.system.DefaultRV32Config.fir@195757.4]
  assign metaArb_io_in_0_bits_data = {2'h0,s2_req_addr[31:12]}; // @[DCache.scala 948:25:freechips.rocketchip.system.DefaultRV32Config.fir@195757.4 DCache.scala 951:30:freechips.rocketchip.system.DefaultRV32Config.fir@195770.4]
  assign metaArb_io_in_1_valid = pma_checker__T_2026 & _T_792; // @[DCache.scala 401:26:freechips.rocketchip.system.DefaultRV32Config.fir@193378.4]
  assign metaArb_io_in_1_bits_addr = {io_cpu_req_bits_addr[31:12],_T_808}; // @[DCache.scala 405:30:freechips.rocketchip.system.DefaultRV32Config.fir@193398.4]
  assign metaArb_io_in_1_bits_idx = s2_probe ? probe_bits_address[11:6] : s2_vaddr[11:6]; // @[DCache.scala 404:29:freechips.rocketchip.system.DefaultRV32Config.fir@193394.4]
  assign metaArb_io_in_1_bits_data = {new_meta_coh_state,s2_meta_corrected_3_tag}; // @[DCache.scala 406:30:freechips.rocketchip.system.DefaultRV32Config.fir@193409.4]
  assign metaArb_io_in_2_valid = s2_valid_hit_pre_data_ecc_and_waw & s2_update_meta; // @[DCache.scala 413:26:freechips.rocketchip.system.DefaultRV32Config.fir@193411.4]
  assign metaArb_io_in_2_bits_addr = {io_cpu_req_bits_addr[31:12],s2_vaddr[11:0]}; // @[DCache.scala 417:30:freechips.rocketchip.system.DefaultRV32Config.fir@193420.4]
  assign metaArb_io_in_2_bits_idx = s2_vaddr[11:6]; // @[DCache.scala 416:29:freechips.rocketchip.system.DefaultRV32Config.fir@193416.4]
  assign metaArb_io_in_2_bits_way_en = s2_hit_valid ? s2_hit_way : _T_633; // @[DCache.scala 415:32:freechips.rocketchip.system.DefaultRV32Config.fir@193414.4]
  assign metaArb_io_in_2_bits_data = {s2_grow_param,s2_req_addr[31:12]}; // @[DCache.scala 418:30:freechips.rocketchip.system.DefaultRV32Config.fir@193427.4]
  assign metaArb_io_in_3_valid = _T_2254 & _T_2255; // @[DCache.scala 684:26:freechips.rocketchip.system.DefaultRV32Config.fir@195207.4]
  assign metaArb_io_in_3_bits_addr = {io_cpu_req_bits_addr[31:12],s2_vaddr[11:0]}; // @[DCache.scala 688:30:freechips.rocketchip.system.DefaultRV32Config.fir@195215.4]
  assign metaArb_io_in_3_bits_idx = s2_vaddr[11:6]; // @[DCache.scala 687:29:freechips.rocketchip.system.DefaultRV32Config.fir@195211.4]
  assign metaArb_io_in_3_bits_way_en = s2_hit_valid ? s2_hit_way : _T_633; // @[DCache.scala 686:32:freechips.rocketchip.system.DefaultRV32Config.fir@195209.4]
  assign metaArb_io_in_3_bits_data = {_T_2329,s2_req_addr[31:12]}; // @[DCache.scala 689:30:freechips.rocketchip.system.DefaultRV32Config.fir@195293.4]
  assign metaArb_io_in_4_valid = _T_2411 | _T_2446; // @[DCache.scala 810:26:freechips.rocketchip.system.DefaultRV32Config.fir@195575.4]
  assign metaArb_io_in_4_bits_addr = {io_cpu_req_bits_addr[31:12],probe_bits_address[11:0]}; // @[DCache.scala 814:30:freechips.rocketchip.system.DefaultRV32Config.fir@195583.4]
  assign metaArb_io_in_4_bits_idx = probe_bits_address[11:6]; // @[DCache.scala 813:29:freechips.rocketchip.system.DefaultRV32Config.fir@195579.4]
  assign metaArb_io_in_4_bits_way_en = _T_2412 ? s2_victim_way : s2_probe_way; // @[DCache.scala 812:32:freechips.rocketchip.system.DefaultRV32Config.fir@195577.4]
  assign metaArb_io_in_4_bits_data = {newCoh_state,probe_bits_address[31:12]}; // @[DCache.scala 815:30:freechips.rocketchip.system.DefaultRV32Config.fir@195590.4]
  assign metaArb_io_in_5_bits_addr = {io_cpu_req_bits_addr[31:12],_T_2542}; // @[DCache.scala 919:30:freechips.rocketchip.system.DefaultRV32Config.fir@195753.4]
  assign metaArb_io_in_5_bits_idx = flushCounter[5:0]; // @[DCache.scala 918:29:freechips.rocketchip.system.DefaultRV32Config.fir@195749.4]
  assign metaArb_io_in_6_valid = _T_2403 | _T_2345; // @[DCache.scala 712:26:freechips.rocketchip.system.DefaultRV32Config.fir@195321.4 DCache.scala 762:30:freechips.rocketchip.system.DefaultRV32Config.fir@195474.6]
  assign metaArb_io_in_6_bits_addr = _GEN_293[31:0]; // @[DCache.scala 716:30:freechips.rocketchip.system.DefaultRV32Config.fir@195333.4 DCache.scala 764:34:freechips.rocketchip.system.DefaultRV32Config.fir@195479.6]
  assign metaArb_io_in_6_bits_idx = _T_2403 ? probe_bits_address[11:6] : auto_out_b_bits_address[11:6]; // @[DCache.scala 715:29:freechips.rocketchip.system.DefaultRV32Config.fir@195330.4 DCache.scala 763:33:freechips.rocketchip.system.DefaultRV32Config.fir@195476.6]
  assign metaArb_io_in_6_bits_way_en = metaArb_io_in_4_bits_way_en; // @[DCache.scala 717:32:freechips.rocketchip.system.DefaultRV32Config.fir@195334.4]
  assign metaArb_io_in_6_bits_data = metaArb_io_in_4_bits_data; // @[DCache.scala 718:30:freechips.rocketchip.system.DefaultRV32Config.fir@195335.4]
  assign metaArb_io_in_7_valid = io_cpu_req_valid; // @[DCache.scala 220:26:freechips.rocketchip.system.DefaultRV32Config.fir@192506.4]
  assign metaArb_io_in_7_bits_addr = io_cpu_req_bits_addr; // @[DCache.scala 223:30:freechips.rocketchip.system.DefaultRV32Config.fir@192510.4]
  assign metaArb_io_in_7_bits_idx = io_cpu_req_bits_addr[11:6]; // @[DCache.scala 222:29:freechips.rocketchip.system.DefaultRV32Config.fir@192509.4]
  assign metaArb_io_in_7_bits_way_en = metaArb_io_in_4_bits_way_en; // @[DCache.scala 224:32:freechips.rocketchip.system.DefaultRV32Config.fir@192511.4]
  assign metaArb_io_in_7_bits_data = metaArb_io_in_4_bits_data; // @[DCache.scala 225:30:freechips.rocketchip.system.DefaultRV32Config.fir@192512.4]
  assign tag_array_RW0_wdata_0 = metaArb_io_out_bits_data; // @[:freechips.rocketchip.system.DefaultRV32Config.fir@192589.8]
  assign tag_array_RW0_wdata_1 = metaArb_io_out_bits_data; // @[:freechips.rocketchip.system.DefaultRV32Config.fir@192592.8]
  assign tag_array_RW0_wdata_2 = metaArb_io_out_bits_data; // @[:freechips.rocketchip.system.DefaultRV32Config.fir@192595.8]
  assign tag_array_RW0_wdata_3 = metaArb_io_out_bits_data; // @[:freechips.rocketchip.system.DefaultRV32Config.fir@192598.8]
  assign tag_array_RW0_wmask_0 = metaArb_io_out_bits_way_en[0]; // @[:freechips.rocketchip.system.DefaultRV32Config.fir@192587.6 :freechips.rocketchip.system.DefaultRV32Config.fir@192589.8]
  assign tag_array_RW0_wmask_1 = metaArb_io_out_bits_way_en[1]; // @[:freechips.rocketchip.system.DefaultRV32Config.fir@192587.6 :freechips.rocketchip.system.DefaultRV32Config.fir@192592.8]
  assign tag_array_RW0_wmask_2 = metaArb_io_out_bits_way_en[2]; // @[:freechips.rocketchip.system.DefaultRV32Config.fir@192587.6 :freechips.rocketchip.system.DefaultRV32Config.fir@192595.8]
  assign tag_array_RW0_wmask_3 = metaArb_io_out_bits_way_en[3]; // @[:freechips.rocketchip.system.DefaultRV32Config.fir@192587.6 :freechips.rocketchip.system.DefaultRV32Config.fir@192598.8]
  assign data_clock = gated_clock; // @[:freechips.rocketchip.system.DefaultRV32Config.fir@192162.4]
  assign data_io_req_valid = dataArb_io_out_valid; // @[DCache.scala 133:15:freechips.rocketchip.system.DefaultRV32Config.fir@192171.4]
  assign data_io_req_bits_addr = dataArb_io_out_bits_addr; // @[DCache.scala 133:15:freechips.rocketchip.system.DefaultRV32Config.fir@192171.4]
  assign data_io_req_bits_write = dataArb_io_out_bits_write; // @[DCache.scala 133:15:freechips.rocketchip.system.DefaultRV32Config.fir@192171.4]
  assign data_io_req_bits_wdata = dataArb_io_out_bits_wdata; // @[DCache.scala 133:15:freechips.rocketchip.system.DefaultRV32Config.fir@192171.4]
  assign data_io_req_bits_eccMask = dataArb_io_out_bits_eccMask; // @[DCache.scala 133:15:freechips.rocketchip.system.DefaultRV32Config.fir@192171.4]
  assign data_io_req_bits_way_en = dataArb_io_out_bits_way_en; // @[DCache.scala 133:15:freechips.rocketchip.system.DefaultRV32Config.fir@192171.4]
  assign dataArb_io_in_0_valid = pstore_drain_structural | _T_1008; // @[DCache.scala 498:26:freechips.rocketchip.system.DefaultRV32Config.fir@193779.4]
  assign dataArb_io_in_0_bits_addr = _T_1068[11:0]; // @[DCache.scala 500:30:freechips.rocketchip.system.DefaultRV32Config.fir@193782.4]
  assign dataArb_io_in_0_bits_write = pstore_drain_structural | _T_1008; // @[DCache.scala 499:31:freechips.rocketchip.system.DefaultRV32Config.fir@193780.4]
  assign dataArb_io_in_0_bits_wdata = {_T_1076,_T_1075}; // @[DCache.scala 502:31:freechips.rocketchip.system.DefaultRV32Config.fir@193793.4]
  assign dataArb_io_in_0_bits_eccMask = {_T_1090,_T_1089}; // @[DCache.scala 504:33:freechips.rocketchip.system.DefaultRV32Config.fir@193809.4]
  assign dataArb_io_in_0_bits_way_en = pstore2_valid ? pstore2_way : pstore1_way; // @[DCache.scala 501:32:freechips.rocketchip.system.DefaultRV32Config.fir@193784.4]
  assign dataArb_io_in_1_valid = _T_2334 ? _GEN_230 : _T_2246; // @[DCache.scala 664:26:freechips.rocketchip.system.DefaultRV32Config.fir@195186.4 DCache.scala 700:32:freechips.rocketchip.system.DefaultRV32Config.fir@195302.8]
  assign dataArb_io_in_1_bits_addr = _T_2251[11:0]; // @[DCache.scala 671:32:freechips.rocketchip.system.DefaultRV32Config.fir@195197.4]
  assign dataArb_io_in_1_bits_write = _T_2334 ? _GEN_231 : 1'h1; // @[DCache.scala 670:33:freechips.rocketchip.system.DefaultRV32Config.fir@195193.4 DCache.scala 701:37:freechips.rocketchip.system.DefaultRV32Config.fir@195303.8]
  assign dataArb_io_in_1_bits_wdata = {_T_327,_T_326}; // @[DCache.scala 132:43:freechips.rocketchip.system.DefaultRV32Config.fir@192168.4 DCache.scala 673:33:freechips.rocketchip.system.DefaultRV32Config.fir@195199.4]
  assign dataArb_io_in_1_bits_way_en = s2_hit_valid ? s2_hit_way : _T_633; // @[DCache.scala 672:34:freechips.rocketchip.system.DefaultRV32Config.fir@195198.4]
  assign dataArb_io_in_2_valid = inWriteback & _T_2436; // @[DCache.scala 803:26:freechips.rocketchip.system.DefaultRV32Config.fir@195559.4]
  assign dataArb_io_in_2_bits_addr = _T_2439 | _GEN_381; // @[DCache.scala 804:25:freechips.rocketchip.system.DefaultRV32Config.fir@195560.4 DCache.scala 806:30:freechips.rocketchip.system.DefaultRV32Config.fir@195567.4]
  assign dataArb_io_in_2_bits_wdata = dataArb_io_in_1_bits_wdata; // @[DCache.scala 132:43:freechips.rocketchip.system.DefaultRV32Config.fir@192169.4 DCache.scala 804:25:freechips.rocketchip.system.DefaultRV32Config.fir@195560.4]
  assign dataArb_io_in_3_valid = io_cpu_req_valid & res; // @[DCache.scala 212:26:freechips.rocketchip.system.DefaultRV32Config.fir@192436.4]
  assign dataArb_io_in_3_bits_addr = io_cpu_req_bits_addr[11:0]; // @[DCache.scala 213:25:freechips.rocketchip.system.DefaultRV32Config.fir@192437.4 DCache.scala 215:30:freechips.rocketchip.system.DefaultRV32Config.fir@192439.4]
  assign dataArb_io_in_3_bits_wdata = dataArb_io_in_1_bits_wdata; // @[DCache.scala 132:43:freechips.rocketchip.system.DefaultRV32Config.fir@192170.4 DCache.scala 213:25:freechips.rocketchip.system.DefaultRV32Config.fir@192437.4]
  assign amoalu_io_mask = pstore1_mask; // @[DCache.scala 882:22:freechips.rocketchip.system.DefaultRV32Config.fir@195711.4]
  assign amoalu_io_cmd = pstore1_cmd; // @[DCache.scala 883:21:freechips.rocketchip.system.DefaultRV32Config.fir@195712.4]
  assign amoalu_io_lhs = {_T_600,_T_599}; // @[DCache.scala 884:21:freechips.rocketchip.system.DefaultRV32Config.fir@195714.4]
  assign amoalu_io_rhs = pstore1_data; // @[DCache.scala 885:21:freechips.rocketchip.system.DefaultRV32Config.fir@195716.4]
  assign _GEN_385 = _T_2217 & grantIsCached; // @[DCache.scala 620:13:freechips.rocketchip.system.DefaultRV32Config.fir@195113.10]
  assign _GEN_388 = _T_2217 & _T_2725; // @[DCache.scala 630:17:freechips.rocketchip.system.DefaultRV32Config.fir@195132.14]
  assign _GEN_389 = _GEN_388 & grantIsUncached; // @[DCache.scala 630:17:freechips.rocketchip.system.DefaultRV32Config.fir@195132.14]
  assign _GEN_390 = _GEN_389 & _T_2222; // @[DCache.scala 630:17:freechips.rocketchip.system.DefaultRV32Config.fir@195132.14]
  assign _GEN_398 = _GEN_388 & _T_2192; // @[DCache.scala 651:13:freechips.rocketchip.system.DefaultRV32Config.fir@195158.14]
  assign _GEN_399 = _GEN_398 & grantIsVoluntary; // @[DCache.scala 651:13:freechips.rocketchip.system.DefaultRV32Config.fir@195158.14]
  assign tag_array_RW0_wmode = metaArb_io_out_bits_write;
  assign tag_array_RW0_clk = gated_clock;
  assign tag_array_RW0_en = s0_clk_en | _T_258;
  assign tag_array_RW0_addr = metaArb_io_out_bits_idx;
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  tlb_sectored_entries_0_tag = _RAND_0[19:0];
  _RAND_1 = {2{`RANDOM}};
  tlb_sectored_entries_0_data_0 = _RAND_1[34:0];
  _RAND_2 = {2{`RANDOM}};
  tlb_sectored_entries_0_data_1 = _RAND_2[34:0];
  _RAND_3 = {2{`RANDOM}};
  tlb_sectored_entries_0_data_2 = _RAND_3[34:0];
  _RAND_4 = {2{`RANDOM}};
  tlb_sectored_entries_0_data_3 = _RAND_4[34:0];
  _RAND_5 = {1{`RANDOM}};
  tlb_sectored_entries_0_valid_0 = _RAND_5[0:0];
  _RAND_6 = {1{`RANDOM}};
  tlb_sectored_entries_0_valid_1 = _RAND_6[0:0];
  _RAND_7 = {1{`RANDOM}};
  tlb_sectored_entries_0_valid_2 = _RAND_7[0:0];
  _RAND_8 = {1{`RANDOM}};
  tlb_sectored_entries_0_valid_3 = _RAND_8[0:0];
  _RAND_9 = {1{`RANDOM}};
  tlb_sectored_entries_1_tag = _RAND_9[19:0];
  _RAND_10 = {2{`RANDOM}};
  tlb_sectored_entries_1_data_0 = _RAND_10[34:0];
  _RAND_11 = {2{`RANDOM}};
  tlb_sectored_entries_1_data_1 = _RAND_11[34:0];
  _RAND_12 = {2{`RANDOM}};
  tlb_sectored_entries_1_data_2 = _RAND_12[34:0];
  _RAND_13 = {2{`RANDOM}};
  tlb_sectored_entries_1_data_3 = _RAND_13[34:0];
  _RAND_14 = {1{`RANDOM}};
  tlb_sectored_entries_1_valid_0 = _RAND_14[0:0];
  _RAND_15 = {1{`RANDOM}};
  tlb_sectored_entries_1_valid_1 = _RAND_15[0:0];
  _RAND_16 = {1{`RANDOM}};
  tlb_sectored_entries_1_valid_2 = _RAND_16[0:0];
  _RAND_17 = {1{`RANDOM}};
  tlb_sectored_entries_1_valid_3 = _RAND_17[0:0];
  _RAND_18 = {1{`RANDOM}};
  tlb_sectored_entries_2_tag = _RAND_18[19:0];
  _RAND_19 = {2{`RANDOM}};
  tlb_sectored_entries_2_data_0 = _RAND_19[34:0];
  _RAND_20 = {2{`RANDOM}};
  tlb_sectored_entries_2_data_1 = _RAND_20[34:0];
  _RAND_21 = {2{`RANDOM}};
  tlb_sectored_entries_2_data_2 = _RAND_21[34:0];
  _RAND_22 = {2{`RANDOM}};
  tlb_sectored_entries_2_data_3 = _RAND_22[34:0];
  _RAND_23 = {1{`RANDOM}};
  tlb_sectored_entries_2_valid_0 = _RAND_23[0:0];
  _RAND_24 = {1{`RANDOM}};
  tlb_sectored_entries_2_valid_1 = _RAND_24[0:0];
  _RAND_25 = {1{`RANDOM}};
  tlb_sectored_entries_2_valid_2 = _RAND_25[0:0];
  _RAND_26 = {1{`RANDOM}};
  tlb_sectored_entries_2_valid_3 = _RAND_26[0:0];
  _RAND_27 = {1{`RANDOM}};
  tlb_sectored_entries_3_tag = _RAND_27[19:0];
  _RAND_28 = {2{`RANDOM}};
  tlb_sectored_entries_3_data_0 = _RAND_28[34:0];
  _RAND_29 = {2{`RANDOM}};
  tlb_sectored_entries_3_data_1 = _RAND_29[34:0];
  _RAND_30 = {2{`RANDOM}};
  tlb_sectored_entries_3_data_2 = _RAND_30[34:0];
  _RAND_31 = {2{`RANDOM}};
  tlb_sectored_entries_3_data_3 = _RAND_31[34:0];
  _RAND_32 = {1{`RANDOM}};
  tlb_sectored_entries_3_valid_0 = _RAND_32[0:0];
  _RAND_33 = {1{`RANDOM}};
  tlb_sectored_entries_3_valid_1 = _RAND_33[0:0];
  _RAND_34 = {1{`RANDOM}};
  tlb_sectored_entries_3_valid_2 = _RAND_34[0:0];
  _RAND_35 = {1{`RANDOM}};
  tlb_sectored_entries_3_valid_3 = _RAND_35[0:0];
  _RAND_36 = {1{`RANDOM}};
  tlb_sectored_entries_4_tag = _RAND_36[19:0];
  _RAND_37 = {2{`RANDOM}};
  tlb_sectored_entries_4_data_0 = _RAND_37[34:0];
  _RAND_38 = {2{`RANDOM}};
  tlb_sectored_entries_4_data_1 = _RAND_38[34:0];
  _RAND_39 = {2{`RANDOM}};
  tlb_sectored_entries_4_data_2 = _RAND_39[34:0];
  _RAND_40 = {2{`RANDOM}};
  tlb_sectored_entries_4_data_3 = _RAND_40[34:0];
  _RAND_41 = {1{`RANDOM}};
  tlb_sectored_entries_4_valid_0 = _RAND_41[0:0];
  _RAND_42 = {1{`RANDOM}};
  tlb_sectored_entries_4_valid_1 = _RAND_42[0:0];
  _RAND_43 = {1{`RANDOM}};
  tlb_sectored_entries_4_valid_2 = _RAND_43[0:0];
  _RAND_44 = {1{`RANDOM}};
  tlb_sectored_entries_4_valid_3 = _RAND_44[0:0];
  _RAND_45 = {1{`RANDOM}};
  tlb_sectored_entries_5_tag = _RAND_45[19:0];
  _RAND_46 = {2{`RANDOM}};
  tlb_sectored_entries_5_data_0 = _RAND_46[34:0];
  _RAND_47 = {2{`RANDOM}};
  tlb_sectored_entries_5_data_1 = _RAND_47[34:0];
  _RAND_48 = {2{`RANDOM}};
  tlb_sectored_entries_5_data_2 = _RAND_48[34:0];
  _RAND_49 = {2{`RANDOM}};
  tlb_sectored_entries_5_data_3 = _RAND_49[34:0];
  _RAND_50 = {1{`RANDOM}};
  tlb_sectored_entries_5_valid_0 = _RAND_50[0:0];
  _RAND_51 = {1{`RANDOM}};
  tlb_sectored_entries_5_valid_1 = _RAND_51[0:0];
  _RAND_52 = {1{`RANDOM}};
  tlb_sectored_entries_5_valid_2 = _RAND_52[0:0];
  _RAND_53 = {1{`RANDOM}};
  tlb_sectored_entries_5_valid_3 = _RAND_53[0:0];
  _RAND_54 = {1{`RANDOM}};
  tlb_sectored_entries_6_tag = _RAND_54[19:0];
  _RAND_55 = {2{`RANDOM}};
  tlb_sectored_entries_6_data_0 = _RAND_55[34:0];
  _RAND_56 = {2{`RANDOM}};
  tlb_sectored_entries_6_data_1 = _RAND_56[34:0];
  _RAND_57 = {2{`RANDOM}};
  tlb_sectored_entries_6_data_2 = _RAND_57[34:0];
  _RAND_58 = {2{`RANDOM}};
  tlb_sectored_entries_6_data_3 = _RAND_58[34:0];
  _RAND_59 = {1{`RANDOM}};
  tlb_sectored_entries_6_valid_0 = _RAND_59[0:0];
  _RAND_60 = {1{`RANDOM}};
  tlb_sectored_entries_6_valid_1 = _RAND_60[0:0];
  _RAND_61 = {1{`RANDOM}};
  tlb_sectored_entries_6_valid_2 = _RAND_61[0:0];
  _RAND_62 = {1{`RANDOM}};
  tlb_sectored_entries_6_valid_3 = _RAND_62[0:0];
  _RAND_63 = {1{`RANDOM}};
  tlb_sectored_entries_7_tag = _RAND_63[19:0];
  _RAND_64 = {2{`RANDOM}};
  tlb_sectored_entries_7_data_0 = _RAND_64[34:0];
  _RAND_65 = {2{`RANDOM}};
  tlb_sectored_entries_7_data_1 = _RAND_65[34:0];
  _RAND_66 = {2{`RANDOM}};
  tlb_sectored_entries_7_data_2 = _RAND_66[34:0];
  _RAND_67 = {2{`RANDOM}};
  tlb_sectored_entries_7_data_3 = _RAND_67[34:0];
  _RAND_68 = {1{`RANDOM}};
  tlb_sectored_entries_7_valid_0 = _RAND_68[0:0];
  _RAND_69 = {1{`RANDOM}};
  tlb_sectored_entries_7_valid_1 = _RAND_69[0:0];
  _RAND_70 = {1{`RANDOM}};
  tlb_sectored_entries_7_valid_2 = _RAND_70[0:0];
  _RAND_71 = {1{`RANDOM}};
  tlb_sectored_entries_7_valid_3 = _RAND_71[0:0];
  _RAND_72 = {1{`RANDOM}};
  tlb_superpage_entries_0_tag = _RAND_72[19:0];
  _RAND_73 = {2{`RANDOM}};
  tlb_superpage_entries_0_data_0 = _RAND_73[34:0];
  _RAND_74 = {1{`RANDOM}};
  tlb_superpage_entries_0_valid_0 = _RAND_74[0:0];
  _RAND_75 = {1{`RANDOM}};
  tlb_superpage_entries_1_tag = _RAND_75[19:0];
  _RAND_76 = {2{`RANDOM}};
  tlb_superpage_entries_1_data_0 = _RAND_76[34:0];
  _RAND_77 = {1{`RANDOM}};
  tlb_superpage_entries_1_valid_0 = _RAND_77[0:0];
  _RAND_78 = {1{`RANDOM}};
  tlb_superpage_entries_2_tag = _RAND_78[19:0];
  _RAND_79 = {2{`RANDOM}};
  tlb_superpage_entries_2_data_0 = _RAND_79[34:0];
  _RAND_80 = {1{`RANDOM}};
  tlb_superpage_entries_2_valid_0 = _RAND_80[0:0];
  _RAND_81 = {1{`RANDOM}};
  tlb_superpage_entries_3_tag = _RAND_81[19:0];
  _RAND_82 = {2{`RANDOM}};
  tlb_superpage_entries_3_data_0 = _RAND_82[34:0];
  _RAND_83 = {1{`RANDOM}};
  tlb_superpage_entries_3_valid_0 = _RAND_83[0:0];
  _RAND_84 = {1{`RANDOM}};
  tlb_special_entry_level = _RAND_84[0:0];
  _RAND_85 = {1{`RANDOM}};
  tlb_special_entry_tag = _RAND_85[19:0];
  _RAND_86 = {2{`RANDOM}};
  tlb_special_entry_data_0 = _RAND_86[34:0];
  _RAND_87 = {1{`RANDOM}};
  tlb_special_entry_valid_0 = _RAND_87[0:0];
  _RAND_88 = {1{`RANDOM}};
  tlb_state = _RAND_88[1:0];
  _RAND_89 = {1{`RANDOM}};
  tlb_r_refill_tag = _RAND_89[19:0];
  _RAND_90 = {1{`RANDOM}};
  tlb_r_superpage_repl_addr = _RAND_90[1:0];
  _RAND_91 = {1{`RANDOM}};
  tlb_r_sectored_repl_addr = _RAND_91[2:0];
  _RAND_92 = {1{`RANDOM}};
  tlb_r_sectored_hit_addr = _RAND_92[2:0];
  _RAND_93 = {1{`RANDOM}};
  tlb_r_sectored_hit = _RAND_93[0:0];
  _RAND_94 = {1{`RANDOM}};
  tlb__T_2007 = _RAND_94[6:0];
  _RAND_95 = {1{`RANDOM}};
  tlb__T_2008 = _RAND_95[2:0];
  _RAND_96 = {1{`RANDOM}};
  s1_valid = _RAND_96[0:0];
  _RAND_97 = {1{`RANDOM}};
  blockProbeAfterGrantCount = _RAND_97[2:0];
  _RAND_98 = {1{`RANDOM}};
  lrscCount = _RAND_98[6:0];
  _RAND_99 = {1{`RANDOM}};
  s1_probe = _RAND_99[0:0];
  _RAND_100 = {1{`RANDOM}};
  s2_probe = _RAND_100[0:0];
  _RAND_101 = {1{`RANDOM}};
  release_state = _RAND_101[2:0];
  _RAND_102 = {1{`RANDOM}};
  release_ack_wait = _RAND_102[0:0];
  _RAND_103 = {1{`RANDOM}};
  release_ack_addr = _RAND_103[31:0];
  _RAND_104 = {1{`RANDOM}};
  grantInProgress = _RAND_104[0:0];
  _RAND_105 = {1{`RANDOM}};
  s2_valid = _RAND_105[0:0];
  _RAND_106 = {1{`RANDOM}};
  probe_bits_param = _RAND_106[1:0];
  _RAND_107 = {1{`RANDOM}};
  probe_bits_size = _RAND_107[3:0];
  _RAND_108 = {1{`RANDOM}};
  probe_bits_source = _RAND_108[0:0];
  _RAND_109 = {1{`RANDOM}};
  probe_bits_address = _RAND_109[31:0];
  _RAND_110 = {1{`RANDOM}};
  s2_probe_state_state = _RAND_110[1:0];
  _RAND_111 = {1{`RANDOM}};
  _T_2362 = _RAND_111[9:0];
  _RAND_112 = {1{`RANDOM}};
  s2_release_data_valid = _RAND_112[0:0];
  _RAND_113 = {1{`RANDOM}};
  s1_req_cmd = _RAND_113[4:0];
  _RAND_114 = {1{`RANDOM}};
  s2_req_cmd = _RAND_114[4:0];
  _RAND_115 = {1{`RANDOM}};
  pstore1_held = _RAND_115[0:0];
  _RAND_116 = {1{`RANDOM}};
  pstore1_addr = _RAND_116[31:0];
  _RAND_117 = {1{`RANDOM}};
  s1_req_addr = _RAND_117[31:0];
  _RAND_118 = {1{`RANDOM}};
  pstore1_mask = _RAND_118[3:0];
  _RAND_119 = {1{`RANDOM}};
  s1_req_size = _RAND_119[1:0];
  _RAND_120 = {1{`RANDOM}};
  pstore2_valid = _RAND_120[0:0];
  _RAND_121 = {1{`RANDOM}};
  pstore2_addr = _RAND_121[31:0];
  _RAND_122 = {1{`RANDOM}};
  mask = _RAND_122[3:0];
  _RAND_123 = {1{`RANDOM}};
  s2_not_nacked_in_s1 = _RAND_123[0:0];
  _RAND_124 = {1{`RANDOM}};
  s2_hit_state_state = _RAND_124[1:0];
  _RAND_125 = {1{`RANDOM}};
  s1_req_tag = _RAND_125[6:0];
  _RAND_126 = {1{`RANDOM}};
  s1_req_signed = _RAND_126[0:0];
  _RAND_127 = {1{`RANDOM}};
  s1_req_dprv = _RAND_127[1:0];
  _RAND_128 = {1{`RANDOM}};
  s1_tlb_req_vaddr = _RAND_128[31:0];
  _RAND_129 = {1{`RANDOM}};
  s1_tlb_req_passthrough = _RAND_129[0:0];
  _RAND_130 = {1{`RANDOM}};
  s1_tlb_req_size = _RAND_130[1:0];
  _RAND_131 = {1{`RANDOM}};
  s1_tlb_req_cmd = _RAND_131[4:0];
  _RAND_132 = {1{`RANDOM}};
  cached_grant_wait = _RAND_132[0:0];
  _RAND_133 = {1{`RANDOM}};
  uncachedInFlight_0 = _RAND_133[0:0];
  _RAND_134 = {1{`RANDOM}};
  uncachedReqs_0_addr = _RAND_134[31:0];
  _RAND_135 = {1{`RANDOM}};
  uncachedReqs_0_tag = _RAND_135[6:0];
  _RAND_136 = {1{`RANDOM}};
  uncachedReqs_0_size = _RAND_136[1:0];
  _RAND_137 = {1{`RANDOM}};
  uncachedReqs_0_signed = _RAND_137[0:0];
  _RAND_138 = {1{`RANDOM}};
  s1_did_read = _RAND_138[0:0];
  _RAND_139 = {1{`RANDOM}};
  s2_hit_way = _RAND_139[3:0];
  _RAND_140 = {1{`RANDOM}};
  _T_632 = _RAND_140[1:0];
  _RAND_141 = {1{`RANDOM}};
  s2_probe_way = _RAND_141[3:0];
  _RAND_142 = {1{`RANDOM}};
  s2_req_addr = _RAND_142[31:0];
  _RAND_143 = {1{`RANDOM}};
  s2_req_tag = _RAND_143[6:0];
  _RAND_144 = {1{`RANDOM}};
  s2_req_size = _RAND_144[1:0];
  _RAND_145 = {1{`RANDOM}};
  s2_req_signed = _RAND_145[0:0];
  _RAND_146 = {1{`RANDOM}};
  s2_req_dprv = _RAND_146[1:0];
  _RAND_147 = {1{`RANDOM}};
  s2_tlb_xcpt_pf_ld = _RAND_147[0:0];
  _RAND_148 = {1{`RANDOM}};
  s2_tlb_xcpt_pf_st = _RAND_148[0:0];
  _RAND_149 = {1{`RANDOM}};
  s2_tlb_xcpt_ae_ld = _RAND_149[0:0];
  _RAND_150 = {1{`RANDOM}};
  s2_tlb_xcpt_ae_st = _RAND_150[0:0];
  _RAND_151 = {1{`RANDOM}};
  s2_tlb_xcpt_ma_ld = _RAND_151[0:0];
  _RAND_152 = {1{`RANDOM}};
  s2_tlb_xcpt_ma_st = _RAND_152[0:0];
  _RAND_153 = {1{`RANDOM}};
  s2_pma_cacheable = _RAND_153[0:0];
  _RAND_154 = {1{`RANDOM}};
  s2_uncached_resp_addr = _RAND_154[31:0];
  _RAND_155 = {1{`RANDOM}};
  _T_377 = _RAND_155[31:0];
  _RAND_156 = {1{`RANDOM}};
  _T_449 = _RAND_156[21:0];
  _RAND_157 = {1{`RANDOM}};
  blockUncachedGrant = _RAND_157[0:0];
  _RAND_158 = {1{`RANDOM}};
  _T_2177 = _RAND_158[9:0];
  _RAND_159 = {1{`RANDOM}};
  s2_data = _RAND_159[31:0];
  _RAND_160 = {1{`RANDOM}};
  _T_637 = _RAND_160[19:0];
  _RAND_161 = {1{`RANDOM}};
  _T_639_state = _RAND_161[1:0];
  _RAND_162 = {1{`RANDOM}};
  lrscAddr = _RAND_162[25:0];
  _RAND_163 = {1{`RANDOM}};
  pstore1_cmd = _RAND_163[4:0];
  _RAND_164 = {1{`RANDOM}};
  pstore1_data = _RAND_164[31:0];
  _RAND_165 = {1{`RANDOM}};
  pstore1_way = _RAND_165[3:0];
  _RAND_166 = {1{`RANDOM}};
  pstore1_rmw = _RAND_166[0:0];
  _RAND_167 = {1{`RANDOM}};
  _T_976 = _RAND_167[0:0];
  _RAND_168 = {1{`RANDOM}};
  pstore2_way = _RAND_168[3:0];
  _RAND_169 = {1{`RANDOM}};
  _T_1032 = _RAND_169[7:0];
  _RAND_170 = {1{`RANDOM}};
  _T_1037 = _RAND_170[7:0];
  _RAND_171 = {1{`RANDOM}};
  _T_1042 = _RAND_171[7:0];
  _RAND_172 = {1{`RANDOM}};
  _T_1047 = _RAND_172[7:0];
  _RAND_173 = {1{`RANDOM}};
  s1_release_data_valid = _RAND_173[0:0];
  _RAND_174 = {1{`RANDOM}};
  _T_2470 = _RAND_174[0:0];
  _RAND_175 = {1{`RANDOM}};
  doUncachedResp = _RAND_175[0:0];
  _RAND_176 = {1{`RANDOM}};
  resetting = _RAND_176[0:0];
  _RAND_177 = {1{`RANDOM}};
  _T_2523 = _RAND_177[0:0];
  _RAND_178 = {1{`RANDOM}};
  flushCounter = _RAND_178[7:0];
  _RAND_179 = {1{`RANDOM}};
  _T_2604 = _RAND_179[9:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge tlb_clock) begin
    if (tlb__T_939) begin
      if (!(tlb__T_961)) begin
        if (!(tlb__T_979)) begin
          if (tlb__T_1045) begin
            tlb_sectored_entries_0_tag <= tlb_r_refill_tag;
          end
        end
      end
    end
    if (tlb__T_939) begin
      if (!(tlb__T_961)) begin
        if (!(tlb__T_979)) begin
          if (tlb__T_1045) begin
            if (2'h0 == tlb__T_1047) begin
              tlb_sectored_entries_0_data_0 <= tlb__T_978;
            end
          end
        end
      end
    end
    if (tlb__T_939) begin
      if (!(tlb__T_961)) begin
        if (!(tlb__T_979)) begin
          if (tlb__T_1045) begin
            if (2'h1 == tlb__T_1047) begin
              tlb_sectored_entries_0_data_1 <= tlb__T_978;
            end
          end
        end
      end
    end
    if (tlb__T_939) begin
      if (!(tlb__T_961)) begin
        if (!(tlb__T_979)) begin
          if (tlb__T_1045) begin
            if (2'h2 == tlb__T_1047) begin
              tlb_sectored_entries_0_data_2 <= tlb__T_978;
            end
          end
        end
      end
    end
    if (tlb__T_939) begin
      if (!(tlb__T_961)) begin
        if (!(tlb__T_979)) begin
          if (tlb__T_1045) begin
            if (2'h3 == tlb__T_1047) begin
              tlb_sectored_entries_0_data_3 <= tlb__T_978;
            end
          end
        end
      end
    end
    if (tlb__T_3753) begin
      tlb_sectored_entries_0_valid_0 <= 1'h0;
    end else if (tlb_io_sfence_valid) begin
      if (tlb_io_sfence_bits_rs1) begin
        if (tlb__T_2353) begin
          if (tlb__T_2356) begin
            tlb_sectored_entries_0_valid_0 <= 1'h0;
          end else if (tlb__T_415) begin
            if (2'h0 == tlb__T_510) begin
              tlb_sectored_entries_0_valid_0 <= 1'h0;
            end else if (tlb__T_939) begin
              if (!(tlb__T_961)) begin
                if (!(tlb__T_979)) begin
                  if (tlb__T_1045) begin
                    tlb_sectored_entries_0_valid_0 <= tlb__GEN_84;
                  end
                end
              end
            end
          end else if (tlb__T_939) begin
            if (!(tlb__T_961)) begin
              if (!(tlb__T_979)) begin
                if (tlb__T_1045) begin
                  tlb_sectored_entries_0_valid_0 <= tlb__GEN_84;
                end
              end
            end
          end
        end else if (tlb__T_415) begin
          if (2'h0 == tlb__T_510) begin
            tlb_sectored_entries_0_valid_0 <= 1'h0;
          end else if (tlb__T_939) begin
            if (!(tlb__T_961)) begin
              if (!(tlb__T_979)) begin
                if (tlb__T_1045) begin
                  tlb_sectored_entries_0_valid_0 <= tlb__GEN_84;
                end
              end
            end
          end
        end else if (tlb__T_939) begin
          if (!(tlb__T_961)) begin
            if (!(tlb__T_979)) begin
              if (tlb__T_1045) begin
                tlb_sectored_entries_0_valid_0 <= tlb__GEN_84;
              end
            end
          end
        end
      end else begin
        tlb_sectored_entries_0_valid_0 <= tlb__GEN_652;
      end
    end else begin
      tlb_sectored_entries_0_valid_0 <= tlb__GEN_472;
    end
    if (tlb__T_3753) begin
      tlb_sectored_entries_0_valid_1 <= 1'h0;
    end else if (tlb_io_sfence_valid) begin
      if (tlb_io_sfence_bits_rs1) begin
        if (tlb__T_2353) begin
          if (tlb__T_2374) begin
            tlb_sectored_entries_0_valid_1 <= 1'h0;
          end else if (tlb__T_415) begin
            if (2'h1 == tlb__T_510) begin
              tlb_sectored_entries_0_valid_1 <= 1'h0;
            end else if (tlb__T_939) begin
              if (!(tlb__T_961)) begin
                if (!(tlb__T_979)) begin
                  if (tlb__T_1045) begin
                    tlb_sectored_entries_0_valid_1 <= tlb__GEN_85;
                  end
                end
              end
            end
          end else if (tlb__T_939) begin
            if (!(tlb__T_961)) begin
              if (!(tlb__T_979)) begin
                if (tlb__T_1045) begin
                  tlb_sectored_entries_0_valid_1 <= tlb__GEN_85;
                end
              end
            end
          end
        end else if (tlb__T_415) begin
          if (2'h1 == tlb__T_510) begin
            tlb_sectored_entries_0_valid_1 <= 1'h0;
          end else if (tlb__T_939) begin
            if (!(tlb__T_961)) begin
              if (!(tlb__T_979)) begin
                if (tlb__T_1045) begin
                  tlb_sectored_entries_0_valid_1 <= tlb__GEN_85;
                end
              end
            end
          end
        end else if (tlb__T_939) begin
          if (!(tlb__T_961)) begin
            if (!(tlb__T_979)) begin
              if (tlb__T_1045) begin
                tlb_sectored_entries_0_valid_1 <= tlb__GEN_85;
              end
            end
          end
        end
      end else begin
        tlb_sectored_entries_0_valid_1 <= tlb__GEN_653;
      end
    end else begin
      tlb_sectored_entries_0_valid_1 <= tlb__GEN_473;
    end
    if (tlb__T_3753) begin
      tlb_sectored_entries_0_valid_2 <= 1'h0;
    end else if (tlb_io_sfence_valid) begin
      if (tlb_io_sfence_bits_rs1) begin
        if (tlb__T_2353) begin
          if (tlb__T_2392) begin
            tlb_sectored_entries_0_valid_2 <= 1'h0;
          end else if (tlb__T_415) begin
            if (2'h2 == tlb__T_510) begin
              tlb_sectored_entries_0_valid_2 <= 1'h0;
            end else if (tlb__T_939) begin
              if (!(tlb__T_961)) begin
                if (!(tlb__T_979)) begin
                  if (tlb__T_1045) begin
                    tlb_sectored_entries_0_valid_2 <= tlb__GEN_86;
                  end
                end
              end
            end
          end else if (tlb__T_939) begin
            if (!(tlb__T_961)) begin
              if (!(tlb__T_979)) begin
                if (tlb__T_1045) begin
                  tlb_sectored_entries_0_valid_2 <= tlb__GEN_86;
                end
              end
            end
          end
        end else if (tlb__T_415) begin
          if (2'h2 == tlb__T_510) begin
            tlb_sectored_entries_0_valid_2 <= 1'h0;
          end else if (tlb__T_939) begin
            if (!(tlb__T_961)) begin
              if (!(tlb__T_979)) begin
                if (tlb__T_1045) begin
                  tlb_sectored_entries_0_valid_2 <= tlb__GEN_86;
                end
              end
            end
          end
        end else if (tlb__T_939) begin
          if (!(tlb__T_961)) begin
            if (!(tlb__T_979)) begin
              if (tlb__T_1045) begin
                tlb_sectored_entries_0_valid_2 <= tlb__GEN_86;
              end
            end
          end
        end
      end else begin
        tlb_sectored_entries_0_valid_2 <= tlb__GEN_654;
      end
    end else begin
      tlb_sectored_entries_0_valid_2 <= tlb__GEN_474;
    end
    if (tlb__T_3753) begin
      tlb_sectored_entries_0_valid_3 <= 1'h0;
    end else if (tlb_io_sfence_valid) begin
      if (tlb_io_sfence_bits_rs1) begin
        if (tlb__T_2353) begin
          if (tlb__T_2410) begin
            tlb_sectored_entries_0_valid_3 <= 1'h0;
          end else if (tlb__T_415) begin
            if (2'h3 == tlb__T_510) begin
              tlb_sectored_entries_0_valid_3 <= 1'h0;
            end else if (tlb__T_939) begin
              if (!(tlb__T_961)) begin
                if (!(tlb__T_979)) begin
                  if (tlb__T_1045) begin
                    tlb_sectored_entries_0_valid_3 <= tlb__GEN_87;
                  end
                end
              end
            end
          end else if (tlb__T_939) begin
            if (!(tlb__T_961)) begin
              if (!(tlb__T_979)) begin
                if (tlb__T_1045) begin
                  tlb_sectored_entries_0_valid_3 <= tlb__GEN_87;
                end
              end
            end
          end
        end else if (tlb__T_415) begin
          if (2'h3 == tlb__T_510) begin
            tlb_sectored_entries_0_valid_3 <= 1'h0;
          end else if (tlb__T_939) begin
            if (!(tlb__T_961)) begin
              if (!(tlb__T_979)) begin
                if (tlb__T_1045) begin
                  tlb_sectored_entries_0_valid_3 <= tlb__GEN_87;
                end
              end
            end
          end
        end else if (tlb__T_939) begin
          if (!(tlb__T_961)) begin
            if (!(tlb__T_979)) begin
              if (tlb__T_1045) begin
                tlb_sectored_entries_0_valid_3 <= tlb__GEN_87;
              end
            end
          end
        end
      end else begin
        tlb_sectored_entries_0_valid_3 <= tlb__GEN_655;
      end
    end else begin
      tlb_sectored_entries_0_valid_3 <= tlb__GEN_475;
    end
    if (tlb__T_939) begin
      if (!(tlb__T_961)) begin
        if (!(tlb__T_979)) begin
          if (tlb__T_1063) begin
            tlb_sectored_entries_1_tag <= tlb_r_refill_tag;
          end
        end
      end
    end
    if (tlb__T_939) begin
      if (!(tlb__T_961)) begin
        if (!(tlb__T_979)) begin
          if (tlb__T_1063) begin
            if (2'h0 == tlb__T_1047) begin
              tlb_sectored_entries_1_data_0 <= tlb__T_978;
            end
          end
        end
      end
    end
    if (tlb__T_939) begin
      if (!(tlb__T_961)) begin
        if (!(tlb__T_979)) begin
          if (tlb__T_1063) begin
            if (2'h1 == tlb__T_1047) begin
              tlb_sectored_entries_1_data_1 <= tlb__T_978;
            end
          end
        end
      end
    end
    if (tlb__T_939) begin
      if (!(tlb__T_961)) begin
        if (!(tlb__T_979)) begin
          if (tlb__T_1063) begin
            if (2'h2 == tlb__T_1047) begin
              tlb_sectored_entries_1_data_2 <= tlb__T_978;
            end
          end
        end
      end
    end
    if (tlb__T_939) begin
      if (!(tlb__T_961)) begin
        if (!(tlb__T_979)) begin
          if (tlb__T_1063) begin
            if (2'h3 == tlb__T_1047) begin
              tlb_sectored_entries_1_data_3 <= tlb__T_978;
            end
          end
        end
      end
    end
    if (tlb__T_3753) begin
      tlb_sectored_entries_1_valid_0 <= 1'h0;
    end else if (tlb_io_sfence_valid) begin
      if (tlb_io_sfence_bits_rs1) begin
        if (tlb__T_2508) begin
          if (tlb__T_2511) begin
            tlb_sectored_entries_1_valid_0 <= 1'h0;
          end else if (tlb__T_421) begin
            if (2'h0 == tlb__T_510) begin
              tlb_sectored_entries_1_valid_0 <= 1'h0;
            end else if (tlb__T_939) begin
              if (!(tlb__T_961)) begin
                if (!(tlb__T_979)) begin
                  if (tlb__T_1063) begin
                    tlb_sectored_entries_1_valid_0 <= tlb__GEN_106;
                  end
                end
              end
            end
          end else if (tlb__T_939) begin
            if (!(tlb__T_961)) begin
              if (!(tlb__T_979)) begin
                if (tlb__T_1063) begin
                  tlb_sectored_entries_1_valid_0 <= tlb__GEN_106;
                end
              end
            end
          end
        end else if (tlb__T_421) begin
          if (2'h0 == tlb__T_510) begin
            tlb_sectored_entries_1_valid_0 <= 1'h0;
          end else if (tlb__T_939) begin
            if (!(tlb__T_961)) begin
              if (!(tlb__T_979)) begin
                if (tlb__T_1063) begin
                  tlb_sectored_entries_1_valid_0 <= tlb__GEN_106;
                end
              end
            end
          end
        end else if (tlb__T_939) begin
          if (!(tlb__T_961)) begin
            if (!(tlb__T_979)) begin
              if (tlb__T_1063) begin
                tlb_sectored_entries_1_valid_0 <= tlb__GEN_106;
              end
            end
          end
        end
      end else begin
        tlb_sectored_entries_1_valid_0 <= tlb__GEN_680;
      end
    end else begin
      tlb_sectored_entries_1_valid_0 <= tlb__GEN_482;
    end
    if (tlb__T_3753) begin
      tlb_sectored_entries_1_valid_1 <= 1'h0;
    end else if (tlb_io_sfence_valid) begin
      if (tlb_io_sfence_bits_rs1) begin
        if (tlb__T_2508) begin
          if (tlb__T_2529) begin
            tlb_sectored_entries_1_valid_1 <= 1'h0;
          end else if (tlb__T_421) begin
            if (2'h1 == tlb__T_510) begin
              tlb_sectored_entries_1_valid_1 <= 1'h0;
            end else if (tlb__T_939) begin
              if (!(tlb__T_961)) begin
                if (!(tlb__T_979)) begin
                  if (tlb__T_1063) begin
                    tlb_sectored_entries_1_valid_1 <= tlb__GEN_107;
                  end
                end
              end
            end
          end else if (tlb__T_939) begin
            if (!(tlb__T_961)) begin
              if (!(tlb__T_979)) begin
                if (tlb__T_1063) begin
                  tlb_sectored_entries_1_valid_1 <= tlb__GEN_107;
                end
              end
            end
          end
        end else if (tlb__T_421) begin
          if (2'h1 == tlb__T_510) begin
            tlb_sectored_entries_1_valid_1 <= 1'h0;
          end else if (tlb__T_939) begin
            if (!(tlb__T_961)) begin
              if (!(tlb__T_979)) begin
                if (tlb__T_1063) begin
                  tlb_sectored_entries_1_valid_1 <= tlb__GEN_107;
                end
              end
            end
          end
        end else if (tlb__T_939) begin
          if (!(tlb__T_961)) begin
            if (!(tlb__T_979)) begin
              if (tlb__T_1063) begin
                tlb_sectored_entries_1_valid_1 <= tlb__GEN_107;
              end
            end
          end
        end
      end else begin
        tlb_sectored_entries_1_valid_1 <= tlb__GEN_681;
      end
    end else begin
      tlb_sectored_entries_1_valid_1 <= tlb__GEN_483;
    end
    if (tlb__T_3753) begin
      tlb_sectored_entries_1_valid_2 <= 1'h0;
    end else if (tlb_io_sfence_valid) begin
      if (tlb_io_sfence_bits_rs1) begin
        if (tlb__T_2508) begin
          if (tlb__T_2547) begin
            tlb_sectored_entries_1_valid_2 <= 1'h0;
          end else if (tlb__T_421) begin
            if (2'h2 == tlb__T_510) begin
              tlb_sectored_entries_1_valid_2 <= 1'h0;
            end else if (tlb__T_939) begin
              if (!(tlb__T_961)) begin
                if (!(tlb__T_979)) begin
                  if (tlb__T_1063) begin
                    tlb_sectored_entries_1_valid_2 <= tlb__GEN_108;
                  end
                end
              end
            end
          end else if (tlb__T_939) begin
            if (!(tlb__T_961)) begin
              if (!(tlb__T_979)) begin
                if (tlb__T_1063) begin
                  tlb_sectored_entries_1_valid_2 <= tlb__GEN_108;
                end
              end
            end
          end
        end else if (tlb__T_421) begin
          if (2'h2 == tlb__T_510) begin
            tlb_sectored_entries_1_valid_2 <= 1'h0;
          end else if (tlb__T_939) begin
            if (!(tlb__T_961)) begin
              if (!(tlb__T_979)) begin
                if (tlb__T_1063) begin
                  tlb_sectored_entries_1_valid_2 <= tlb__GEN_108;
                end
              end
            end
          end
        end else if (tlb__T_939) begin
          if (!(tlb__T_961)) begin
            if (!(tlb__T_979)) begin
              if (tlb__T_1063) begin
                tlb_sectored_entries_1_valid_2 <= tlb__GEN_108;
              end
            end
          end
        end
      end else begin
        tlb_sectored_entries_1_valid_2 <= tlb__GEN_682;
      end
    end else begin
      tlb_sectored_entries_1_valid_2 <= tlb__GEN_484;
    end
    if (tlb__T_3753) begin
      tlb_sectored_entries_1_valid_3 <= 1'h0;
    end else if (tlb_io_sfence_valid) begin
      if (tlb_io_sfence_bits_rs1) begin
        if (tlb__T_2508) begin
          if (tlb__T_2565) begin
            tlb_sectored_entries_1_valid_3 <= 1'h0;
          end else if (tlb__T_421) begin
            if (2'h3 == tlb__T_510) begin
              tlb_sectored_entries_1_valid_3 <= 1'h0;
            end else if (tlb__T_939) begin
              if (!(tlb__T_961)) begin
                if (!(tlb__T_979)) begin
                  if (tlb__T_1063) begin
                    tlb_sectored_entries_1_valid_3 <= tlb__GEN_109;
                  end
                end
              end
            end
          end else if (tlb__T_939) begin
            if (!(tlb__T_961)) begin
              if (!(tlb__T_979)) begin
                if (tlb__T_1063) begin
                  tlb_sectored_entries_1_valid_3 <= tlb__GEN_109;
                end
              end
            end
          end
        end else if (tlb__T_421) begin
          if (2'h3 == tlb__T_510) begin
            tlb_sectored_entries_1_valid_3 <= 1'h0;
          end else if (tlb__T_939) begin
            if (!(tlb__T_961)) begin
              if (!(tlb__T_979)) begin
                if (tlb__T_1063) begin
                  tlb_sectored_entries_1_valid_3 <= tlb__GEN_109;
                end
              end
            end
          end
        end else if (tlb__T_939) begin
          if (!(tlb__T_961)) begin
            if (!(tlb__T_979)) begin
              if (tlb__T_1063) begin
                tlb_sectored_entries_1_valid_3 <= tlb__GEN_109;
              end
            end
          end
        end
      end else begin
        tlb_sectored_entries_1_valid_3 <= tlb__GEN_683;
      end
    end else begin
      tlb_sectored_entries_1_valid_3 <= tlb__GEN_485;
    end
    if (tlb__T_939) begin
      if (!(tlb__T_961)) begin
        if (!(tlb__T_979)) begin
          if (tlb__T_1081) begin
            tlb_sectored_entries_2_tag <= tlb_r_refill_tag;
          end
        end
      end
    end
    if (tlb__T_939) begin
      if (!(tlb__T_961)) begin
        if (!(tlb__T_979)) begin
          if (tlb__T_1081) begin
            if (2'h0 == tlb__T_1047) begin
              tlb_sectored_entries_2_data_0 <= tlb__T_978;
            end
          end
        end
      end
    end
    if (tlb__T_939) begin
      if (!(tlb__T_961)) begin
        if (!(tlb__T_979)) begin
          if (tlb__T_1081) begin
            if (2'h1 == tlb__T_1047) begin
              tlb_sectored_entries_2_data_1 <= tlb__T_978;
            end
          end
        end
      end
    end
    if (tlb__T_939) begin
      if (!(tlb__T_961)) begin
        if (!(tlb__T_979)) begin
          if (tlb__T_1081) begin
            if (2'h2 == tlb__T_1047) begin
              tlb_sectored_entries_2_data_2 <= tlb__T_978;
            end
          end
        end
      end
    end
    if (tlb__T_939) begin
      if (!(tlb__T_961)) begin
        if (!(tlb__T_979)) begin
          if (tlb__T_1081) begin
            if (2'h3 == tlb__T_1047) begin
              tlb_sectored_entries_2_data_3 <= tlb__T_978;
            end
          end
        end
      end
    end
    if (tlb__T_3753) begin
      tlb_sectored_entries_2_valid_0 <= 1'h0;
    end else if (tlb_io_sfence_valid) begin
      if (tlb_io_sfence_bits_rs1) begin
        if (tlb__T_2663) begin
          if (tlb__T_2666) begin
            tlb_sectored_entries_2_valid_0 <= 1'h0;
          end else if (tlb__T_427) begin
            if (2'h0 == tlb__T_510) begin
              tlb_sectored_entries_2_valid_0 <= 1'h0;
            end else if (tlb__T_939) begin
              if (!(tlb__T_961)) begin
                if (!(tlb__T_979)) begin
                  if (tlb__T_1081) begin
                    tlb_sectored_entries_2_valid_0 <= tlb__GEN_128;
                  end
                end
              end
            end
          end else if (tlb__T_939) begin
            if (!(tlb__T_961)) begin
              if (!(tlb__T_979)) begin
                if (tlb__T_1081) begin
                  tlb_sectored_entries_2_valid_0 <= tlb__GEN_128;
                end
              end
            end
          end
        end else if (tlb__T_427) begin
          if (2'h0 == tlb__T_510) begin
            tlb_sectored_entries_2_valid_0 <= 1'h0;
          end else if (tlb__T_939) begin
            if (!(tlb__T_961)) begin
              if (!(tlb__T_979)) begin
                if (tlb__T_1081) begin
                  tlb_sectored_entries_2_valid_0 <= tlb__GEN_128;
                end
              end
            end
          end
        end else if (tlb__T_939) begin
          if (!(tlb__T_961)) begin
            if (!(tlb__T_979)) begin
              if (tlb__T_1081) begin
                tlb_sectored_entries_2_valid_0 <= tlb__GEN_128;
              end
            end
          end
        end
      end else begin
        tlb_sectored_entries_2_valid_0 <= tlb__GEN_708;
      end
    end else begin
      tlb_sectored_entries_2_valid_0 <= tlb__GEN_492;
    end
    if (tlb__T_3753) begin
      tlb_sectored_entries_2_valid_1 <= 1'h0;
    end else if (tlb_io_sfence_valid) begin
      if (tlb_io_sfence_bits_rs1) begin
        if (tlb__T_2663) begin
          if (tlb__T_2684) begin
            tlb_sectored_entries_2_valid_1 <= 1'h0;
          end else if (tlb__T_427) begin
            if (2'h1 == tlb__T_510) begin
              tlb_sectored_entries_2_valid_1 <= 1'h0;
            end else if (tlb__T_939) begin
              if (!(tlb__T_961)) begin
                if (!(tlb__T_979)) begin
                  if (tlb__T_1081) begin
                    tlb_sectored_entries_2_valid_1 <= tlb__GEN_129;
                  end
                end
              end
            end
          end else if (tlb__T_939) begin
            if (!(tlb__T_961)) begin
              if (!(tlb__T_979)) begin
                if (tlb__T_1081) begin
                  tlb_sectored_entries_2_valid_1 <= tlb__GEN_129;
                end
              end
            end
          end
        end else if (tlb__T_427) begin
          if (2'h1 == tlb__T_510) begin
            tlb_sectored_entries_2_valid_1 <= 1'h0;
          end else if (tlb__T_939) begin
            if (!(tlb__T_961)) begin
              if (!(tlb__T_979)) begin
                if (tlb__T_1081) begin
                  tlb_sectored_entries_2_valid_1 <= tlb__GEN_129;
                end
              end
            end
          end
        end else if (tlb__T_939) begin
          if (!(tlb__T_961)) begin
            if (!(tlb__T_979)) begin
              if (tlb__T_1081) begin
                tlb_sectored_entries_2_valid_1 <= tlb__GEN_129;
              end
            end
          end
        end
      end else begin
        tlb_sectored_entries_2_valid_1 <= tlb__GEN_709;
      end
    end else begin
      tlb_sectored_entries_2_valid_1 <= tlb__GEN_493;
    end
    if (tlb__T_3753) begin
      tlb_sectored_entries_2_valid_2 <= 1'h0;
    end else if (tlb_io_sfence_valid) begin
      if (tlb_io_sfence_bits_rs1) begin
        if (tlb__T_2663) begin
          if (tlb__T_2702) begin
            tlb_sectored_entries_2_valid_2 <= 1'h0;
          end else if (tlb__T_427) begin
            if (2'h2 == tlb__T_510) begin
              tlb_sectored_entries_2_valid_2 <= 1'h0;
            end else if (tlb__T_939) begin
              if (!(tlb__T_961)) begin
                if (!(tlb__T_979)) begin
                  if (tlb__T_1081) begin
                    tlb_sectored_entries_2_valid_2 <= tlb__GEN_130;
                  end
                end
              end
            end
          end else if (tlb__T_939) begin
            if (!(tlb__T_961)) begin
              if (!(tlb__T_979)) begin
                if (tlb__T_1081) begin
                  tlb_sectored_entries_2_valid_2 <= tlb__GEN_130;
                end
              end
            end
          end
        end else if (tlb__T_427) begin
          if (2'h2 == tlb__T_510) begin
            tlb_sectored_entries_2_valid_2 <= 1'h0;
          end else if (tlb__T_939) begin
            if (!(tlb__T_961)) begin
              if (!(tlb__T_979)) begin
                if (tlb__T_1081) begin
                  tlb_sectored_entries_2_valid_2 <= tlb__GEN_130;
                end
              end
            end
          end
        end else if (tlb__T_939) begin
          if (!(tlb__T_961)) begin
            if (!(tlb__T_979)) begin
              if (tlb__T_1081) begin
                tlb_sectored_entries_2_valid_2 <= tlb__GEN_130;
              end
            end
          end
        end
      end else begin
        tlb_sectored_entries_2_valid_2 <= tlb__GEN_710;
      end
    end else begin
      tlb_sectored_entries_2_valid_2 <= tlb__GEN_494;
    end
    if (tlb__T_3753) begin
      tlb_sectored_entries_2_valid_3 <= 1'h0;
    end else if (tlb_io_sfence_valid) begin
      if (tlb_io_sfence_bits_rs1) begin
        if (tlb__T_2663) begin
          if (tlb__T_2720) begin
            tlb_sectored_entries_2_valid_3 <= 1'h0;
          end else if (tlb__T_427) begin
            if (2'h3 == tlb__T_510) begin
              tlb_sectored_entries_2_valid_3 <= 1'h0;
            end else if (tlb__T_939) begin
              if (!(tlb__T_961)) begin
                if (!(tlb__T_979)) begin
                  if (tlb__T_1081) begin
                    tlb_sectored_entries_2_valid_3 <= tlb__GEN_131;
                  end
                end
              end
            end
          end else if (tlb__T_939) begin
            if (!(tlb__T_961)) begin
              if (!(tlb__T_979)) begin
                if (tlb__T_1081) begin
                  tlb_sectored_entries_2_valid_3 <= tlb__GEN_131;
                end
              end
            end
          end
        end else if (tlb__T_427) begin
          if (2'h3 == tlb__T_510) begin
            tlb_sectored_entries_2_valid_3 <= 1'h0;
          end else if (tlb__T_939) begin
            if (!(tlb__T_961)) begin
              if (!(tlb__T_979)) begin
                if (tlb__T_1081) begin
                  tlb_sectored_entries_2_valid_3 <= tlb__GEN_131;
                end
              end
            end
          end
        end else if (tlb__T_939) begin
          if (!(tlb__T_961)) begin
            if (!(tlb__T_979)) begin
              if (tlb__T_1081) begin
                tlb_sectored_entries_2_valid_3 <= tlb__GEN_131;
              end
            end
          end
        end
      end else begin
        tlb_sectored_entries_2_valid_3 <= tlb__GEN_711;
      end
    end else begin
      tlb_sectored_entries_2_valid_3 <= tlb__GEN_495;
    end
    if (tlb__T_939) begin
      if (!(tlb__T_961)) begin
        if (!(tlb__T_979)) begin
          if (tlb__T_1099) begin
            tlb_sectored_entries_3_tag <= tlb_r_refill_tag;
          end
        end
      end
    end
    if (tlb__T_939) begin
      if (!(tlb__T_961)) begin
        if (!(tlb__T_979)) begin
          if (tlb__T_1099) begin
            if (2'h0 == tlb__T_1047) begin
              tlb_sectored_entries_3_data_0 <= tlb__T_978;
            end
          end
        end
      end
    end
    if (tlb__T_939) begin
      if (!(tlb__T_961)) begin
        if (!(tlb__T_979)) begin
          if (tlb__T_1099) begin
            if (2'h1 == tlb__T_1047) begin
              tlb_sectored_entries_3_data_1 <= tlb__T_978;
            end
          end
        end
      end
    end
    if (tlb__T_939) begin
      if (!(tlb__T_961)) begin
        if (!(tlb__T_979)) begin
          if (tlb__T_1099) begin
            if (2'h2 == tlb__T_1047) begin
              tlb_sectored_entries_3_data_2 <= tlb__T_978;
            end
          end
        end
      end
    end
    if (tlb__T_939) begin
      if (!(tlb__T_961)) begin
        if (!(tlb__T_979)) begin
          if (tlb__T_1099) begin
            if (2'h3 == tlb__T_1047) begin
              tlb_sectored_entries_3_data_3 <= tlb__T_978;
            end
          end
        end
      end
    end
    if (tlb__T_3753) begin
      tlb_sectored_entries_3_valid_0 <= 1'h0;
    end else if (tlb_io_sfence_valid) begin
      if (tlb_io_sfence_bits_rs1) begin
        if (tlb__T_2818) begin
          if (tlb__T_2821) begin
            tlb_sectored_entries_3_valid_0 <= 1'h0;
          end else if (tlb__T_433) begin
            if (2'h0 == tlb__T_510) begin
              tlb_sectored_entries_3_valid_0 <= 1'h0;
            end else if (tlb__T_939) begin
              if (!(tlb__T_961)) begin
                if (!(tlb__T_979)) begin
                  if (tlb__T_1099) begin
                    tlb_sectored_entries_3_valid_0 <= tlb__GEN_150;
                  end
                end
              end
            end
          end else if (tlb__T_939) begin
            if (!(tlb__T_961)) begin
              if (!(tlb__T_979)) begin
                if (tlb__T_1099) begin
                  tlb_sectored_entries_3_valid_0 <= tlb__GEN_150;
                end
              end
            end
          end
        end else if (tlb__T_433) begin
          if (2'h0 == tlb__T_510) begin
            tlb_sectored_entries_3_valid_0 <= 1'h0;
          end else if (tlb__T_939) begin
            if (!(tlb__T_961)) begin
              if (!(tlb__T_979)) begin
                if (tlb__T_1099) begin
                  tlb_sectored_entries_3_valid_0 <= tlb__GEN_150;
                end
              end
            end
          end
        end else if (tlb__T_939) begin
          if (!(tlb__T_961)) begin
            if (!(tlb__T_979)) begin
              if (tlb__T_1099) begin
                tlb_sectored_entries_3_valid_0 <= tlb__GEN_150;
              end
            end
          end
        end
      end else begin
        tlb_sectored_entries_3_valid_0 <= tlb__GEN_736;
      end
    end else begin
      tlb_sectored_entries_3_valid_0 <= tlb__GEN_502;
    end
    if (tlb__T_3753) begin
      tlb_sectored_entries_3_valid_1 <= 1'h0;
    end else if (tlb_io_sfence_valid) begin
      if (tlb_io_sfence_bits_rs1) begin
        if (tlb__T_2818) begin
          if (tlb__T_2839) begin
            tlb_sectored_entries_3_valid_1 <= 1'h0;
          end else if (tlb__T_433) begin
            if (2'h1 == tlb__T_510) begin
              tlb_sectored_entries_3_valid_1 <= 1'h0;
            end else if (tlb__T_939) begin
              if (!(tlb__T_961)) begin
                if (!(tlb__T_979)) begin
                  if (tlb__T_1099) begin
                    tlb_sectored_entries_3_valid_1 <= tlb__GEN_151;
                  end
                end
              end
            end
          end else if (tlb__T_939) begin
            if (!(tlb__T_961)) begin
              if (!(tlb__T_979)) begin
                if (tlb__T_1099) begin
                  tlb_sectored_entries_3_valid_1 <= tlb__GEN_151;
                end
              end
            end
          end
        end else if (tlb__T_433) begin
          if (2'h1 == tlb__T_510) begin
            tlb_sectored_entries_3_valid_1 <= 1'h0;
          end else if (tlb__T_939) begin
            if (!(tlb__T_961)) begin
              if (!(tlb__T_979)) begin
                if (tlb__T_1099) begin
                  tlb_sectored_entries_3_valid_1 <= tlb__GEN_151;
                end
              end
            end
          end
        end else if (tlb__T_939) begin
          if (!(tlb__T_961)) begin
            if (!(tlb__T_979)) begin
              if (tlb__T_1099) begin
                tlb_sectored_entries_3_valid_1 <= tlb__GEN_151;
              end
            end
          end
        end
      end else begin
        tlb_sectored_entries_3_valid_1 <= tlb__GEN_737;
      end
    end else begin
      tlb_sectored_entries_3_valid_1 <= tlb__GEN_503;
    end
    if (tlb__T_3753) begin
      tlb_sectored_entries_3_valid_2 <= 1'h0;
    end else if (tlb_io_sfence_valid) begin
      if (tlb_io_sfence_bits_rs1) begin
        if (tlb__T_2818) begin
          if (tlb__T_2857) begin
            tlb_sectored_entries_3_valid_2 <= 1'h0;
          end else if (tlb__T_433) begin
            if (2'h2 == tlb__T_510) begin
              tlb_sectored_entries_3_valid_2 <= 1'h0;
            end else if (tlb__T_939) begin
              if (!(tlb__T_961)) begin
                if (!(tlb__T_979)) begin
                  if (tlb__T_1099) begin
                    tlb_sectored_entries_3_valid_2 <= tlb__GEN_152;
                  end
                end
              end
            end
          end else if (tlb__T_939) begin
            if (!(tlb__T_961)) begin
              if (!(tlb__T_979)) begin
                if (tlb__T_1099) begin
                  tlb_sectored_entries_3_valid_2 <= tlb__GEN_152;
                end
              end
            end
          end
        end else if (tlb__T_433) begin
          if (2'h2 == tlb__T_510) begin
            tlb_sectored_entries_3_valid_2 <= 1'h0;
          end else if (tlb__T_939) begin
            if (!(tlb__T_961)) begin
              if (!(tlb__T_979)) begin
                if (tlb__T_1099) begin
                  tlb_sectored_entries_3_valid_2 <= tlb__GEN_152;
                end
              end
            end
          end
        end else if (tlb__T_939) begin
          if (!(tlb__T_961)) begin
            if (!(tlb__T_979)) begin
              if (tlb__T_1099) begin
                tlb_sectored_entries_3_valid_2 <= tlb__GEN_152;
              end
            end
          end
        end
      end else begin
        tlb_sectored_entries_3_valid_2 <= tlb__GEN_738;
      end
    end else begin
      tlb_sectored_entries_3_valid_2 <= tlb__GEN_504;
    end
    if (tlb__T_3753) begin
      tlb_sectored_entries_3_valid_3 <= 1'h0;
    end else if (tlb_io_sfence_valid) begin
      if (tlb_io_sfence_bits_rs1) begin
        if (tlb__T_2818) begin
          if (tlb__T_2875) begin
            tlb_sectored_entries_3_valid_3 <= 1'h0;
          end else if (tlb__T_433) begin
            if (2'h3 == tlb__T_510) begin
              tlb_sectored_entries_3_valid_3 <= 1'h0;
            end else if (tlb__T_939) begin
              if (!(tlb__T_961)) begin
                if (!(tlb__T_979)) begin
                  if (tlb__T_1099) begin
                    tlb_sectored_entries_3_valid_3 <= tlb__GEN_153;
                  end
                end
              end
            end
          end else if (tlb__T_939) begin
            if (!(tlb__T_961)) begin
              if (!(tlb__T_979)) begin
                if (tlb__T_1099) begin
                  tlb_sectored_entries_3_valid_3 <= tlb__GEN_153;
                end
              end
            end
          end
        end else if (tlb__T_433) begin
          if (2'h3 == tlb__T_510) begin
            tlb_sectored_entries_3_valid_3 <= 1'h0;
          end else if (tlb__T_939) begin
            if (!(tlb__T_961)) begin
              if (!(tlb__T_979)) begin
                if (tlb__T_1099) begin
                  tlb_sectored_entries_3_valid_3 <= tlb__GEN_153;
                end
              end
            end
          end
        end else if (tlb__T_939) begin
          if (!(tlb__T_961)) begin
            if (!(tlb__T_979)) begin
              if (tlb__T_1099) begin
                tlb_sectored_entries_3_valid_3 <= tlb__GEN_153;
              end
            end
          end
        end
      end else begin
        tlb_sectored_entries_3_valid_3 <= tlb__GEN_739;
      end
    end else begin
      tlb_sectored_entries_3_valid_3 <= tlb__GEN_505;
    end
    if (tlb__T_939) begin
      if (!(tlb__T_961)) begin
        if (!(tlb__T_979)) begin
          if (tlb__T_1117) begin
            tlb_sectored_entries_4_tag <= tlb_r_refill_tag;
          end
        end
      end
    end
    if (tlb__T_939) begin
      if (!(tlb__T_961)) begin
        if (!(tlb__T_979)) begin
          if (tlb__T_1117) begin
            if (2'h0 == tlb__T_1047) begin
              tlb_sectored_entries_4_data_0 <= tlb__T_978;
            end
          end
        end
      end
    end
    if (tlb__T_939) begin
      if (!(tlb__T_961)) begin
        if (!(tlb__T_979)) begin
          if (tlb__T_1117) begin
            if (2'h1 == tlb__T_1047) begin
              tlb_sectored_entries_4_data_1 <= tlb__T_978;
            end
          end
        end
      end
    end
    if (tlb__T_939) begin
      if (!(tlb__T_961)) begin
        if (!(tlb__T_979)) begin
          if (tlb__T_1117) begin
            if (2'h2 == tlb__T_1047) begin
              tlb_sectored_entries_4_data_2 <= tlb__T_978;
            end
          end
        end
      end
    end
    if (tlb__T_939) begin
      if (!(tlb__T_961)) begin
        if (!(tlb__T_979)) begin
          if (tlb__T_1117) begin
            if (2'h3 == tlb__T_1047) begin
              tlb_sectored_entries_4_data_3 <= tlb__T_978;
            end
          end
        end
      end
    end
    if (tlb__T_3753) begin
      tlb_sectored_entries_4_valid_0 <= 1'h0;
    end else if (tlb_io_sfence_valid) begin
      if (tlb_io_sfence_bits_rs1) begin
        if (tlb__T_2973) begin
          if (tlb__T_2976) begin
            tlb_sectored_entries_4_valid_0 <= 1'h0;
          end else if (tlb__T_439) begin
            if (2'h0 == tlb__T_510) begin
              tlb_sectored_entries_4_valid_0 <= 1'h0;
            end else if (tlb__T_939) begin
              if (!(tlb__T_961)) begin
                if (!(tlb__T_979)) begin
                  if (tlb__T_1117) begin
                    tlb_sectored_entries_4_valid_0 <= tlb__GEN_172;
                  end
                end
              end
            end
          end else if (tlb__T_939) begin
            if (!(tlb__T_961)) begin
              if (!(tlb__T_979)) begin
                if (tlb__T_1117) begin
                  tlb_sectored_entries_4_valid_0 <= tlb__GEN_172;
                end
              end
            end
          end
        end else if (tlb__T_439) begin
          if (2'h0 == tlb__T_510) begin
            tlb_sectored_entries_4_valid_0 <= 1'h0;
          end else if (tlb__T_939) begin
            if (!(tlb__T_961)) begin
              if (!(tlb__T_979)) begin
                if (tlb__T_1117) begin
                  tlb_sectored_entries_4_valid_0 <= tlb__GEN_172;
                end
              end
            end
          end
        end else if (tlb__T_939) begin
          if (!(tlb__T_961)) begin
            if (!(tlb__T_979)) begin
              if (tlb__T_1117) begin
                tlb_sectored_entries_4_valid_0 <= tlb__GEN_172;
              end
            end
          end
        end
      end else begin
        tlb_sectored_entries_4_valid_0 <= tlb__GEN_764;
      end
    end else begin
      tlb_sectored_entries_4_valid_0 <= tlb__GEN_512;
    end
    if (tlb__T_3753) begin
      tlb_sectored_entries_4_valid_1 <= 1'h0;
    end else if (tlb_io_sfence_valid) begin
      if (tlb_io_sfence_bits_rs1) begin
        if (tlb__T_2973) begin
          if (tlb__T_2994) begin
            tlb_sectored_entries_4_valid_1 <= 1'h0;
          end else if (tlb__T_439) begin
            if (2'h1 == tlb__T_510) begin
              tlb_sectored_entries_4_valid_1 <= 1'h0;
            end else if (tlb__T_939) begin
              if (!(tlb__T_961)) begin
                if (!(tlb__T_979)) begin
                  if (tlb__T_1117) begin
                    tlb_sectored_entries_4_valid_1 <= tlb__GEN_173;
                  end
                end
              end
            end
          end else if (tlb__T_939) begin
            if (!(tlb__T_961)) begin
              if (!(tlb__T_979)) begin
                if (tlb__T_1117) begin
                  tlb_sectored_entries_4_valid_1 <= tlb__GEN_173;
                end
              end
            end
          end
        end else if (tlb__T_439) begin
          if (2'h1 == tlb__T_510) begin
            tlb_sectored_entries_4_valid_1 <= 1'h0;
          end else if (tlb__T_939) begin
            if (!(tlb__T_961)) begin
              if (!(tlb__T_979)) begin
                if (tlb__T_1117) begin
                  tlb_sectored_entries_4_valid_1 <= tlb__GEN_173;
                end
              end
            end
          end
        end else if (tlb__T_939) begin
          if (!(tlb__T_961)) begin
            if (!(tlb__T_979)) begin
              if (tlb__T_1117) begin
                tlb_sectored_entries_4_valid_1 <= tlb__GEN_173;
              end
            end
          end
        end
      end else begin
        tlb_sectored_entries_4_valid_1 <= tlb__GEN_765;
      end
    end else begin
      tlb_sectored_entries_4_valid_1 <= tlb__GEN_513;
    end
    if (tlb__T_3753) begin
      tlb_sectored_entries_4_valid_2 <= 1'h0;
    end else if (tlb_io_sfence_valid) begin
      if (tlb_io_sfence_bits_rs1) begin
        if (tlb__T_2973) begin
          if (tlb__T_3012) begin
            tlb_sectored_entries_4_valid_2 <= 1'h0;
          end else if (tlb__T_439) begin
            if (2'h2 == tlb__T_510) begin
              tlb_sectored_entries_4_valid_2 <= 1'h0;
            end else if (tlb__T_939) begin
              if (!(tlb__T_961)) begin
                if (!(tlb__T_979)) begin
                  if (tlb__T_1117) begin
                    tlb_sectored_entries_4_valid_2 <= tlb__GEN_174;
                  end
                end
              end
            end
          end else if (tlb__T_939) begin
            if (!(tlb__T_961)) begin
              if (!(tlb__T_979)) begin
                if (tlb__T_1117) begin
                  tlb_sectored_entries_4_valid_2 <= tlb__GEN_174;
                end
              end
            end
          end
        end else if (tlb__T_439) begin
          if (2'h2 == tlb__T_510) begin
            tlb_sectored_entries_4_valid_2 <= 1'h0;
          end else if (tlb__T_939) begin
            if (!(tlb__T_961)) begin
              if (!(tlb__T_979)) begin
                if (tlb__T_1117) begin
                  tlb_sectored_entries_4_valid_2 <= tlb__GEN_174;
                end
              end
            end
          end
        end else if (tlb__T_939) begin
          if (!(tlb__T_961)) begin
            if (!(tlb__T_979)) begin
              if (tlb__T_1117) begin
                tlb_sectored_entries_4_valid_2 <= tlb__GEN_174;
              end
            end
          end
        end
      end else begin
        tlb_sectored_entries_4_valid_2 <= tlb__GEN_766;
      end
    end else begin
      tlb_sectored_entries_4_valid_2 <= tlb__GEN_514;
    end
    if (tlb__T_3753) begin
      tlb_sectored_entries_4_valid_3 <= 1'h0;
    end else if (tlb_io_sfence_valid) begin
      if (tlb_io_sfence_bits_rs1) begin
        if (tlb__T_2973) begin
          if (tlb__T_3030) begin
            tlb_sectored_entries_4_valid_3 <= 1'h0;
          end else if (tlb__T_439) begin
            if (2'h3 == tlb__T_510) begin
              tlb_sectored_entries_4_valid_3 <= 1'h0;
            end else if (tlb__T_939) begin
              if (!(tlb__T_961)) begin
                if (!(tlb__T_979)) begin
                  if (tlb__T_1117) begin
                    tlb_sectored_entries_4_valid_3 <= tlb__GEN_175;
                  end
                end
              end
            end
          end else if (tlb__T_939) begin
            if (!(tlb__T_961)) begin
              if (!(tlb__T_979)) begin
                if (tlb__T_1117) begin
                  tlb_sectored_entries_4_valid_3 <= tlb__GEN_175;
                end
              end
            end
          end
        end else if (tlb__T_439) begin
          if (2'h3 == tlb__T_510) begin
            tlb_sectored_entries_4_valid_3 <= 1'h0;
          end else if (tlb__T_939) begin
            if (!(tlb__T_961)) begin
              if (!(tlb__T_979)) begin
                if (tlb__T_1117) begin
                  tlb_sectored_entries_4_valid_3 <= tlb__GEN_175;
                end
              end
            end
          end
        end else if (tlb__T_939) begin
          if (!(tlb__T_961)) begin
            if (!(tlb__T_979)) begin
              if (tlb__T_1117) begin
                tlb_sectored_entries_4_valid_3 <= tlb__GEN_175;
              end
            end
          end
        end
      end else begin
        tlb_sectored_entries_4_valid_3 <= tlb__GEN_767;
      end
    end else begin
      tlb_sectored_entries_4_valid_3 <= tlb__GEN_515;
    end
    if (tlb__T_939) begin
      if (!(tlb__T_961)) begin
        if (!(tlb__T_979)) begin
          if (tlb__T_1135) begin
            tlb_sectored_entries_5_tag <= tlb_r_refill_tag;
          end
        end
      end
    end
    if (tlb__T_939) begin
      if (!(tlb__T_961)) begin
        if (!(tlb__T_979)) begin
          if (tlb__T_1135) begin
            if (2'h0 == tlb__T_1047) begin
              tlb_sectored_entries_5_data_0 <= tlb__T_978;
            end
          end
        end
      end
    end
    if (tlb__T_939) begin
      if (!(tlb__T_961)) begin
        if (!(tlb__T_979)) begin
          if (tlb__T_1135) begin
            if (2'h1 == tlb__T_1047) begin
              tlb_sectored_entries_5_data_1 <= tlb__T_978;
            end
          end
        end
      end
    end
    if (tlb__T_939) begin
      if (!(tlb__T_961)) begin
        if (!(tlb__T_979)) begin
          if (tlb__T_1135) begin
            if (2'h2 == tlb__T_1047) begin
              tlb_sectored_entries_5_data_2 <= tlb__T_978;
            end
          end
        end
      end
    end
    if (tlb__T_939) begin
      if (!(tlb__T_961)) begin
        if (!(tlb__T_979)) begin
          if (tlb__T_1135) begin
            if (2'h3 == tlb__T_1047) begin
              tlb_sectored_entries_5_data_3 <= tlb__T_978;
            end
          end
        end
      end
    end
    if (tlb__T_3753) begin
      tlb_sectored_entries_5_valid_0 <= 1'h0;
    end else if (tlb_io_sfence_valid) begin
      if (tlb_io_sfence_bits_rs1) begin
        if (tlb__T_3128) begin
          if (tlb__T_3131) begin
            tlb_sectored_entries_5_valid_0 <= 1'h0;
          end else if (tlb__T_445) begin
            if (2'h0 == tlb__T_510) begin
              tlb_sectored_entries_5_valid_0 <= 1'h0;
            end else if (tlb__T_939) begin
              if (!(tlb__T_961)) begin
                if (!(tlb__T_979)) begin
                  if (tlb__T_1135) begin
                    tlb_sectored_entries_5_valid_0 <= tlb__GEN_194;
                  end
                end
              end
            end
          end else if (tlb__T_939) begin
            if (!(tlb__T_961)) begin
              if (!(tlb__T_979)) begin
                if (tlb__T_1135) begin
                  tlb_sectored_entries_5_valid_0 <= tlb__GEN_194;
                end
              end
            end
          end
        end else if (tlb__T_445) begin
          if (2'h0 == tlb__T_510) begin
            tlb_sectored_entries_5_valid_0 <= 1'h0;
          end else if (tlb__T_939) begin
            if (!(tlb__T_961)) begin
              if (!(tlb__T_979)) begin
                if (tlb__T_1135) begin
                  tlb_sectored_entries_5_valid_0 <= tlb__GEN_194;
                end
              end
            end
          end
        end else if (tlb__T_939) begin
          if (!(tlb__T_961)) begin
            if (!(tlb__T_979)) begin
              if (tlb__T_1135) begin
                tlb_sectored_entries_5_valid_0 <= tlb__GEN_194;
              end
            end
          end
        end
      end else begin
        tlb_sectored_entries_5_valid_0 <= tlb__GEN_792;
      end
    end else begin
      tlb_sectored_entries_5_valid_0 <= tlb__GEN_522;
    end
    if (tlb__T_3753) begin
      tlb_sectored_entries_5_valid_1 <= 1'h0;
    end else if (tlb_io_sfence_valid) begin
      if (tlb_io_sfence_bits_rs1) begin
        if (tlb__T_3128) begin
          if (tlb__T_3149) begin
            tlb_sectored_entries_5_valid_1 <= 1'h0;
          end else if (tlb__T_445) begin
            if (2'h1 == tlb__T_510) begin
              tlb_sectored_entries_5_valid_1 <= 1'h0;
            end else if (tlb__T_939) begin
              if (!(tlb__T_961)) begin
                if (!(tlb__T_979)) begin
                  if (tlb__T_1135) begin
                    tlb_sectored_entries_5_valid_1 <= tlb__GEN_195;
                  end
                end
              end
            end
          end else if (tlb__T_939) begin
            if (!(tlb__T_961)) begin
              if (!(tlb__T_979)) begin
                if (tlb__T_1135) begin
                  tlb_sectored_entries_5_valid_1 <= tlb__GEN_195;
                end
              end
            end
          end
        end else if (tlb__T_445) begin
          if (2'h1 == tlb__T_510) begin
            tlb_sectored_entries_5_valid_1 <= 1'h0;
          end else if (tlb__T_939) begin
            if (!(tlb__T_961)) begin
              if (!(tlb__T_979)) begin
                if (tlb__T_1135) begin
                  tlb_sectored_entries_5_valid_1 <= tlb__GEN_195;
                end
              end
            end
          end
        end else if (tlb__T_939) begin
          if (!(tlb__T_961)) begin
            if (!(tlb__T_979)) begin
              if (tlb__T_1135) begin
                tlb_sectored_entries_5_valid_1 <= tlb__GEN_195;
              end
            end
          end
        end
      end else begin
        tlb_sectored_entries_5_valid_1 <= tlb__GEN_793;
      end
    end else begin
      tlb_sectored_entries_5_valid_1 <= tlb__GEN_523;
    end
    if (tlb__T_3753) begin
      tlb_sectored_entries_5_valid_2 <= 1'h0;
    end else if (tlb_io_sfence_valid) begin
      if (tlb_io_sfence_bits_rs1) begin
        if (tlb__T_3128) begin
          if (tlb__T_3167) begin
            tlb_sectored_entries_5_valid_2 <= 1'h0;
          end else if (tlb__T_445) begin
            if (2'h2 == tlb__T_510) begin
              tlb_sectored_entries_5_valid_2 <= 1'h0;
            end else if (tlb__T_939) begin
              if (!(tlb__T_961)) begin
                if (!(tlb__T_979)) begin
                  if (tlb__T_1135) begin
                    tlb_sectored_entries_5_valid_2 <= tlb__GEN_196;
                  end
                end
              end
            end
          end else if (tlb__T_939) begin
            if (!(tlb__T_961)) begin
              if (!(tlb__T_979)) begin
                if (tlb__T_1135) begin
                  tlb_sectored_entries_5_valid_2 <= tlb__GEN_196;
                end
              end
            end
          end
        end else if (tlb__T_445) begin
          if (2'h2 == tlb__T_510) begin
            tlb_sectored_entries_5_valid_2 <= 1'h0;
          end else if (tlb__T_939) begin
            if (!(tlb__T_961)) begin
              if (!(tlb__T_979)) begin
                if (tlb__T_1135) begin
                  tlb_sectored_entries_5_valid_2 <= tlb__GEN_196;
                end
              end
            end
          end
        end else if (tlb__T_939) begin
          if (!(tlb__T_961)) begin
            if (!(tlb__T_979)) begin
              if (tlb__T_1135) begin
                tlb_sectored_entries_5_valid_2 <= tlb__GEN_196;
              end
            end
          end
        end
      end else begin
        tlb_sectored_entries_5_valid_2 <= tlb__GEN_794;
      end
    end else begin
      tlb_sectored_entries_5_valid_2 <= tlb__GEN_524;
    end
    if (tlb__T_3753) begin
      tlb_sectored_entries_5_valid_3 <= 1'h0;
    end else if (tlb_io_sfence_valid) begin
      if (tlb_io_sfence_bits_rs1) begin
        if (tlb__T_3128) begin
          if (tlb__T_3185) begin
            tlb_sectored_entries_5_valid_3 <= 1'h0;
          end else if (tlb__T_445) begin
            if (2'h3 == tlb__T_510) begin
              tlb_sectored_entries_5_valid_3 <= 1'h0;
            end else if (tlb__T_939) begin
              if (!(tlb__T_961)) begin
                if (!(tlb__T_979)) begin
                  if (tlb__T_1135) begin
                    tlb_sectored_entries_5_valid_3 <= tlb__GEN_197;
                  end
                end
              end
            end
          end else if (tlb__T_939) begin
            if (!(tlb__T_961)) begin
              if (!(tlb__T_979)) begin
                if (tlb__T_1135) begin
                  tlb_sectored_entries_5_valid_3 <= tlb__GEN_197;
                end
              end
            end
          end
        end else if (tlb__T_445) begin
          if (2'h3 == tlb__T_510) begin
            tlb_sectored_entries_5_valid_3 <= 1'h0;
          end else if (tlb__T_939) begin
            if (!(tlb__T_961)) begin
              if (!(tlb__T_979)) begin
                if (tlb__T_1135) begin
                  tlb_sectored_entries_5_valid_3 <= tlb__GEN_197;
                end
              end
            end
          end
        end else if (tlb__T_939) begin
          if (!(tlb__T_961)) begin
            if (!(tlb__T_979)) begin
              if (tlb__T_1135) begin
                tlb_sectored_entries_5_valid_3 <= tlb__GEN_197;
              end
            end
          end
        end
      end else begin
        tlb_sectored_entries_5_valid_3 <= tlb__GEN_795;
      end
    end else begin
      tlb_sectored_entries_5_valid_3 <= tlb__GEN_525;
    end
    if (tlb__T_939) begin
      if (!(tlb__T_961)) begin
        if (!(tlb__T_979)) begin
          if (tlb__T_1153) begin
            tlb_sectored_entries_6_tag <= tlb_r_refill_tag;
          end
        end
      end
    end
    if (tlb__T_939) begin
      if (!(tlb__T_961)) begin
        if (!(tlb__T_979)) begin
          if (tlb__T_1153) begin
            if (2'h0 == tlb__T_1047) begin
              tlb_sectored_entries_6_data_0 <= tlb__T_978;
            end
          end
        end
      end
    end
    if (tlb__T_939) begin
      if (!(tlb__T_961)) begin
        if (!(tlb__T_979)) begin
          if (tlb__T_1153) begin
            if (2'h1 == tlb__T_1047) begin
              tlb_sectored_entries_6_data_1 <= tlb__T_978;
            end
          end
        end
      end
    end
    if (tlb__T_939) begin
      if (!(tlb__T_961)) begin
        if (!(tlb__T_979)) begin
          if (tlb__T_1153) begin
            if (2'h2 == tlb__T_1047) begin
              tlb_sectored_entries_6_data_2 <= tlb__T_978;
            end
          end
        end
      end
    end
    if (tlb__T_939) begin
      if (!(tlb__T_961)) begin
        if (!(tlb__T_979)) begin
          if (tlb__T_1153) begin
            if (2'h3 == tlb__T_1047) begin
              tlb_sectored_entries_6_data_3 <= tlb__T_978;
            end
          end
        end
      end
    end
    if (tlb__T_3753) begin
      tlb_sectored_entries_6_valid_0 <= 1'h0;
    end else if (tlb_io_sfence_valid) begin
      if (tlb_io_sfence_bits_rs1) begin
        if (tlb__T_3283) begin
          if (tlb__T_3286) begin
            tlb_sectored_entries_6_valid_0 <= 1'h0;
          end else if (tlb__T_451) begin
            if (2'h0 == tlb__T_510) begin
              tlb_sectored_entries_6_valid_0 <= 1'h0;
            end else if (tlb__T_939) begin
              if (!(tlb__T_961)) begin
                if (!(tlb__T_979)) begin
                  if (tlb__T_1153) begin
                    tlb_sectored_entries_6_valid_0 <= tlb__GEN_216;
                  end
                end
              end
            end
          end else if (tlb__T_939) begin
            if (!(tlb__T_961)) begin
              if (!(tlb__T_979)) begin
                if (tlb__T_1153) begin
                  tlb_sectored_entries_6_valid_0 <= tlb__GEN_216;
                end
              end
            end
          end
        end else if (tlb__T_451) begin
          if (2'h0 == tlb__T_510) begin
            tlb_sectored_entries_6_valid_0 <= 1'h0;
          end else if (tlb__T_939) begin
            if (!(tlb__T_961)) begin
              if (!(tlb__T_979)) begin
                if (tlb__T_1153) begin
                  tlb_sectored_entries_6_valid_0 <= tlb__GEN_216;
                end
              end
            end
          end
        end else if (tlb__T_939) begin
          if (!(tlb__T_961)) begin
            if (!(tlb__T_979)) begin
              if (tlb__T_1153) begin
                tlb_sectored_entries_6_valid_0 <= tlb__GEN_216;
              end
            end
          end
        end
      end else begin
        tlb_sectored_entries_6_valid_0 <= tlb__GEN_820;
      end
    end else begin
      tlb_sectored_entries_6_valid_0 <= tlb__GEN_532;
    end
    if (tlb__T_3753) begin
      tlb_sectored_entries_6_valid_1 <= 1'h0;
    end else if (tlb_io_sfence_valid) begin
      if (tlb_io_sfence_bits_rs1) begin
        if (tlb__T_3283) begin
          if (tlb__T_3304) begin
            tlb_sectored_entries_6_valid_1 <= 1'h0;
          end else if (tlb__T_451) begin
            if (2'h1 == tlb__T_510) begin
              tlb_sectored_entries_6_valid_1 <= 1'h0;
            end else if (tlb__T_939) begin
              if (!(tlb__T_961)) begin
                if (!(tlb__T_979)) begin
                  if (tlb__T_1153) begin
                    tlb_sectored_entries_6_valid_1 <= tlb__GEN_217;
                  end
                end
              end
            end
          end else if (tlb__T_939) begin
            if (!(tlb__T_961)) begin
              if (!(tlb__T_979)) begin
                if (tlb__T_1153) begin
                  tlb_sectored_entries_6_valid_1 <= tlb__GEN_217;
                end
              end
            end
          end
        end else if (tlb__T_451) begin
          if (2'h1 == tlb__T_510) begin
            tlb_sectored_entries_6_valid_1 <= 1'h0;
          end else if (tlb__T_939) begin
            if (!(tlb__T_961)) begin
              if (!(tlb__T_979)) begin
                if (tlb__T_1153) begin
                  tlb_sectored_entries_6_valid_1 <= tlb__GEN_217;
                end
              end
            end
          end
        end else if (tlb__T_939) begin
          if (!(tlb__T_961)) begin
            if (!(tlb__T_979)) begin
              if (tlb__T_1153) begin
                tlb_sectored_entries_6_valid_1 <= tlb__GEN_217;
              end
            end
          end
        end
      end else begin
        tlb_sectored_entries_6_valid_1 <= tlb__GEN_821;
      end
    end else begin
      tlb_sectored_entries_6_valid_1 <= tlb__GEN_533;
    end
    if (tlb__T_3753) begin
      tlb_sectored_entries_6_valid_2 <= 1'h0;
    end else if (tlb_io_sfence_valid) begin
      if (tlb_io_sfence_bits_rs1) begin
        if (tlb__T_3283) begin
          if (tlb__T_3322) begin
            tlb_sectored_entries_6_valid_2 <= 1'h0;
          end else if (tlb__T_451) begin
            if (2'h2 == tlb__T_510) begin
              tlb_sectored_entries_6_valid_2 <= 1'h0;
            end else if (tlb__T_939) begin
              if (!(tlb__T_961)) begin
                if (!(tlb__T_979)) begin
                  if (tlb__T_1153) begin
                    tlb_sectored_entries_6_valid_2 <= tlb__GEN_218;
                  end
                end
              end
            end
          end else if (tlb__T_939) begin
            if (!(tlb__T_961)) begin
              if (!(tlb__T_979)) begin
                if (tlb__T_1153) begin
                  tlb_sectored_entries_6_valid_2 <= tlb__GEN_218;
                end
              end
            end
          end
        end else if (tlb__T_451) begin
          if (2'h2 == tlb__T_510) begin
            tlb_sectored_entries_6_valid_2 <= 1'h0;
          end else if (tlb__T_939) begin
            if (!(tlb__T_961)) begin
              if (!(tlb__T_979)) begin
                if (tlb__T_1153) begin
                  tlb_sectored_entries_6_valid_2 <= tlb__GEN_218;
                end
              end
            end
          end
        end else if (tlb__T_939) begin
          if (!(tlb__T_961)) begin
            if (!(tlb__T_979)) begin
              if (tlb__T_1153) begin
                tlb_sectored_entries_6_valid_2 <= tlb__GEN_218;
              end
            end
          end
        end
      end else begin
        tlb_sectored_entries_6_valid_2 <= tlb__GEN_822;
      end
    end else begin
      tlb_sectored_entries_6_valid_2 <= tlb__GEN_534;
    end
    if (tlb__T_3753) begin
      tlb_sectored_entries_6_valid_3 <= 1'h0;
    end else if (tlb_io_sfence_valid) begin
      if (tlb_io_sfence_bits_rs1) begin
        if (tlb__T_3283) begin
          if (tlb__T_3340) begin
            tlb_sectored_entries_6_valid_3 <= 1'h0;
          end else if (tlb__T_451) begin
            if (2'h3 == tlb__T_510) begin
              tlb_sectored_entries_6_valid_3 <= 1'h0;
            end else if (tlb__T_939) begin
              if (!(tlb__T_961)) begin
                if (!(tlb__T_979)) begin
                  if (tlb__T_1153) begin
                    tlb_sectored_entries_6_valid_3 <= tlb__GEN_219;
                  end
                end
              end
            end
          end else if (tlb__T_939) begin
            if (!(tlb__T_961)) begin
              if (!(tlb__T_979)) begin
                if (tlb__T_1153) begin
                  tlb_sectored_entries_6_valid_3 <= tlb__GEN_219;
                end
              end
            end
          end
        end else if (tlb__T_451) begin
          if (2'h3 == tlb__T_510) begin
            tlb_sectored_entries_6_valid_3 <= 1'h0;
          end else if (tlb__T_939) begin
            if (!(tlb__T_961)) begin
              if (!(tlb__T_979)) begin
                if (tlb__T_1153) begin
                  tlb_sectored_entries_6_valid_3 <= tlb__GEN_219;
                end
              end
            end
          end
        end else if (tlb__T_939) begin
          if (!(tlb__T_961)) begin
            if (!(tlb__T_979)) begin
              if (tlb__T_1153) begin
                tlb_sectored_entries_6_valid_3 <= tlb__GEN_219;
              end
            end
          end
        end
      end else begin
        tlb_sectored_entries_6_valid_3 <= tlb__GEN_823;
      end
    end else begin
      tlb_sectored_entries_6_valid_3 <= tlb__GEN_535;
    end
    if (tlb__T_939) begin
      if (!(tlb__T_961)) begin
        if (!(tlb__T_979)) begin
          if (tlb__T_1171) begin
            tlb_sectored_entries_7_tag <= tlb_r_refill_tag;
          end
        end
      end
    end
    if (tlb__T_939) begin
      if (!(tlb__T_961)) begin
        if (!(tlb__T_979)) begin
          if (tlb__T_1171) begin
            if (2'h0 == tlb__T_1047) begin
              tlb_sectored_entries_7_data_0 <= tlb__T_978;
            end
          end
        end
      end
    end
    if (tlb__T_939) begin
      if (!(tlb__T_961)) begin
        if (!(tlb__T_979)) begin
          if (tlb__T_1171) begin
            if (2'h1 == tlb__T_1047) begin
              tlb_sectored_entries_7_data_1 <= tlb__T_978;
            end
          end
        end
      end
    end
    if (tlb__T_939) begin
      if (!(tlb__T_961)) begin
        if (!(tlb__T_979)) begin
          if (tlb__T_1171) begin
            if (2'h2 == tlb__T_1047) begin
              tlb_sectored_entries_7_data_2 <= tlb__T_978;
            end
          end
        end
      end
    end
    if (tlb__T_939) begin
      if (!(tlb__T_961)) begin
        if (!(tlb__T_979)) begin
          if (tlb__T_1171) begin
            if (2'h3 == tlb__T_1047) begin
              tlb_sectored_entries_7_data_3 <= tlb__T_978;
            end
          end
        end
      end
    end
    if (tlb__T_3753) begin
      tlb_sectored_entries_7_valid_0 <= 1'h0;
    end else if (tlb_io_sfence_valid) begin
      if (tlb_io_sfence_bits_rs1) begin
        if (tlb__T_3438) begin
          if (tlb__T_3441) begin
            tlb_sectored_entries_7_valid_0 <= 1'h0;
          end else if (tlb__T_457) begin
            if (2'h0 == tlb__T_510) begin
              tlb_sectored_entries_7_valid_0 <= 1'h0;
            end else if (tlb__T_939) begin
              if (!(tlb__T_961)) begin
                if (!(tlb__T_979)) begin
                  if (tlb__T_1171) begin
                    tlb_sectored_entries_7_valid_0 <= tlb__GEN_238;
                  end
                end
              end
            end
          end else if (tlb__T_939) begin
            if (!(tlb__T_961)) begin
              if (!(tlb__T_979)) begin
                if (tlb__T_1171) begin
                  tlb_sectored_entries_7_valid_0 <= tlb__GEN_238;
                end
              end
            end
          end
        end else if (tlb__T_457) begin
          if (2'h0 == tlb__T_510) begin
            tlb_sectored_entries_7_valid_0 <= 1'h0;
          end else if (tlb__T_939) begin
            if (!(tlb__T_961)) begin
              if (!(tlb__T_979)) begin
                if (tlb__T_1171) begin
                  tlb_sectored_entries_7_valid_0 <= tlb__GEN_238;
                end
              end
            end
          end
        end else if (tlb__T_939) begin
          if (!(tlb__T_961)) begin
            if (!(tlb__T_979)) begin
              if (tlb__T_1171) begin
                tlb_sectored_entries_7_valid_0 <= tlb__GEN_238;
              end
            end
          end
        end
      end else begin
        tlb_sectored_entries_7_valid_0 <= tlb__GEN_848;
      end
    end else begin
      tlb_sectored_entries_7_valid_0 <= tlb__GEN_542;
    end
    if (tlb__T_3753) begin
      tlb_sectored_entries_7_valid_1 <= 1'h0;
    end else if (tlb_io_sfence_valid) begin
      if (tlb_io_sfence_bits_rs1) begin
        if (tlb__T_3438) begin
          if (tlb__T_3459) begin
            tlb_sectored_entries_7_valid_1 <= 1'h0;
          end else if (tlb__T_457) begin
            if (2'h1 == tlb__T_510) begin
              tlb_sectored_entries_7_valid_1 <= 1'h0;
            end else if (tlb__T_939) begin
              if (!(tlb__T_961)) begin
                if (!(tlb__T_979)) begin
                  if (tlb__T_1171) begin
                    tlb_sectored_entries_7_valid_1 <= tlb__GEN_239;
                  end
                end
              end
            end
          end else if (tlb__T_939) begin
            if (!(tlb__T_961)) begin
              if (!(tlb__T_979)) begin
                if (tlb__T_1171) begin
                  tlb_sectored_entries_7_valid_1 <= tlb__GEN_239;
                end
              end
            end
          end
        end else if (tlb__T_457) begin
          if (2'h1 == tlb__T_510) begin
            tlb_sectored_entries_7_valid_1 <= 1'h0;
          end else if (tlb__T_939) begin
            if (!(tlb__T_961)) begin
              if (!(tlb__T_979)) begin
                if (tlb__T_1171) begin
                  tlb_sectored_entries_7_valid_1 <= tlb__GEN_239;
                end
              end
            end
          end
        end else if (tlb__T_939) begin
          if (!(tlb__T_961)) begin
            if (!(tlb__T_979)) begin
              if (tlb__T_1171) begin
                tlb_sectored_entries_7_valid_1 <= tlb__GEN_239;
              end
            end
          end
        end
      end else begin
        tlb_sectored_entries_7_valid_1 <= tlb__GEN_849;
      end
    end else begin
      tlb_sectored_entries_7_valid_1 <= tlb__GEN_543;
    end
    if (tlb__T_3753) begin
      tlb_sectored_entries_7_valid_2 <= 1'h0;
    end else if (tlb_io_sfence_valid) begin
      if (tlb_io_sfence_bits_rs1) begin
        if (tlb__T_3438) begin
          if (tlb__T_3477) begin
            tlb_sectored_entries_7_valid_2 <= 1'h0;
          end else if (tlb__T_457) begin
            if (2'h2 == tlb__T_510) begin
              tlb_sectored_entries_7_valid_2 <= 1'h0;
            end else if (tlb__T_939) begin
              if (!(tlb__T_961)) begin
                if (!(tlb__T_979)) begin
                  if (tlb__T_1171) begin
                    tlb_sectored_entries_7_valid_2 <= tlb__GEN_240;
                  end
                end
              end
            end
          end else if (tlb__T_939) begin
            if (!(tlb__T_961)) begin
              if (!(tlb__T_979)) begin
                if (tlb__T_1171) begin
                  tlb_sectored_entries_7_valid_2 <= tlb__GEN_240;
                end
              end
            end
          end
        end else if (tlb__T_457) begin
          if (2'h2 == tlb__T_510) begin
            tlb_sectored_entries_7_valid_2 <= 1'h0;
          end else if (tlb__T_939) begin
            if (!(tlb__T_961)) begin
              if (!(tlb__T_979)) begin
                if (tlb__T_1171) begin
                  tlb_sectored_entries_7_valid_2 <= tlb__GEN_240;
                end
              end
            end
          end
        end else if (tlb__T_939) begin
          if (!(tlb__T_961)) begin
            if (!(tlb__T_979)) begin
              if (tlb__T_1171) begin
                tlb_sectored_entries_7_valid_2 <= tlb__GEN_240;
              end
            end
          end
        end
      end else begin
        tlb_sectored_entries_7_valid_2 <= tlb__GEN_850;
      end
    end else begin
      tlb_sectored_entries_7_valid_2 <= tlb__GEN_544;
    end
    if (tlb__T_3753) begin
      tlb_sectored_entries_7_valid_3 <= 1'h0;
    end else if (tlb_io_sfence_valid) begin
      if (tlb_io_sfence_bits_rs1) begin
        if (tlb__T_3438) begin
          if (tlb__T_3495) begin
            tlb_sectored_entries_7_valid_3 <= 1'h0;
          end else if (tlb__T_457) begin
            if (2'h3 == tlb__T_510) begin
              tlb_sectored_entries_7_valid_3 <= 1'h0;
            end else if (tlb__T_939) begin
              if (!(tlb__T_961)) begin
                if (!(tlb__T_979)) begin
                  if (tlb__T_1171) begin
                    tlb_sectored_entries_7_valid_3 <= tlb__GEN_241;
                  end
                end
              end
            end
          end else if (tlb__T_939) begin
            if (!(tlb__T_961)) begin
              if (!(tlb__T_979)) begin
                if (tlb__T_1171) begin
                  tlb_sectored_entries_7_valid_3 <= tlb__GEN_241;
                end
              end
            end
          end
        end else if (tlb__T_457) begin
          if (2'h3 == tlb__T_510) begin
            tlb_sectored_entries_7_valid_3 <= 1'h0;
          end else if (tlb__T_939) begin
            if (!(tlb__T_961)) begin
              if (!(tlb__T_979)) begin
                if (tlb__T_1171) begin
                  tlb_sectored_entries_7_valid_3 <= tlb__GEN_241;
                end
              end
            end
          end
        end else if (tlb__T_939) begin
          if (!(tlb__T_961)) begin
            if (!(tlb__T_979)) begin
              if (tlb__T_1171) begin
                tlb_sectored_entries_7_valid_3 <= tlb__GEN_241;
              end
            end
          end
        end
      end else begin
        tlb_sectored_entries_7_valid_3 <= tlb__GEN_851;
      end
    end else begin
      tlb_sectored_entries_7_valid_3 <= tlb__GEN_545;
    end
    if (tlb__T_939) begin
      if (!(tlb__T_961)) begin
        if (tlb__T_979) begin
          if (tlb__T_980) begin
            tlb_superpage_entries_0_tag <= tlb_r_refill_tag;
          end
        end
      end
    end
    if (tlb__T_939) begin
      if (!(tlb__T_961)) begin
        if (tlb__T_979) begin
          if (tlb__T_980) begin
            tlb_superpage_entries_0_data_0 <= tlb__T_978;
          end
        end
      end
    end
    if (tlb__T_3753) begin
      tlb_superpage_entries_0_valid_0 <= 1'h0;
    end else if (tlb_io_sfence_valid) begin
      if (tlb_io_sfence_bits_rs1) begin
        if (tlb__T_464) begin
          tlb_superpage_entries_0_valid_0 <= 1'h0;
        end else if (tlb__T_939) begin
          if (!(tlb__T_961)) begin
            if (tlb__T_979) begin
              tlb_superpage_entries_0_valid_0 <= tlb__GEN_66;
            end
          end
        end
      end else begin
        tlb_superpage_entries_0_valid_0 <= tlb__GEN_858;
      end
    end else if (tlb__T_939) begin
      if (!(tlb__T_961)) begin
        if (tlb__T_979) begin
          tlb_superpage_entries_0_valid_0 <= tlb__GEN_66;
        end
      end
    end
    if (tlb__T_939) begin
      if (!(tlb__T_961)) begin
        if (tlb__T_979) begin
          if (tlb__T_996) begin
            tlb_superpage_entries_1_tag <= tlb_r_refill_tag;
          end
        end
      end
    end
    if (tlb__T_939) begin
      if (!(tlb__T_961)) begin
        if (tlb__T_979) begin
          if (tlb__T_996) begin
            tlb_superpage_entries_1_data_0 <= tlb__T_978;
          end
        end
      end
    end
    if (tlb__T_3753) begin
      tlb_superpage_entries_1_valid_0 <= 1'h0;
    end else if (tlb_io_sfence_valid) begin
      if (tlb_io_sfence_bits_rs1) begin
        if (tlb__T_477) begin
          tlb_superpage_entries_1_valid_0 <= 1'h0;
        end else if (tlb__T_939) begin
          if (!(tlb__T_961)) begin
            if (tlb__T_979) begin
              tlb_superpage_entries_1_valid_0 <= tlb__GEN_70;
            end
          end
        end
      end else begin
        tlb_superpage_entries_1_valid_0 <= tlb__GEN_862;
      end
    end else if (tlb__T_939) begin
      if (!(tlb__T_961)) begin
        if (tlb__T_979) begin
          tlb_superpage_entries_1_valid_0 <= tlb__GEN_70;
        end
      end
    end
    if (tlb__T_939) begin
      if (!(tlb__T_961)) begin
        if (tlb__T_979) begin
          if (tlb__T_1012) begin
            tlb_superpage_entries_2_tag <= tlb_r_refill_tag;
          end
        end
      end
    end
    if (tlb__T_939) begin
      if (!(tlb__T_961)) begin
        if (tlb__T_979) begin
          if (tlb__T_1012) begin
            tlb_superpage_entries_2_data_0 <= tlb__T_978;
          end
        end
      end
    end
    if (tlb__T_3753) begin
      tlb_superpage_entries_2_valid_0 <= 1'h0;
    end else if (tlb_io_sfence_valid) begin
      if (tlb_io_sfence_bits_rs1) begin
        if (tlb__T_490) begin
          tlb_superpage_entries_2_valid_0 <= 1'h0;
        end else if (tlb__T_939) begin
          if (!(tlb__T_961)) begin
            if (tlb__T_979) begin
              tlb_superpage_entries_2_valid_0 <= tlb__GEN_74;
            end
          end
        end
      end else begin
        tlb_superpage_entries_2_valid_0 <= tlb__GEN_866;
      end
    end else if (tlb__T_939) begin
      if (!(tlb__T_961)) begin
        if (tlb__T_979) begin
          tlb_superpage_entries_2_valid_0 <= tlb__GEN_74;
        end
      end
    end
    if (tlb__T_939) begin
      if (!(tlb__T_961)) begin
        if (tlb__T_979) begin
          if (tlb__T_1028) begin
            tlb_superpage_entries_3_tag <= tlb_r_refill_tag;
          end
        end
      end
    end
    if (tlb__T_939) begin
      if (!(tlb__T_961)) begin
        if (tlb__T_979) begin
          if (tlb__T_1028) begin
            tlb_superpage_entries_3_data_0 <= tlb__T_978;
          end
        end
      end
    end
    if (tlb__T_3753) begin
      tlb_superpage_entries_3_valid_0 <= 1'h0;
    end else if (tlb_io_sfence_valid) begin
      if (tlb_io_sfence_bits_rs1) begin
        if (tlb__T_503) begin
          tlb_superpage_entries_3_valid_0 <= 1'h0;
        end else if (tlb__T_939) begin
          if (!(tlb__T_961)) begin
            if (tlb__T_979) begin
              tlb_superpage_entries_3_valid_0 <= tlb__GEN_78;
            end
          end
        end
      end else begin
        tlb_superpage_entries_3_valid_0 <= tlb__GEN_870;
      end
    end else if (tlb__T_939) begin
      if (!(tlb__T_961)) begin
        if (tlb__T_979) begin
          tlb_superpage_entries_3_valid_0 <= tlb__GEN_78;
        end
      end
    end
    if (tlb__T_939) begin
      if (tlb__T_961) begin
        tlb_special_entry_level <= tlb_io_ptw_resp_bits_level;
      end
    end
    if (tlb__T_939) begin
      if (tlb__T_961) begin
        tlb_special_entry_tag <= tlb_r_refill_tag;
      end
    end
    if (tlb__T_939) begin
      if (tlb__T_961) begin
        tlb_special_entry_data_0 <= tlb__T_978;
      end
    end
    if (tlb__T_3753) begin
      tlb_special_entry_valid_0 <= 1'h0;
    end else if (tlb_io_sfence_valid) begin
      if (tlb_io_sfence_bits_rs1) begin
        if (tlb__T_619) begin
          tlb_special_entry_valid_0 <= 1'h0;
        end else if (tlb__T_939) begin
          tlb_special_entry_valid_0 <= tlb__GEN_354;
        end
      end else begin
        tlb_special_entry_valid_0 <= tlb__GEN_874;
      end
    end else if (tlb__T_939) begin
      tlb_special_entry_valid_0 <= tlb__GEN_354;
    end
    if (tlb_reset) begin
      tlb_state <= 2'h0;
    end else if (tlb_io_ptw_resp_valid) begin
      tlb_state <= 2'h0;
    end else if (tlb__T_2339) begin
      tlb_state <= 2'h3;
    end else if (tlb__T_4) begin
      if (tlb_io_ptw_req_ready) begin
        if (tlb_io_sfence_valid) begin
          tlb_state <= 2'h3;
        end else begin
          tlb_state <= 2'h2;
        end
      end else if (tlb_io_sfence_valid) begin
        tlb_state <= 2'h0;
      end else if (tlb__T_2222) begin
        tlb_state <= 2'h1;
      end
    end else if (tlb__T_2222) begin
      tlb_state <= 2'h1;
    end
    if (tlb__T_2222) begin
      tlb_r_refill_tag <= tlb_vpn;
    end
    if (tlb__T_2222) begin
      if (tlb__T_2233) begin
        tlb_r_superpage_repl_addr <= tlb__T_2229;
      end else if (tlb__T_2235) begin
        tlb_r_superpage_repl_addr <= 2'h0;
      end else if (tlb__T_2236) begin
        tlb_r_superpage_repl_addr <= 2'h1;
      end else if (tlb__T_2237) begin
        tlb_r_superpage_repl_addr <= 2'h2;
      end else begin
        tlb_r_superpage_repl_addr <= 2'h3;
      end
    end
    if (tlb__T_2222) begin
      if (tlb__T_2293) begin
        tlb_r_sectored_repl_addr <= tlb__T_2261;
      end else if (tlb__T_2295) begin
        tlb_r_sectored_repl_addr <= 3'h0;
      end else if (tlb__T_2296) begin
        tlb_r_sectored_repl_addr <= 3'h1;
      end else if (tlb__T_2297) begin
        tlb_r_sectored_repl_addr <= 3'h2;
      end else if (tlb__T_2298) begin
        tlb_r_sectored_repl_addr <= 3'h3;
      end else if (tlb__T_2299) begin
        tlb_r_sectored_repl_addr <= 3'h4;
      end else if (tlb__T_2300) begin
        tlb_r_sectored_repl_addr <= 3'h5;
      end else if (tlb__T_2301) begin
        tlb_r_sectored_repl_addr <= 3'h6;
      end else begin
        tlb_r_sectored_repl_addr <= 3'h7;
      end
    end
    if (tlb__T_2222) begin
      tlb_r_sectored_hit_addr <= tlb__T_2034;
    end
    if (tlb__T_2222) begin
      tlb_r_sectored_hit <= tlb__T_2016;
    end
    if (tlb__T_2009) begin
      if (tlb__T_2016) begin
        tlb__T_2007 <= tlb__T_2073;
      end
    end
    if (tlb__T_2009) begin
      if (tlb__T_2076) begin
        tlb__T_2008 <= tlb__T_2100;
      end
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (tlb_io_sfence_valid & tlb__T_2346) begin
          $fwrite(32'h80000002,"Assertion failed\n    at TLB.scala:376 assert(!io.sfence.bits.rs1 || (io.sfence.bits.addr >> pgIdxBits) === vpn)\n"); // @[TLB.scala 376:13:freechips.rocketchip.system.DefaultRV32Config.fir@180461.8]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (tlb_io_sfence_valid & tlb__T_2346) begin
          $fatal; // @[TLB.scala 376:13:freechips.rocketchip.system.DefaultRV32Config.fir@180462.8]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
  end
  always @(posedge gated_clock) begin
    if (reset) begin
      s1_valid <= 1'h0;
    end else begin
      s1_valid <= _T_16;
    end
    if (reset) begin
      blockProbeAfterGrantCount <= 3'h0;
    end else if (_T_2217) begin
      if (grantIsCached) begin
        if (d_last) begin
          blockProbeAfterGrantCount <= 3'h7;
        end else if (_T_2338) begin
          blockProbeAfterGrantCount <= _T_2205;
        end
      end else if (_T_2338) begin
        blockProbeAfterGrantCount <= _T_2205;
      end
    end else if (_T_2338) begin
      blockProbeAfterGrantCount <= _T_2205;
    end
    if (reset) begin
      lrscCount <= 7'h0;
    end else if (s1_probe) begin
      lrscCount <= 7'h0;
    end else if (_T_839) begin
      lrscCount <= 7'h3;
    end else if (_T_823) begin
      lrscCount <= _T_838;
    end else if (_T_831) begin
      if (s2_hit) begin
        lrscCount <= 7'h4f;
      end else begin
        lrscCount <= 7'h0;
      end
    end
    if (reset) begin
      s1_probe <= 1'h0;
    end else if (_T_2403) begin
      s1_probe <= _GEN_290;
    end else begin
      s1_probe <= _T_17;
    end
    if (reset) begin
      s2_probe <= 1'h0;
    end else begin
      s2_probe <= s1_probe;
    end
    if (reset) begin
      release_state <= 3'h0;
    end else if (_T_2455) begin
      release_state <= 3'h0;
    end else if (_T_2412) begin
      if (releaseDone) begin
        release_state <= 3'h6;
      end else if (_T_2409) begin
        if (releaseDone) begin
          release_state <= 3'h7;
        end else if (_T_2408) begin
          if (releaseDone) begin
            release_state <= 3'h7;
          end else if (_T_2407) begin
            if (releaseDone) begin
              release_state <= 3'h0;
            end else if (_T_2403) begin
              if (metaArb_io_in_6_ready) begin
                release_state <= 3'h0;
              end else if (s2_probe) begin
                if (pma_checker__T_2026) begin
                  release_state <= 3'h4;
                end else if (s2_prb_ack_data) begin
                  release_state <= 3'h2;
                end else if (_T_2399) begin
                  if (releaseDone) begin
                    release_state <= 3'h7;
                  end else begin
                    release_state <= 3'h3;
                  end
                end else if (releaseDone) begin
                  release_state <= 3'h0;
                end else begin
                  release_state <= 3'h5;
                end
              end else if (s2_want_victimize) begin
                if (_T_2394) begin
                  release_state <= 3'h1;
                end else begin
                  release_state <= 3'h6;
                end
              end
            end else if (s2_probe) begin
              if (pma_checker__T_2026) begin
                release_state <= 3'h4;
              end else if (s2_prb_ack_data) begin
                release_state <= 3'h2;
              end else if (_T_2399) begin
                if (releaseDone) begin
                  release_state <= 3'h7;
                end else begin
                  release_state <= 3'h3;
                end
              end else if (releaseDone) begin
                release_state <= 3'h0;
              end else begin
                release_state <= 3'h5;
              end
            end else if (s2_want_victimize) begin
              if (_T_2394) begin
                release_state <= 3'h1;
              end else begin
                release_state <= 3'h6;
              end
            end
          end else if (_T_2403) begin
            if (metaArb_io_in_6_ready) begin
              release_state <= 3'h0;
            end else if (s2_probe) begin
              if (pma_checker__T_2026) begin
                release_state <= 3'h4;
              end else if (s2_prb_ack_data) begin
                release_state <= 3'h2;
              end else if (_T_2399) begin
                if (releaseDone) begin
                  release_state <= 3'h7;
                end else begin
                  release_state <= 3'h3;
                end
              end else if (releaseDone) begin
                release_state <= 3'h0;
              end else begin
                release_state <= 3'h5;
              end
            end else if (s2_want_victimize) begin
              if (_T_2394) begin
                release_state <= 3'h1;
              end else begin
                release_state <= 3'h6;
              end
            end
          end else if (s2_probe) begin
            if (pma_checker__T_2026) begin
              release_state <= 3'h4;
            end else if (s2_prb_ack_data) begin
              release_state <= 3'h2;
            end else if (_T_2399) begin
              if (releaseDone) begin
                release_state <= 3'h7;
              end else begin
                release_state <= 3'h3;
              end
            end else if (releaseDone) begin
              release_state <= 3'h0;
            end else begin
              release_state <= 3'h5;
            end
          end else if (s2_want_victimize) begin
            if (_T_2394) begin
              release_state <= 3'h1;
            end else begin
              release_state <= 3'h6;
            end
          end
        end else if (_T_2407) begin
          if (releaseDone) begin
            release_state <= 3'h0;
          end else if (_T_2403) begin
            if (metaArb_io_in_6_ready) begin
              release_state <= 3'h0;
            end else begin
              release_state <= _GEN_279;
            end
          end else begin
            release_state <= _GEN_279;
          end
        end else if (_T_2403) begin
          if (metaArb_io_in_6_ready) begin
            release_state <= 3'h0;
          end else begin
            release_state <= _GEN_279;
          end
        end else begin
          release_state <= _GEN_279;
        end
      end else if (_T_2408) begin
        if (releaseDone) begin
          release_state <= 3'h7;
        end else if (_T_2407) begin
          if (releaseDone) begin
            release_state <= 3'h0;
          end else begin
            release_state <= _GEN_294;
          end
        end else begin
          release_state <= _GEN_294;
        end
      end else if (_T_2407) begin
        if (releaseDone) begin
          release_state <= 3'h0;
        end else begin
          release_state <= _GEN_294;
        end
      end else begin
        release_state <= _GEN_294;
      end
    end else if (_T_2409) begin
      if (releaseDone) begin
        release_state <= 3'h7;
      end else if (_T_2408) begin
        if (releaseDone) begin
          release_state <= 3'h7;
        end else begin
          release_state <= _GEN_298;
        end
      end else begin
        release_state <= _GEN_298;
      end
    end else if (_T_2408) begin
      if (releaseDone) begin
        release_state <= 3'h7;
      end else begin
        release_state <= _GEN_298;
      end
    end else begin
      release_state <= _GEN_298;
    end
    if (reset) begin
      release_ack_wait <= 1'h0;
    end else if (_T_2412) begin
      release_ack_wait <= _GEN_319;
    end else if (_T_2217) begin
      if (!(grantIsCached)) begin
        if (!(grantIsUncached)) begin
          if (grantIsVoluntary) begin
            release_ack_wait <= 1'h0;
          end
        end
      end
    end
    if (_T_2412) begin
      if (_T_2434) begin
        release_ack_addr <= probe_bits_address;
      end
    end
    if (reset) begin
      grantInProgress <= 1'h0;
    end else if (_T_2217) begin
      if (grantIsCached) begin
        if (d_last) begin
          grantInProgress <= 1'h0;
        end else begin
          grantInProgress <= 1'h1;
        end
      end
    end
    if (reset) begin
      s2_valid <= 1'h0;
    end else begin
      s2_valid <= _T_357;
    end
    if (s2_want_victimize) begin
      probe_bits_param <= 2'h0;
    end else if (_T_17) begin
      probe_bits_param <= auto_out_b_bits_param;
    end
    if (s2_want_victimize) begin
      probe_bits_size <= 4'h0;
    end else if (_T_17) begin
      probe_bits_size <= auto_out_b_bits_size;
    end
    if (s2_want_victimize) begin
      probe_bits_source <= 1'h0;
    end else if (_T_17) begin
      probe_bits_source <= auto_out_b_bits_source;
    end
    if (s2_want_victimize) begin
      probe_bits_address <= res_2_address;
    end else if (_T_17) begin
      probe_bits_address <= auto_out_b_bits_address;
    end
    if (s1_probe) begin
      s2_probe_state_state <= s1_meta_hit_state_state;
    end
    if (reset) begin
      _T_2362 <= 10'h0;
    end else if (_T_2354) begin
      if (c_first) begin
        if (tl_out__c_bits_opcode[0]) begin
          _T_2362 <= _T_2358[11:2];
        end else begin
          _T_2362 <= 10'h0;
        end
      end else begin
        _T_2362 <= _T_2364;
      end
    end
    s2_release_data_valid <= s1_release_data_valid & _T_2370;
    if (s0_clk_en) begin
      s1_req_cmd <= io_cpu_req_bits_cmd;
    end
    if (_T_2217) begin
      if (grantIsCached) begin
        if (s1_valid_not_nacked) begin
          s2_req_cmd <= s1_req_cmd;
        end
      end else if (grantIsUncached) begin
        if (grantIsUncachedData) begin
          s2_req_cmd <= 5'h0;
        end else if (s1_valid_not_nacked) begin
          s2_req_cmd <= s1_req_cmd;
        end
      end else if (s1_valid_not_nacked) begin
        s2_req_cmd <= s1_req_cmd;
      end
    end else if (s1_valid_not_nacked) begin
      s2_req_cmd <= s1_req_cmd;
    end
    pstore1_held <= _T_1018 & _T_1019;
    if (_T_847) begin
      pstore1_addr <= s1_req_addr;
    end
    if (s0_clk_en) begin
      s1_req_addr <= s0_req_addr;
    end
    if (_T_847) begin
      if (_T_53) begin
        pstore1_mask <= io_cpu_s1_data_mask;
      end else begin
        pstore1_mask <= s1_mask_xwr;
      end
    end
    if (s0_clk_en) begin
      s1_req_size <= io_cpu_req_bits_size;
    end
    pstore2_valid <= _T_1024 | advance_pstore1;
    if (advance_pstore1) begin
      pstore2_addr <= pstore1_addr;
    end
    if (advance_pstore1) begin
      mask <= _T_1054;
    end
    s2_not_nacked_in_s1 <= ~s1_nack;
    if (s1_valid_not_nacked) begin
      s2_hit_state_state <= s1_meta_hit_state_state;
    end
    if (s0_clk_en) begin
      s1_req_tag <= io_cpu_req_bits_tag;
    end
    if (s0_clk_en) begin
      s1_req_signed <= io_cpu_req_bits_signed;
    end
    if (s0_clk_en) begin
      s1_req_dprv <= io_cpu_req_bits_dprv;
    end
    if (s0_clk_en) begin
      s1_tlb_req_vaddr <= s0_req_addr;
    end
    if (s0_clk_en) begin
      s1_tlb_req_passthrough <= s0_req_phys;
    end
    if (s0_clk_en) begin
      s1_tlb_req_size <= io_cpu_req_bits_size;
    end
    if (s0_clk_en) begin
      s1_tlb_req_cmd <= io_cpu_req_bits_cmd;
    end
    if (reset) begin
      cached_grant_wait <= 1'h0;
    end else if (_T_2217) begin
      if (grantIsCached) begin
        if (d_last) begin
          cached_grant_wait <= 1'h0;
        end else if (_T_2164) begin
          if (!(s2_uncached)) begin
            cached_grant_wait <= 1'h1;
          end
        end
      end else if (_T_2164) begin
        if (!(s2_uncached)) begin
          cached_grant_wait <= 1'h1;
        end
      end
    end else if (_T_2164) begin
      if (!(s2_uncached)) begin
        cached_grant_wait <= 1'h1;
      end
    end
    if (reset) begin
      uncachedInFlight_0 <= 1'h0;
    end else if (_T_2217) begin
      if (grantIsCached) begin
        if (_T_2164) begin
          if (s2_uncached) begin
            uncachedInFlight_0 <= _GEN_139;
          end
        end
      end else if (grantIsUncached) begin
        if (_T_2222) begin
          uncachedInFlight_0 <= 1'h0;
        end else if (_T_2164) begin
          if (s2_uncached) begin
            uncachedInFlight_0 <= _GEN_139;
          end
        end
      end else if (_T_2164) begin
        if (s2_uncached) begin
          uncachedInFlight_0 <= _GEN_139;
        end
      end
    end else if (_T_2164) begin
      if (s2_uncached) begin
        uncachedInFlight_0 <= _GEN_139;
      end
    end
    if (_T_2164) begin
      if (s2_uncached) begin
        if (a_sel) begin
          uncachedReqs_0_addr <= s2_req_addr;
        end
      end
    end
    if (_T_2164) begin
      if (s2_uncached) begin
        if (a_sel) begin
          uncachedReqs_0_tag <= s2_req_tag;
        end
      end
    end
    if (_T_2164) begin
      if (s2_uncached) begin
        if (a_sel) begin
          uncachedReqs_0_size <= s2_req_size;
        end
      end
    end
    if (_T_2164) begin
      if (s2_uncached) begin
        if (a_sel) begin
          uncachedReqs_0_signed <= s2_req_signed;
        end
      end
    end
    if (s0_clk_en) begin
      s1_did_read <= _T_224;
    end
    if (s1_valid_not_nacked) begin
      s2_hit_way <= s1_meta_hit_way;
    end
    if (s1_valid_not_nacked) begin
      _T_632 <= s1_victim_way;
    end
    if (s1_probe) begin
      s2_probe_way <= s1_meta_hit_way;
    end
    if (_T_2217) begin
      if (grantIsCached) begin
        if (s1_valid_not_nacked) begin
          s2_req_addr <= s1_paddr;
        end
      end else if (grantIsUncached) begin
        if (grantIsUncachedData) begin
          s2_req_addr <= _T_2229;
        end else if (s1_valid_not_nacked) begin
          s2_req_addr <= s1_paddr;
        end
      end else if (s1_valid_not_nacked) begin
        s2_req_addr <= s1_paddr;
      end
    end else if (s1_valid_not_nacked) begin
      s2_req_addr <= s1_paddr;
    end
    if (_T_2217) begin
      if (grantIsCached) begin
        if (s1_valid_not_nacked) begin
          s2_req_tag <= s1_req_tag;
        end
      end else if (grantIsUncached) begin
        if (grantIsUncachedData) begin
          s2_req_tag <= uncachedReqs_0_tag;
        end else if (s1_valid_not_nacked) begin
          s2_req_tag <= s1_req_tag;
        end
      end else if (s1_valid_not_nacked) begin
        s2_req_tag <= s1_req_tag;
      end
    end else if (s1_valid_not_nacked) begin
      s2_req_tag <= s1_req_tag;
    end
    if (_T_2217) begin
      if (grantIsCached) begin
        if (s1_valid_not_nacked) begin
          s2_req_size <= s1_req_size;
        end
      end else if (grantIsUncached) begin
        if (grantIsUncachedData) begin
          s2_req_size <= uncachedReqs_0_size;
        end else if (s1_valid_not_nacked) begin
          s2_req_size <= s1_req_size;
        end
      end else if (s1_valid_not_nacked) begin
        s2_req_size <= s1_req_size;
      end
    end else if (s1_valid_not_nacked) begin
      s2_req_size <= s1_req_size;
    end
    if (_T_2217) begin
      if (grantIsCached) begin
        if (s1_valid_not_nacked) begin
          s2_req_signed <= s1_req_signed;
        end
      end else if (grantIsUncached) begin
        if (grantIsUncachedData) begin
          s2_req_signed <= uncachedReqs_0_signed;
        end else if (s1_valid_not_nacked) begin
          s2_req_signed <= s1_req_signed;
        end
      end else if (s1_valid_not_nacked) begin
        s2_req_signed <= s1_req_signed;
      end
    end else if (s1_valid_not_nacked) begin
      s2_req_signed <= s1_req_signed;
    end
    if (s1_valid_not_nacked) begin
      s2_req_dprv <= s1_req_dprv;
    end
    if (s1_valid_not_nacked) begin
      s2_tlb_xcpt_pf_ld <= tlb_io_resp_pf_ld;
    end
    if (s1_valid_not_nacked) begin
      s2_tlb_xcpt_pf_st <= tlb_io_resp_pf_st;
    end
    if (s1_valid_not_nacked) begin
      s2_tlb_xcpt_ae_ld <= tlb_io_resp_ae_ld;
    end
    if (s1_valid_not_nacked) begin
      s2_tlb_xcpt_ae_st <= tlb_io_resp_ae_st;
    end
    if (s1_valid_not_nacked) begin
      s2_tlb_xcpt_ma_ld <= tlb_io_resp_ma_ld;
    end
    if (s1_valid_not_nacked) begin
      s2_tlb_xcpt_ma_st <= tlb_io_resp_ma_st;
    end
    if (s1_valid_not_nacked) begin
      s2_pma_cacheable <= tlb_io_resp_cacheable;
    end
    if (_T_2217) begin
      if (!(grantIsCached)) begin
        if (grantIsUncached) begin
          if (grantIsUncachedData) begin
            s2_uncached_resp_addr <= uncachedReqs_0_addr;
          end
        end
      end
    end
    if (s1_valid_not_nacked) begin
      _T_377 <= s1_req_addr;
    end
    if (s1_meta_clk_en) begin
      _T_449 <= tag_array_RW0_rdata_3;
    end
    if (_T_2334) begin
      if (auto_out_d_valid) begin
        blockUncachedGrant <= _T_2247;
      end else begin
        blockUncachedGrant <= dataArb_io_out_valid;
      end
    end else begin
      blockUncachedGrant <= dataArb_io_out_valid;
    end
    if (reset) begin
      _T_2177 <= 10'h0;
    end else if (_T_2217) begin
      if (d_first) begin
        if (auto_out_d_bits_opcode[0]) begin
          _T_2177 <= _T_2173[11:2];
        end else begin
          _T_2177 <= 10'h0;
        end
      end else begin
        _T_2177 <= _T_2179;
      end
    end
    if (en) begin
      s2_data <= _T_474;
    end
    if (s1_valid_not_nacked) begin
      if (_T_320) begin
        _T_637 <= s1_meta_uncorrected_3_tag;
      end else if (_T_318) begin
        _T_637 <= s1_meta_uncorrected_2_tag;
      end else if (_T_316) begin
        _T_637 <= s1_meta_uncorrected_1_tag;
      end else begin
        _T_637 <= s1_meta_uncorrected_0_tag;
      end
    end
    if (s1_valid_not_nacked) begin
      if (_T_320) begin
        _T_639_state <= s1_meta_uncorrected_3_coh_state;
      end else if (_T_318) begin
        _T_639_state <= s1_meta_uncorrected_2_coh_state;
      end else if (_T_316) begin
        _T_639_state <= s1_meta_uncorrected_1_coh_state;
      end else begin
        _T_639_state <= s1_meta_uncorrected_0_coh_state;
      end
    end
    if (_T_831) begin
      lrscAddr <= s2_req_addr[31:6];
    end
    if (_T_847) begin
      pstore1_cmd <= s1_req_cmd;
    end
    if (_T_847) begin
      pstore1_data <= io_cpu_s1_data_data;
    end
    if (_T_847) begin
      pstore1_way <= s1_meta_hit_way;
    end
    if (_T_847) begin
      pstore1_rmw <= _T_902;
    end
    _T_976 <= io_cpu_s2_nack;
    if (advance_pstore1) begin
      pstore2_way <= pstore1_way;
    end
    if (advance_pstore1) begin
      _T_1032 <= pstore1_storegen_data[7:0];
    end
    if (advance_pstore1) begin
      _T_1037 <= pstore1_storegen_data[15:8];
    end
    if (advance_pstore1) begin
      _T_1042 <= pstore1_storegen_data[23:16];
    end
    if (advance_pstore1) begin
      _T_1047 <= pstore1_storegen_data[31:24];
    end
    s1_release_data_valid <= dataArb_io_in_2_ready & dataArb_io_in_2_valid;
    _T_2470 <= tlb_io_req_valid & _T_20;
    doUncachedResp <= io_cpu_replay_next;
    if (reset) begin
      resetting <= 1'h0;
    end else if (resetting) begin
      if (flushDone) begin
        resetting <= 1'h0;
      end else begin
        resetting <= _GEN_337;
      end
    end else begin
      resetting <= _GEN_337;
    end
    _T_2523 <= reset;
    if (reset) begin
      flushCounter <= 8'hc0;
    end else begin
      flushCounter <= _GEN_339[7:0];
    end
    if (reset) begin
      _T_2604 <= 10'h0;
    end else if (_T_2354) begin
      if (_T_2607) begin
        if (tl_out__c_bits_opcode[0]) begin
          _T_2604 <= _T_2358[11:2];
        end else begin
          _T_2604 <= 10'h0;
        end
      end else begin
        _T_2604 <= _T_2606;
      end
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_166) begin
          $fwrite(32'h80000002,"Assertion failed\n    at DCache.scala:1081 assert(!needsRead(req) || res)\n"); // @[DCache.scala 1081:11:freechips.rocketchip.system.DefaultRV32Config.fir@192432.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_166) begin
          $fatal; // @[DCache.scala 1081:11:freechips.rocketchip.system.DefaultRV32Config.fir@192433.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_355) begin
          $fwrite(32'h80000002,"Assertion failed\n    at DCache.scala:281 assert(!(s1_valid_masked && s1_req.cmd === M_PWR) || (s1_mask_xwr | ~io.cpu.s1_data.mask).andR)\n"); // @[DCache.scala 281:9:freechips.rocketchip.system.DefaultRV32Config.fir@192751.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_355) begin
          $fatal; // @[DCache.scala 281:9:freechips.rocketchip.system.DefaultRV32Config.fir@192752.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_166) begin
          $fwrite(32'h80000002,"Assertion failed\n    at DCache.scala:1081 assert(!needsRead(req) || res)\n"); // @[DCache.scala 1081:11:freechips.rocketchip.system.DefaultRV32Config.fir@193635.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_166) begin
          $fatal; // @[DCache.scala 1081:11:freechips.rocketchip.system.DefaultRV32Config.fir@193636.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_995) begin
          $fwrite(32'h80000002,"Assertion failed\n    at DCache.scala:461 assert(pstore1_rmw || pstore1_valid_not_rmw(io.cpu.s2_kill) === pstore1_valid)\n"); // @[DCache.scala 461:9:freechips.rocketchip.system.DefaultRV32Config.fir@193671.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_995) begin
          $fatal; // @[DCache.scala 461:9:freechips.rocketchip.system.DefaultRV32Config.fir@193672.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_385 & _T_2220) begin
          $fwrite(32'h80000002,"Assertion failed: A GrantData was unexpected by the dcache.\n    at DCache.scala:620 assert(cached_grant_wait, \"A GrantData was unexpected by the dcache.\")\n"); // @[DCache.scala 620:13:freechips.rocketchip.system.DefaultRV32Config.fir@195113.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_385 & _T_2220) begin
          $fatal; // @[DCache.scala 620:13:freechips.rocketchip.system.DefaultRV32Config.fir@195114.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_390 & _T_2225) begin
          $fwrite(32'h80000002,"Assertion failed: An AccessAck was unexpected by the dcache.\n    at DCache.scala:630 assert(f, \"An AccessAck was unexpected by the dcache.\") // TODO must handle Ack coming back on same cycle!\n"); // @[DCache.scala 630:17:freechips.rocketchip.system.DefaultRV32Config.fir@195132.14]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_390 & _T_2225) begin
          $fatal; // @[DCache.scala 630:17:freechips.rocketchip.system.DefaultRV32Config.fir@195133.14]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_399 & _T_2232) begin
          $fwrite(32'h80000002,"Assertion failed: A ReleaseAck was unexpected by the dcache.\n    at DCache.scala:651 assert(release_ack_wait, \"A ReleaseAck was unexpected by the dcache.\") // TODO should handle Ack coming back on same cycle!\n"); // @[DCache.scala 651:13:freechips.rocketchip.system.DefaultRV32Config.fir@195158.14]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_399 & _T_2232) begin
          $fatal; // @[DCache.scala 651:13:freechips.rocketchip.system.DefaultRV32Config.fir@195159.14]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2244) begin
          $fwrite(32'h80000002,"Assertion failed\n    at DCache.scala:659 assert(tl_out.e.fire() === (tl_out.d.fire() && d_first && grantIsCached))\n"); // @[DCache.scala 659:9:freechips.rocketchip.system.DefaultRV32Config.fir@195181.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_2244) begin
          $fatal; // @[DCache.scala 659:9:freechips.rocketchip.system.DefaultRV32Config.fir@195182.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (s2_want_victimize & _T_2388) begin
          $fwrite(32'h80000002,"Assertion failed\n    at DCache.scala:739 assert(s2_valid_flush_line || s2_flush_valid || io.cpu.s2_nack)\n"); // @[DCache.scala 739:13:freechips.rocketchip.system.DefaultRV32Config.fir@195421.8]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (s2_want_victimize & _T_2388) begin
          $fatal; // @[DCache.scala 739:13:freechips.rocketchip.system.DefaultRV32Config.fir@195422.8]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (doUncachedResp & _T_2484) begin
          $fwrite(32'h80000002,"Assertion failed\n    at DCache.scala:851 assert(!s2_valid_hit)\n"); // @[DCache.scala 851:11:freechips.rocketchip.system.DefaultRV32Config.fir@195659.8]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (doUncachedResp & _T_2484) begin
          $fatal; // @[DCache.scala 851:11:freechips.rocketchip.system.DefaultRV32Config.fir@195660.8]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
  end
endmodule
