module OptimizationBarrier_118( // @[:freechips.rocketchip.system.DefaultRV32Config.fir@214059.2]
  input  [53:0] io_x_ppn, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@214062.4]
  input         io_x_d, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@214062.4]
  input         io_x_a, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@214062.4]
  input         io_x_g, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@214062.4]
  input         io_x_u, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@214062.4]
  input         io_x_x, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@214062.4]
  input         io_x_w, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@214062.4]
  input         io_x_r, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@214062.4]
  input         io_x_v, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@214062.4]
  output [53:0] io_y_ppn, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@214062.4]
  output        io_y_d, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@214062.4]
  output        io_y_a, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@214062.4]
  output        io_y_g, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@214062.4]
  output        io_y_u, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@214062.4]
  output        io_y_x, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@214062.4]
  output        io_y_w, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@214062.4]
  output        io_y_r, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@214062.4]
  output        io_y_v // @[:freechips.rocketchip.system.DefaultRV32Config.fir@214062.4]
);
  assign io_y_ppn = io_x_ppn; // @[package.scala 236:12:freechips.rocketchip.system.DefaultRV32Config.fir@214067.4]
  assign io_y_d = io_x_d; // @[package.scala 236:12:freechips.rocketchip.system.DefaultRV32Config.fir@214067.4]
  assign io_y_a = io_x_a; // @[package.scala 236:12:freechips.rocketchip.system.DefaultRV32Config.fir@214067.4]
  assign io_y_g = io_x_g; // @[package.scala 236:12:freechips.rocketchip.system.DefaultRV32Config.fir@214067.4]
  assign io_y_u = io_x_u; // @[package.scala 236:12:freechips.rocketchip.system.DefaultRV32Config.fir@214067.4]
  assign io_y_x = io_x_x; // @[package.scala 236:12:freechips.rocketchip.system.DefaultRV32Config.fir@214067.4]
  assign io_y_w = io_x_w; // @[package.scala 236:12:freechips.rocketchip.system.DefaultRV32Config.fir@214067.4]
  assign io_y_r = io_x_r; // @[package.scala 236:12:freechips.rocketchip.system.DefaultRV32Config.fir@214067.4]
  assign io_y_v = io_x_v; // @[package.scala 236:12:freechips.rocketchip.system.DefaultRV32Config.fir@214067.4]
endmodule
