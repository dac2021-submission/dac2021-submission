module RecFNToIN( // @[:freechips.rocketchip.system.DefaultRV32Config.fir@211878.2]
  input  [32:0] io_in, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@211879.4]
  input  [2:0]  io_roundingMode, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@211879.4]
  input         io_signedOut, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@211879.4]
  output [31:0] io_out, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@211879.4]
  output [2:0]  io_intExceptionFlags // @[:freechips.rocketchip.system.DefaultRV32Config.fir@211879.4]
);
  wire  rawIn_isZero; // @[rawFloatFromRecFN.scala 51:54:freechips.rocketchip.system.DefaultRV32Config.fir@211884.4]
  wire  _T_4; // @[rawFloatFromRecFN.scala 52:54:freechips.rocketchip.system.DefaultRV32Config.fir@211886.4]
  wire  rawIn_isNaN; // @[rawFloatFromRecFN.scala 55:33:freechips.rocketchip.system.DefaultRV32Config.fir@211890.4]
  wire  _T_8; // @[rawFloatFromRecFN.scala 56:36:freechips.rocketchip.system.DefaultRV32Config.fir@211893.4]
  wire  rawIn_isInf; // @[rawFloatFromRecFN.scala 56:33:freechips.rocketchip.system.DefaultRV32Config.fir@211894.4]
  wire  rawIn_sign; // @[rawFloatFromRecFN.scala 58:25:freechips.rocketchip.system.DefaultRV32Config.fir@211897.4]
  wire [9:0] rawIn_sExp; // @[rawFloatFromRecFN.scala 59:27:freechips.rocketchip.system.DefaultRV32Config.fir@211899.4]
  wire  _T_12; // @[rawFloatFromRecFN.scala 60:39:freechips.rocketchip.system.DefaultRV32Config.fir@211901.4]
  wire [24:0] rawIn_sig; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@211904.4]
  wire  magGeOne; // @[RecFNToIN.scala 58:30:freechips.rocketchip.system.DefaultRV32Config.fir@211906.4]
  wire [7:0] posExp; // @[RecFNToIN.scala 59:28:freechips.rocketchip.system.DefaultRV32Config.fir@211907.4]
  wire  _T_16; // @[RecFNToIN.scala 60:27:freechips.rocketchip.system.DefaultRV32Config.fir@211908.4]
  wire  _T_17; // @[RecFNToIN.scala 60:47:freechips.rocketchip.system.DefaultRV32Config.fir@211909.4]
  wire  magJustBelowOne; // @[RecFNToIN.scala 60:37:freechips.rocketchip.system.DefaultRV32Config.fir@211910.4]
  wire  roundingMode_near_even; // @[RecFNToIN.scala 64:53:freechips.rocketchip.system.DefaultRV32Config.fir@211911.4]
  wire  roundingMode_min; // @[RecFNToIN.scala 66:53:freechips.rocketchip.system.DefaultRV32Config.fir@211913.4]
  wire  roundingMode_max; // @[RecFNToIN.scala 67:53:freechips.rocketchip.system.DefaultRV32Config.fir@211914.4]
  wire  roundingMode_near_maxMag; // @[RecFNToIN.scala 68:53:freechips.rocketchip.system.DefaultRV32Config.fir@211915.4]
  wire  roundingMode_odd; // @[RecFNToIN.scala 69:53:freechips.rocketchip.system.DefaultRV32Config.fir@211916.4]
  wire [23:0] _T_19; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@211918.4]
  wire [4:0] _T_21; // @[RecFNToIN.scala 81:16:freechips.rocketchip.system.DefaultRV32Config.fir@211920.4]
  wire [54:0] _GEN_0; // @[RecFNToIN.scala 80:50:freechips.rocketchip.system.DefaultRV32Config.fir@211921.4]
  wire [54:0] shiftedSig; // @[RecFNToIN.scala 80:50:freechips.rocketchip.system.DefaultRV32Config.fir@211921.4]
  wire  _T_24; // @[RecFNToIN.scala 86:69:freechips.rocketchip.system.DefaultRV32Config.fir@211924.4]
  wire [33:0] alignedSig; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@211925.4]
  wire [31:0] unroundedInt; // @[RecFNToIN.scala 87:54:freechips.rocketchip.system.DefaultRV32Config.fir@211926.4]
  wire  _T_27; // @[RecFNToIN.scala 89:57:freechips.rocketchip.system.DefaultRV32Config.fir@211929.4]
  wire  common_inexact; // @[RecFNToIN.scala 89:29:freechips.rocketchip.system.DefaultRV32Config.fir@211931.4]
  wire  _T_30; // @[RecFNToIN.scala 91:46:freechips.rocketchip.system.DefaultRV32Config.fir@211933.4]
  wire  _T_32; // @[RecFNToIN.scala 91:71:freechips.rocketchip.system.DefaultRV32Config.fir@211935.4]
  wire  _T_33; // @[RecFNToIN.scala 91:51:freechips.rocketchip.system.DefaultRV32Config.fir@211936.4]
  wire  _T_34; // @[RecFNToIN.scala 91:25:freechips.rocketchip.system.DefaultRV32Config.fir@211937.4]
  wire  _T_37; // @[RecFNToIN.scala 92:26:freechips.rocketchip.system.DefaultRV32Config.fir@211940.4]
  wire  roundIncr_near_even; // @[RecFNToIN.scala 91:78:freechips.rocketchip.system.DefaultRV32Config.fir@211941.4]
  wire  _T_39; // @[RecFNToIN.scala 93:43:freechips.rocketchip.system.DefaultRV32Config.fir@211943.4]
  wire  roundIncr_near_maxMag; // @[RecFNToIN.scala 93:61:freechips.rocketchip.system.DefaultRV32Config.fir@211944.4]
  wire  _T_40; // @[RecFNToIN.scala 95:35:freechips.rocketchip.system.DefaultRV32Config.fir@211945.4]
  wire  _T_41; // @[RecFNToIN.scala 96:35:freechips.rocketchip.system.DefaultRV32Config.fir@211946.4]
  wire  _T_42; // @[RecFNToIN.scala 95:61:freechips.rocketchip.system.DefaultRV32Config.fir@211947.4]
  wire  _T_43; // @[RecFNToIN.scala 97:28:freechips.rocketchip.system.DefaultRV32Config.fir@211948.4]
  wire  _T_44; // @[RecFNToIN.scala 98:26:freechips.rocketchip.system.DefaultRV32Config.fir@211949.4]
  wire  _T_45; // @[RecFNToIN.scala 97:49:freechips.rocketchip.system.DefaultRV32Config.fir@211950.4]
  wire  _T_46; // @[RecFNToIN.scala 96:61:freechips.rocketchip.system.DefaultRV32Config.fir@211951.4]
  wire  _T_47; // @[RecFNToIN.scala 99:31:freechips.rocketchip.system.DefaultRV32Config.fir@211952.4]
  wire  _T_48; // @[RecFNToIN.scala 99:43:freechips.rocketchip.system.DefaultRV32Config.fir@211953.4]
  wire  _T_49; // @[RecFNToIN.scala 99:27:freechips.rocketchip.system.DefaultRV32Config.fir@211954.4]
  wire  roundIncr; // @[RecFNToIN.scala 98:46:freechips.rocketchip.system.DefaultRV32Config.fir@211955.4]
  wire [31:0] _T_50; // @[RecFNToIN.scala 100:45:freechips.rocketchip.system.DefaultRV32Config.fir@211956.4]
  wire [31:0] complUnroundedInt; // @[RecFNToIN.scala 100:32:freechips.rocketchip.system.DefaultRV32Config.fir@211957.4]
  wire  _T_51; // @[RecFNToIN.scala 102:23:freechips.rocketchip.system.DefaultRV32Config.fir@211958.4]
  wire [31:0] _T_53; // @[RecFNToIN.scala 103:31:freechips.rocketchip.system.DefaultRV32Config.fir@211960.4]
  wire [31:0] _T_54; // @[RecFNToIN.scala 102:12:freechips.rocketchip.system.DefaultRV32Config.fir@211961.4]
  wire  _T_55; // @[RecFNToIN.scala 105:31:freechips.rocketchip.system.DefaultRV32Config.fir@211962.4]
  wire [31:0] _GEN_1; // @[RecFNToIN.scala 105:11:freechips.rocketchip.system.DefaultRV32Config.fir@211963.4]
  wire [31:0] roundedInt; // @[RecFNToIN.scala 105:11:freechips.rocketchip.system.DefaultRV32Config.fir@211963.4]
  wire  magGeOne_atOverflowEdge; // @[RecFNToIN.scala 107:43:freechips.rocketchip.system.DefaultRV32Config.fir@211964.4]
  wire  _T_57; // @[RecFNToIN.scala 110:56:freechips.rocketchip.system.DefaultRV32Config.fir@211966.4]
  wire  roundCarryBut2; // @[RecFNToIN.scala 110:61:freechips.rocketchip.system.DefaultRV32Config.fir@211967.4]
  wire  _T_58; // @[RecFNToIN.scala 113:21:freechips.rocketchip.system.DefaultRV32Config.fir@211968.4]
  wire  _T_60; // @[RecFNToIN.scala 117:60:freechips.rocketchip.system.DefaultRV32Config.fir@211970.4]
  wire  _T_61; // @[RecFNToIN.scala 117:64:freechips.rocketchip.system.DefaultRV32Config.fir@211971.4]
  wire  _T_62; // @[RecFNToIN.scala 116:49:freechips.rocketchip.system.DefaultRV32Config.fir@211972.4]
  wire  _T_63; // @[RecFNToIN.scala 119:38:freechips.rocketchip.system.DefaultRV32Config.fir@211973.4]
  wire  _T_64; // @[RecFNToIN.scala 119:62:freechips.rocketchip.system.DefaultRV32Config.fir@211974.4]
  wire  _T_65; // @[RecFNToIN.scala 118:49:freechips.rocketchip.system.DefaultRV32Config.fir@211975.4]
  wire  _T_66; // @[RecFNToIN.scala 115:24:freechips.rocketchip.system.DefaultRV32Config.fir@211976.4]
  wire  _T_68; // @[RecFNToIN.scala 122:50:freechips.rocketchip.system.DefaultRV32Config.fir@211978.4]
  wire  _T_69; // @[RecFNToIN.scala 123:57:freechips.rocketchip.system.DefaultRV32Config.fir@211979.4]
  wire  _T_70; // @[RecFNToIN.scala 121:32:freechips.rocketchip.system.DefaultRV32Config.fir@211980.4]
  wire  _T_71; // @[RecFNToIN.scala 114:20:freechips.rocketchip.system.DefaultRV32Config.fir@211981.4]
  wire  _T_72; // @[RecFNToIN.scala 113:40:freechips.rocketchip.system.DefaultRV32Config.fir@211982.4]
  wire  _T_73; // @[RecFNToIN.scala 125:13:freechips.rocketchip.system.DefaultRV32Config.fir@211983.4]
  wire  _T_74; // @[RecFNToIN.scala 125:27:freechips.rocketchip.system.DefaultRV32Config.fir@211984.4]
  wire  _T_75; // @[RecFNToIN.scala 125:41:freechips.rocketchip.system.DefaultRV32Config.fir@211985.4]
  wire  common_overflow; // @[RecFNToIN.scala 112:12:freechips.rocketchip.system.DefaultRV32Config.fir@211986.4]
  wire  invalidExc; // @[RecFNToIN.scala 130:34:freechips.rocketchip.system.DefaultRV32Config.fir@211987.4]
  wire  _T_76; // @[RecFNToIN.scala 131:20:freechips.rocketchip.system.DefaultRV32Config.fir@211988.4]
  wire  overflow; // @[RecFNToIN.scala 131:32:freechips.rocketchip.system.DefaultRV32Config.fir@211989.4]
  wire  _T_78; // @[RecFNToIN.scala 132:35:freechips.rocketchip.system.DefaultRV32Config.fir@211991.4]
  wire  _T_79; // @[RecFNToIN.scala 132:32:freechips.rocketchip.system.DefaultRV32Config.fir@211992.4]
  wire  inexact; // @[RecFNToIN.scala 132:52:freechips.rocketchip.system.DefaultRV32Config.fir@211993.4]
  wire  _T_80; // @[RecFNToIN.scala 134:19:freechips.rocketchip.system.DefaultRV32Config.fir@211994.4]
  wire  excSign; // @[RecFNToIN.scala 134:32:freechips.rocketchip.system.DefaultRV32Config.fir@211995.4]
  wire  _T_81; // @[RecFNToIN.scala 136:27:freechips.rocketchip.system.DefaultRV32Config.fir@211996.4]
  wire [31:0] _T_82; // @[RecFNToIN.scala 136:12:freechips.rocketchip.system.DefaultRV32Config.fir@211997.4]
  wire  _T_83; // @[RecFNToIN.scala 140:13:freechips.rocketchip.system.DefaultRV32Config.fir@211998.4]
  wire [30:0] _T_84; // @[RecFNToIN.scala 140:12:freechips.rocketchip.system.DefaultRV32Config.fir@211999.4]
  wire [31:0] _GEN_2; // @[RecFNToIN.scala 139:11:freechips.rocketchip.system.DefaultRV32Config.fir@212000.4]
  wire [31:0] excOut; // @[RecFNToIN.scala 139:11:freechips.rocketchip.system.DefaultRV32Config.fir@212000.4]
  wire  _T_85; // @[RecFNToIN.scala 142:30:freechips.rocketchip.system.DefaultRV32Config.fir@212001.4]
  wire [1:0] _T_87; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@212004.4]
  assign rawIn_isZero = io_in[31:29] == 3'h0; // @[rawFloatFromRecFN.scala 51:54:freechips.rocketchip.system.DefaultRV32Config.fir@211884.4]
  assign _T_4 = io_in[31:30] == 2'h3; // @[rawFloatFromRecFN.scala 52:54:freechips.rocketchip.system.DefaultRV32Config.fir@211886.4]
  assign rawIn_isNaN = _T_4 & io_in[29]; // @[rawFloatFromRecFN.scala 55:33:freechips.rocketchip.system.DefaultRV32Config.fir@211890.4]
  assign _T_8 = ~io_in[29]; // @[rawFloatFromRecFN.scala 56:36:freechips.rocketchip.system.DefaultRV32Config.fir@211893.4]
  assign rawIn_isInf = _T_4 & _T_8; // @[rawFloatFromRecFN.scala 56:33:freechips.rocketchip.system.DefaultRV32Config.fir@211894.4]
  assign rawIn_sign = io_in[32]; // @[rawFloatFromRecFN.scala 58:25:freechips.rocketchip.system.DefaultRV32Config.fir@211897.4]
  assign rawIn_sExp = {1'b0,$signed(io_in[31:23])}; // @[rawFloatFromRecFN.scala 59:27:freechips.rocketchip.system.DefaultRV32Config.fir@211899.4]
  assign _T_12 = ~rawIn_isZero; // @[rawFloatFromRecFN.scala 60:39:freechips.rocketchip.system.DefaultRV32Config.fir@211901.4]
  assign rawIn_sig = {1'h0,_T_12,io_in[22:0]}; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@211904.4]
  assign magGeOne = rawIn_sExp[8]; // @[RecFNToIN.scala 58:30:freechips.rocketchip.system.DefaultRV32Config.fir@211906.4]
  assign posExp = rawIn_sExp[7:0]; // @[RecFNToIN.scala 59:28:freechips.rocketchip.system.DefaultRV32Config.fir@211907.4]
  assign _T_16 = ~magGeOne; // @[RecFNToIN.scala 60:27:freechips.rocketchip.system.DefaultRV32Config.fir@211908.4]
  assign _T_17 = &posExp; // @[RecFNToIN.scala 60:47:freechips.rocketchip.system.DefaultRV32Config.fir@211909.4]
  assign magJustBelowOne = _T_16 & _T_17; // @[RecFNToIN.scala 60:37:freechips.rocketchip.system.DefaultRV32Config.fir@211910.4]
  assign roundingMode_near_even = io_roundingMode == 3'h0; // @[RecFNToIN.scala 64:53:freechips.rocketchip.system.DefaultRV32Config.fir@211911.4]
  assign roundingMode_min = io_roundingMode == 3'h2; // @[RecFNToIN.scala 66:53:freechips.rocketchip.system.DefaultRV32Config.fir@211913.4]
  assign roundingMode_max = io_roundingMode == 3'h3; // @[RecFNToIN.scala 67:53:freechips.rocketchip.system.DefaultRV32Config.fir@211914.4]
  assign roundingMode_near_maxMag = io_roundingMode == 3'h4; // @[RecFNToIN.scala 68:53:freechips.rocketchip.system.DefaultRV32Config.fir@211915.4]
  assign roundingMode_odd = io_roundingMode == 3'h6; // @[RecFNToIN.scala 69:53:freechips.rocketchip.system.DefaultRV32Config.fir@211916.4]
  assign _T_19 = {magGeOne,rawIn_sig[22:0]}; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@211918.4]
  assign _T_21 = magGeOne ? rawIn_sExp[4:0] : 5'h0; // @[RecFNToIN.scala 81:16:freechips.rocketchip.system.DefaultRV32Config.fir@211920.4]
  assign _GEN_0 = {{31'd0}, _T_19}; // @[RecFNToIN.scala 80:50:freechips.rocketchip.system.DefaultRV32Config.fir@211921.4]
  assign shiftedSig = _GEN_0 << _T_21; // @[RecFNToIN.scala 80:50:freechips.rocketchip.system.DefaultRV32Config.fir@211921.4]
  assign _T_24 = |shiftedSig[21:0]; // @[RecFNToIN.scala 86:69:freechips.rocketchip.system.DefaultRV32Config.fir@211924.4]
  assign alignedSig = {shiftedSig[54:22],_T_24}; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@211925.4]
  assign unroundedInt = alignedSig[33:2]; // @[RecFNToIN.scala 87:54:freechips.rocketchip.system.DefaultRV32Config.fir@211926.4]
  assign _T_27 = |alignedSig[1:0]; // @[RecFNToIN.scala 89:57:freechips.rocketchip.system.DefaultRV32Config.fir@211929.4]
  assign common_inexact = magGeOne ? _T_27 : _T_12; // @[RecFNToIN.scala 89:29:freechips.rocketchip.system.DefaultRV32Config.fir@211931.4]
  assign _T_30 = &alignedSig[2:1]; // @[RecFNToIN.scala 91:46:freechips.rocketchip.system.DefaultRV32Config.fir@211933.4]
  assign _T_32 = &alignedSig[1:0]; // @[RecFNToIN.scala 91:71:freechips.rocketchip.system.DefaultRV32Config.fir@211935.4]
  assign _T_33 = _T_30 | _T_32; // @[RecFNToIN.scala 91:51:freechips.rocketchip.system.DefaultRV32Config.fir@211936.4]
  assign _T_34 = magGeOne & _T_33; // @[RecFNToIN.scala 91:25:freechips.rocketchip.system.DefaultRV32Config.fir@211937.4]
  assign _T_37 = magJustBelowOne & _T_27; // @[RecFNToIN.scala 92:26:freechips.rocketchip.system.DefaultRV32Config.fir@211940.4]
  assign roundIncr_near_even = _T_34 | _T_37; // @[RecFNToIN.scala 91:78:freechips.rocketchip.system.DefaultRV32Config.fir@211941.4]
  assign _T_39 = magGeOne & alignedSig[1]; // @[RecFNToIN.scala 93:43:freechips.rocketchip.system.DefaultRV32Config.fir@211943.4]
  assign roundIncr_near_maxMag = _T_39 | magJustBelowOne; // @[RecFNToIN.scala 93:61:freechips.rocketchip.system.DefaultRV32Config.fir@211944.4]
  assign _T_40 = roundingMode_near_even & roundIncr_near_even; // @[RecFNToIN.scala 95:35:freechips.rocketchip.system.DefaultRV32Config.fir@211945.4]
  assign _T_41 = roundingMode_near_maxMag & roundIncr_near_maxMag; // @[RecFNToIN.scala 96:35:freechips.rocketchip.system.DefaultRV32Config.fir@211946.4]
  assign _T_42 = _T_40 | _T_41; // @[RecFNToIN.scala 95:61:freechips.rocketchip.system.DefaultRV32Config.fir@211947.4]
  assign _T_43 = roundingMode_min | roundingMode_odd; // @[RecFNToIN.scala 97:28:freechips.rocketchip.system.DefaultRV32Config.fir@211948.4]
  assign _T_44 = rawIn_sign & common_inexact; // @[RecFNToIN.scala 98:26:freechips.rocketchip.system.DefaultRV32Config.fir@211949.4]
  assign _T_45 = _T_43 & _T_44; // @[RecFNToIN.scala 97:49:freechips.rocketchip.system.DefaultRV32Config.fir@211950.4]
  assign _T_46 = _T_42 | _T_45; // @[RecFNToIN.scala 96:61:freechips.rocketchip.system.DefaultRV32Config.fir@211951.4]
  assign _T_47 = ~rawIn_sign; // @[RecFNToIN.scala 99:31:freechips.rocketchip.system.DefaultRV32Config.fir@211952.4]
  assign _T_48 = _T_47 & common_inexact; // @[RecFNToIN.scala 99:43:freechips.rocketchip.system.DefaultRV32Config.fir@211953.4]
  assign _T_49 = roundingMode_max & _T_48; // @[RecFNToIN.scala 99:27:freechips.rocketchip.system.DefaultRV32Config.fir@211954.4]
  assign roundIncr = _T_46 | _T_49; // @[RecFNToIN.scala 98:46:freechips.rocketchip.system.DefaultRV32Config.fir@211955.4]
  assign _T_50 = ~unroundedInt; // @[RecFNToIN.scala 100:45:freechips.rocketchip.system.DefaultRV32Config.fir@211956.4]
  assign complUnroundedInt = rawIn_sign ? _T_50 : unroundedInt; // @[RecFNToIN.scala 100:32:freechips.rocketchip.system.DefaultRV32Config.fir@211957.4]
  assign _T_51 = roundIncr ^ rawIn_sign; // @[RecFNToIN.scala 102:23:freechips.rocketchip.system.DefaultRV32Config.fir@211958.4]
  assign _T_53 = complUnroundedInt + 32'h1; // @[RecFNToIN.scala 103:31:freechips.rocketchip.system.DefaultRV32Config.fir@211960.4]
  assign _T_54 = _T_51 ? _T_53 : complUnroundedInt; // @[RecFNToIN.scala 102:12:freechips.rocketchip.system.DefaultRV32Config.fir@211961.4]
  assign _T_55 = roundingMode_odd & common_inexact; // @[RecFNToIN.scala 105:31:freechips.rocketchip.system.DefaultRV32Config.fir@211962.4]
  assign _GEN_1 = {{31'd0}, _T_55}; // @[RecFNToIN.scala 105:11:freechips.rocketchip.system.DefaultRV32Config.fir@211963.4]
  assign roundedInt = _T_54 | _GEN_1; // @[RecFNToIN.scala 105:11:freechips.rocketchip.system.DefaultRV32Config.fir@211963.4]
  assign magGeOne_atOverflowEdge = posExp == 8'h1f; // @[RecFNToIN.scala 107:43:freechips.rocketchip.system.DefaultRV32Config.fir@211964.4]
  assign _T_57 = &unroundedInt[29:0]; // @[RecFNToIN.scala 110:56:freechips.rocketchip.system.DefaultRV32Config.fir@211966.4]
  assign roundCarryBut2 = _T_57 & roundIncr; // @[RecFNToIN.scala 110:61:freechips.rocketchip.system.DefaultRV32Config.fir@211967.4]
  assign _T_58 = posExp >= 8'h20; // @[RecFNToIN.scala 113:21:freechips.rocketchip.system.DefaultRV32Config.fir@211968.4]
  assign _T_60 = |unroundedInt[30:0]; // @[RecFNToIN.scala 117:60:freechips.rocketchip.system.DefaultRV32Config.fir@211970.4]
  assign _T_61 = _T_60 | roundIncr; // @[RecFNToIN.scala 117:64:freechips.rocketchip.system.DefaultRV32Config.fir@211971.4]
  assign _T_62 = magGeOne_atOverflowEdge & _T_61; // @[RecFNToIN.scala 116:49:freechips.rocketchip.system.DefaultRV32Config.fir@211972.4]
  assign _T_63 = posExp == 8'h1e; // @[RecFNToIN.scala 119:38:freechips.rocketchip.system.DefaultRV32Config.fir@211973.4]
  assign _T_64 = _T_63 & roundCarryBut2; // @[RecFNToIN.scala 119:62:freechips.rocketchip.system.DefaultRV32Config.fir@211974.4]
  assign _T_65 = magGeOne_atOverflowEdge | _T_64; // @[RecFNToIN.scala 118:49:freechips.rocketchip.system.DefaultRV32Config.fir@211975.4]
  assign _T_66 = rawIn_sign ? _T_62 : _T_65; // @[RecFNToIN.scala 115:24:freechips.rocketchip.system.DefaultRV32Config.fir@211976.4]
  assign _T_68 = magGeOne_atOverflowEdge & unroundedInt[30]; // @[RecFNToIN.scala 122:50:freechips.rocketchip.system.DefaultRV32Config.fir@211978.4]
  assign _T_69 = _T_68 & roundCarryBut2; // @[RecFNToIN.scala 123:57:freechips.rocketchip.system.DefaultRV32Config.fir@211979.4]
  assign _T_70 = rawIn_sign | _T_69; // @[RecFNToIN.scala 121:32:freechips.rocketchip.system.DefaultRV32Config.fir@211980.4]
  assign _T_71 = io_signedOut ? _T_66 : _T_70; // @[RecFNToIN.scala 114:20:freechips.rocketchip.system.DefaultRV32Config.fir@211981.4]
  assign _T_72 = _T_58 | _T_71; // @[RecFNToIN.scala 113:40:freechips.rocketchip.system.DefaultRV32Config.fir@211982.4]
  assign _T_73 = ~io_signedOut; // @[RecFNToIN.scala 125:13:freechips.rocketchip.system.DefaultRV32Config.fir@211983.4]
  assign _T_74 = _T_73 & rawIn_sign; // @[RecFNToIN.scala 125:27:freechips.rocketchip.system.DefaultRV32Config.fir@211984.4]
  assign _T_75 = _T_74 & roundIncr; // @[RecFNToIN.scala 125:41:freechips.rocketchip.system.DefaultRV32Config.fir@211985.4]
  assign common_overflow = magGeOne ? _T_72 : _T_75; // @[RecFNToIN.scala 112:12:freechips.rocketchip.system.DefaultRV32Config.fir@211986.4]
  assign invalidExc = rawIn_isNaN | rawIn_isInf; // @[RecFNToIN.scala 130:34:freechips.rocketchip.system.DefaultRV32Config.fir@211987.4]
  assign _T_76 = ~invalidExc; // @[RecFNToIN.scala 131:20:freechips.rocketchip.system.DefaultRV32Config.fir@211988.4]
  assign overflow = _T_76 & common_overflow; // @[RecFNToIN.scala 131:32:freechips.rocketchip.system.DefaultRV32Config.fir@211989.4]
  assign _T_78 = ~common_overflow; // @[RecFNToIN.scala 132:35:freechips.rocketchip.system.DefaultRV32Config.fir@211991.4]
  assign _T_79 = _T_76 & _T_78; // @[RecFNToIN.scala 132:32:freechips.rocketchip.system.DefaultRV32Config.fir@211992.4]
  assign inexact = _T_79 & common_inexact; // @[RecFNToIN.scala 132:52:freechips.rocketchip.system.DefaultRV32Config.fir@211993.4]
  assign _T_80 = ~rawIn_isNaN; // @[RecFNToIN.scala 134:19:freechips.rocketchip.system.DefaultRV32Config.fir@211994.4]
  assign excSign = _T_80 & rawIn_sign; // @[RecFNToIN.scala 134:32:freechips.rocketchip.system.DefaultRV32Config.fir@211995.4]
  assign _T_81 = io_signedOut == excSign; // @[RecFNToIN.scala 136:27:freechips.rocketchip.system.DefaultRV32Config.fir@211996.4]
  assign _T_82 = _T_81 ? 32'h80000000 : 32'h0; // @[RecFNToIN.scala 136:12:freechips.rocketchip.system.DefaultRV32Config.fir@211997.4]
  assign _T_83 = ~excSign; // @[RecFNToIN.scala 140:13:freechips.rocketchip.system.DefaultRV32Config.fir@211998.4]
  assign _T_84 = _T_83 ? 31'h7fffffff : 31'h0; // @[RecFNToIN.scala 140:12:freechips.rocketchip.system.DefaultRV32Config.fir@211999.4]
  assign _GEN_2 = {{1'd0}, _T_84}; // @[RecFNToIN.scala 139:11:freechips.rocketchip.system.DefaultRV32Config.fir@212000.4]
  assign excOut = _T_82 | _GEN_2; // @[RecFNToIN.scala 139:11:freechips.rocketchip.system.DefaultRV32Config.fir@212000.4]
  assign _T_85 = invalidExc | common_overflow; // @[RecFNToIN.scala 142:30:freechips.rocketchip.system.DefaultRV32Config.fir@212001.4]
  assign _T_87 = {invalidExc,overflow}; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@212004.4]
  assign io_out = _T_85 ? excOut : roundedInt; // @[RecFNToIN.scala 142:12:freechips.rocketchip.system.DefaultRV32Config.fir@212003.4]
  assign io_intExceptionFlags = {_T_87,inexact}; // @[RecFNToIN.scala 143:26:freechips.rocketchip.system.DefaultRV32Config.fir@212006.4]
endmodule
