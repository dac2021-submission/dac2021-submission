module Arbiter( // @[:freechips.rocketchip.system.DefaultRV32Config.fir@214027.2]
  output        io_in_0_ready, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@214030.4]
  input         io_in_0_valid, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@214030.4]
  input  [19:0] io_in_0_bits_bits_addr, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@214030.4]
  output        io_in_1_ready, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@214030.4]
  input         io_in_1_valid, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@214030.4]
  input         io_in_1_bits_valid, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@214030.4]
  input  [19:0] io_in_1_bits_bits_addr, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@214030.4]
  input         io_out_ready, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@214030.4]
  output        io_out_valid, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@214030.4]
  output        io_out_bits_valid, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@214030.4]
  output [19:0] io_out_bits_bits_addr, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@214030.4]
  output        io_chosen // @[:freechips.rocketchip.system.DefaultRV32Config.fir@214030.4]
);
  wire  grant_1; // @[Arbiter.scala 31:78:freechips.rocketchip.system.DefaultRV32Config.fir@214040.4]
  wire  _T_2; // @[Arbiter.scala 135:19:freechips.rocketchip.system.DefaultRV32Config.fir@214045.4]
  assign grant_1 = ~io_in_0_valid; // @[Arbiter.scala 31:78:freechips.rocketchip.system.DefaultRV32Config.fir@214040.4]
  assign _T_2 = ~grant_1; // @[Arbiter.scala 135:19:freechips.rocketchip.system.DefaultRV32Config.fir@214045.4]
  assign io_in_0_ready = io_out_ready; // @[Arbiter.scala 134:14:freechips.rocketchip.system.DefaultRV32Config.fir@214042.4]
  assign io_in_1_ready = grant_1 & io_out_ready; // @[Arbiter.scala 134:14:freechips.rocketchip.system.DefaultRV32Config.fir@214044.4]
  assign io_out_valid = _T_2 | io_in_1_valid; // @[Arbiter.scala 135:16:freechips.rocketchip.system.DefaultRV32Config.fir@214047.4]
  assign io_out_bits_valid = io_in_0_valid | io_in_1_bits_valid; // @[Arbiter.scala 124:15:freechips.rocketchip.system.DefaultRV32Config.fir@214034.4 Arbiter.scala 128:19:freechips.rocketchip.system.DefaultRV32Config.fir@214038.6]
  assign io_out_bits_bits_addr = io_in_0_valid ? io_in_0_bits_bits_addr : io_in_1_bits_bits_addr; // @[Arbiter.scala 124:15:freechips.rocketchip.system.DefaultRV32Config.fir@214033.4 Arbiter.scala 128:19:freechips.rocketchip.system.DefaultRV32Config.fir@214037.6]
  assign io_chosen = io_in_0_valid ? 1'h0 : 1'h1; // @[Arbiter.scala 123:13:freechips.rocketchip.system.DefaultRV32Config.fir@214032.4 Arbiter.scala 127:17:freechips.rocketchip.system.DefaultRV32Config.fir@214036.6]
endmodule
