module TLMonitor_41( // @[:freechips.rocketchip.system.DefaultRV32Config.fir@99790.2]
  input        clock, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@99791.4]
  input        reset, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@99792.4]
  input        io_in_a_ready, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@99793.4]
  input        io_in_a_valid, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@99793.4]
  input  [2:0] io_in_a_bits_opcode, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@99793.4]
  input  [8:0] io_in_a_bits_address, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@99793.4]
  input  [3:0] io_in_a_bits_mask, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@99793.4]
  input        io_in_d_ready, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@99793.4]
  input        io_in_d_valid, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@99793.4]
  input  [2:0] io_in_d_bits_opcode, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@99793.4]
  input  [1:0] io_in_d_bits_param, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@99793.4]
  input  [1:0] io_in_d_bits_size, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@99793.4]
  input        io_in_d_bits_source, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@99793.4]
  input        io_in_d_bits_sink, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@99793.4]
  input        io_in_d_bits_denied, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@99793.4]
  input        io_in_d_bits_corrupt // @[:freechips.rocketchip.system.DefaultRV32Config.fir@99793.4]
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
`endif // RANDOMIZE_REG_INIT
  wire [31:0] plusarg_reader_out; // @[PlusArg.scala 80:11:freechips.rocketchip.system.DefaultRV32Config.fir@101288.4]
  wire [8:0] _T_10; // @[Edges.scala 22:16:freechips.rocketchip.system.DefaultRV32Config.fir@99812.6]
  wire  _T_11; // @[Edges.scala 22:24:freechips.rocketchip.system.DefaultRV32Config.fir@99813.6]
  wire [9:0] _T_48; // @[Parameters.scala 137:49:freechips.rocketchip.system.DefaultRV32Config.fir@99850.6]
  wire  _T_56; // @[Monitor.scala 79:25:freechips.rocketchip.system.DefaultRV32Config.fir@99862.6]
  wire [9:0] _T_61; // @[Parameters.scala 137:52:freechips.rocketchip.system.DefaultRV32Config.fir@99868.8]
  wire  _T_62; // @[Parameters.scala 137:67:freechips.rocketchip.system.DefaultRV32Config.fir@99869.8]
  wire [8:0] _T_63; // @[Parameters.scala 137:31:freechips.rocketchip.system.DefaultRV32Config.fir@99870.8]
  wire [9:0] _T_64; // @[Parameters.scala 137:49:freechips.rocketchip.system.DefaultRV32Config.fir@99871.8]
  wire [9:0] _T_66; // @[Parameters.scala 137:52:freechips.rocketchip.system.DefaultRV32Config.fir@99873.8]
  wire  _T_67; // @[Parameters.scala 137:67:freechips.rocketchip.system.DefaultRV32Config.fir@99874.8]
  wire [8:0] _T_68; // @[Parameters.scala 137:31:freechips.rocketchip.system.DefaultRV32Config.fir@99875.8]
  wire [9:0] _T_69; // @[Parameters.scala 137:49:freechips.rocketchip.system.DefaultRV32Config.fir@99876.8]
  wire [9:0] _T_71; // @[Parameters.scala 137:52:freechips.rocketchip.system.DefaultRV32Config.fir@99878.8]
  wire  _T_72; // @[Parameters.scala 137:67:freechips.rocketchip.system.DefaultRV32Config.fir@99879.8]
  wire [8:0] _T_73; // @[Parameters.scala 137:31:freechips.rocketchip.system.DefaultRV32Config.fir@99880.8]
  wire [9:0] _T_74; // @[Parameters.scala 137:49:freechips.rocketchip.system.DefaultRV32Config.fir@99881.8]
  wire [9:0] _T_76; // @[Parameters.scala 137:52:freechips.rocketchip.system.DefaultRV32Config.fir@99883.8]
  wire  _T_77; // @[Parameters.scala 137:67:freechips.rocketchip.system.DefaultRV32Config.fir@99884.8]
  wire [8:0] _T_78; // @[Parameters.scala 137:31:freechips.rocketchip.system.DefaultRV32Config.fir@99885.8]
  wire [9:0] _T_79; // @[Parameters.scala 137:49:freechips.rocketchip.system.DefaultRV32Config.fir@99886.8]
  wire [9:0] _T_81; // @[Parameters.scala 137:52:freechips.rocketchip.system.DefaultRV32Config.fir@99888.8]
  wire  _T_82; // @[Parameters.scala 137:67:freechips.rocketchip.system.DefaultRV32Config.fir@99889.8]
  wire [8:0] _T_83; // @[Parameters.scala 137:31:freechips.rocketchip.system.DefaultRV32Config.fir@99890.8]
  wire [9:0] _T_84; // @[Parameters.scala 137:49:freechips.rocketchip.system.DefaultRV32Config.fir@99891.8]
  wire [9:0] _T_86; // @[Parameters.scala 137:52:freechips.rocketchip.system.DefaultRV32Config.fir@99893.8]
  wire  _T_87; // @[Parameters.scala 137:67:freechips.rocketchip.system.DefaultRV32Config.fir@99894.8]
  wire  _T_88; // @[Parameters.scala 552:42:freechips.rocketchip.system.DefaultRV32Config.fir@99895.8]
  wire  _T_89; // @[Parameters.scala 552:42:freechips.rocketchip.system.DefaultRV32Config.fir@99896.8]
  wire  _T_90; // @[Parameters.scala 552:42:freechips.rocketchip.system.DefaultRV32Config.fir@99897.8]
  wire  _T_91; // @[Parameters.scala 552:42:freechips.rocketchip.system.DefaultRV32Config.fir@99898.8]
  wire  _T_92; // @[Parameters.scala 552:42:freechips.rocketchip.system.DefaultRV32Config.fir@99899.8]
  wire  _T_97; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@99904.8]
  wire  _T_109; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@99932.8]
  wire  _T_110; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@99933.8]
  wire [3:0] _T_115; // @[Monitor.scala 86:18:freechips.rocketchip.system.DefaultRV32Config.fir@99946.8]
  wire  _T_116; // @[Monitor.scala 86:31:freechips.rocketchip.system.DefaultRV32Config.fir@99947.8]
  wire  _T_118; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@99949.8]
  wire  _T_119; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@99950.8]
  wire  _T_124; // @[Monitor.scala 90:25:freechips.rocketchip.system.DefaultRV32Config.fir@99964.6]
  wire  _T_196; // @[Monitor.scala 102:25:freechips.rocketchip.system.DefaultRV32Config.fir@100074.6]
  wire  _T_239; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@100118.8]
  wire  _T_240; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@100119.8]
  wire  _T_251; // @[Monitor.scala 107:30:freechips.rocketchip.system.DefaultRV32Config.fir@100146.8]
  wire  _T_253; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@100148.8]
  wire  _T_254; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@100149.8]
  wire  _T_259; // @[Monitor.scala 111:25:freechips.rocketchip.system.DefaultRV32Config.fir@100163.6]
  wire  _T_318; // @[Monitor.scala 119:25:freechips.rocketchip.system.DefaultRV32Config.fir@100244.6]
  wire  _T_379; // @[Monitor.scala 127:25:freechips.rocketchip.system.DefaultRV32Config.fir@100327.6]
  wire  _T_435; // @[Monitor.scala 135:25:freechips.rocketchip.system.DefaultRV32Config.fir@100405.6]
  wire  _T_491; // @[Monitor.scala 143:25:freechips.rocketchip.system.DefaultRV32Config.fir@100483.6]
  wire  _T_551; // @[Bundles.scala 44:24:freechips.rocketchip.system.DefaultRV32Config.fir@100571.6]
  wire  _T_553; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@100573.6]
  wire  _T_554; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@100574.6]
  wire  _T_555; // @[Parameters.scala 47:9:freechips.rocketchip.system.DefaultRV32Config.fir@100579.6]
  wire  _T_558; // @[Monitor.scala 307:25:freechips.rocketchip.system.DefaultRV32Config.fir@100584.6]
  wire  _T_560; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@100587.8]
  wire  _T_561; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@100588.8]
  wire  _T_562; // @[Monitor.scala 309:27:freechips.rocketchip.system.DefaultRV32Config.fir@100593.8]
  wire  _T_564; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@100595.8]
  wire  _T_565; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@100596.8]
  wire  _T_566; // @[Monitor.scala 310:28:freechips.rocketchip.system.DefaultRV32Config.fir@100601.8]
  wire  _T_568; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@100603.8]
  wire  _T_569; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@100604.8]
  wire  _T_570; // @[Monitor.scala 311:15:freechips.rocketchip.system.DefaultRV32Config.fir@100609.8]
  wire  _T_572; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@100611.8]
  wire  _T_573; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@100612.8]
  wire  _T_574; // @[Monitor.scala 312:15:freechips.rocketchip.system.DefaultRV32Config.fir@100617.8]
  wire  _T_576; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@100619.8]
  wire  _T_577; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@100620.8]
  wire  _T_578; // @[Monitor.scala 315:25:freechips.rocketchip.system.DefaultRV32Config.fir@100626.6]
  wire  _T_589; // @[Bundles.scala 104:26:freechips.rocketchip.system.DefaultRV32Config.fir@100650.8]
  wire  _T_591; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@100652.8]
  wire  _T_592; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@100653.8]
  wire  _T_593; // @[Monitor.scala 320:28:freechips.rocketchip.system.DefaultRV32Config.fir@100658.8]
  wire  _T_595; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@100660.8]
  wire  _T_596; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@100661.8]
  wire  _T_606; // @[Monitor.scala 325:25:freechips.rocketchip.system.DefaultRV32Config.fir@100684.6]
  wire  _T_626; // @[Monitor.scala 331:30:freechips.rocketchip.system.DefaultRV32Config.fir@100725.8]
  wire  _T_628; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@100727.8]
  wire  _T_629; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@100728.8]
  wire  _T_635; // @[Monitor.scala 335:25:freechips.rocketchip.system.DefaultRV32Config.fir@100743.6]
  wire  _T_652; // @[Monitor.scala 343:25:freechips.rocketchip.system.DefaultRV32Config.fir@100778.6]
  wire  _T_670; // @[Monitor.scala 351:25:freechips.rocketchip.system.DefaultRV32Config.fir@100814.6]
  wire  _T_702; // @[Decoupled.scala 40:37:freechips.rocketchip.system.DefaultRV32Config.fir@100880.4]
  reg  _T_711; // @[Edges.scala 230:27:freechips.rocketchip.system.DefaultRV32Config.fir@100889.4]
  wire  _T_713; // @[Edges.scala 231:28:freechips.rocketchip.system.DefaultRV32Config.fir@100891.4]
  wire  _T_714; // @[Edges.scala 232:25:freechips.rocketchip.system.DefaultRV32Config.fir@100892.4]
  reg [2:0] _T_722; // @[Monitor.scala 381:22:freechips.rocketchip.system.DefaultRV32Config.fir@100903.4]
  reg [8:0] _T_726; // @[Monitor.scala 385:22:freechips.rocketchip.system.DefaultRV32Config.fir@100907.4]
  wire  _T_727; // @[Monitor.scala 386:22:freechips.rocketchip.system.DefaultRV32Config.fir@100908.4]
  wire  _T_728; // @[Monitor.scala 386:19:freechips.rocketchip.system.DefaultRV32Config.fir@100909.4]
  wire  _T_729; // @[Monitor.scala 387:32:freechips.rocketchip.system.DefaultRV32Config.fir@100911.6]
  wire  _T_731; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@100913.6]
  wire  _T_732; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@100914.6]
  wire  _T_745; // @[Monitor.scala 391:32:freechips.rocketchip.system.DefaultRV32Config.fir@100943.6]
  wire  _T_747; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@100945.6]
  wire  _T_748; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@100946.6]
  wire  _T_750; // @[Monitor.scala 393:20:freechips.rocketchip.system.DefaultRV32Config.fir@100953.4]
  wire  _T_751; // @[Decoupled.scala 40:37:freechips.rocketchip.system.DefaultRV32Config.fir@100961.4]
  reg  _T_759; // @[Edges.scala 230:27:freechips.rocketchip.system.DefaultRV32Config.fir@100969.4]
  wire  _T_761; // @[Edges.scala 231:28:freechips.rocketchip.system.DefaultRV32Config.fir@100971.4]
  wire  _T_762; // @[Edges.scala 232:25:freechips.rocketchip.system.DefaultRV32Config.fir@100972.4]
  reg [2:0] _T_770; // @[Monitor.scala 532:22:freechips.rocketchip.system.DefaultRV32Config.fir@100983.4]
  reg [1:0] _T_771; // @[Monitor.scala 533:22:freechips.rocketchip.system.DefaultRV32Config.fir@100984.4]
  reg [1:0] _T_772; // @[Monitor.scala 534:22:freechips.rocketchip.system.DefaultRV32Config.fir@100985.4]
  reg  _T_773; // @[Monitor.scala 535:22:freechips.rocketchip.system.DefaultRV32Config.fir@100986.4]
  reg  _T_774; // @[Monitor.scala 536:22:freechips.rocketchip.system.DefaultRV32Config.fir@100987.4]
  reg  _T_775; // @[Monitor.scala 537:22:freechips.rocketchip.system.DefaultRV32Config.fir@100988.4]
  wire  _T_776; // @[Monitor.scala 538:22:freechips.rocketchip.system.DefaultRV32Config.fir@100989.4]
  wire  _T_777; // @[Monitor.scala 538:19:freechips.rocketchip.system.DefaultRV32Config.fir@100990.4]
  wire  _T_778; // @[Monitor.scala 539:29:freechips.rocketchip.system.DefaultRV32Config.fir@100992.6]
  wire  _T_780; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@100994.6]
  wire  _T_781; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@100995.6]
  wire  _T_782; // @[Monitor.scala 540:29:freechips.rocketchip.system.DefaultRV32Config.fir@101000.6]
  wire  _T_784; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@101002.6]
  wire  _T_785; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@101003.6]
  wire  _T_786; // @[Monitor.scala 541:29:freechips.rocketchip.system.DefaultRV32Config.fir@101008.6]
  wire  _T_788; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@101010.6]
  wire  _T_789; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@101011.6]
  wire  _T_790; // @[Monitor.scala 542:29:freechips.rocketchip.system.DefaultRV32Config.fir@101016.6]
  wire  _T_792; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@101018.6]
  wire  _T_793; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@101019.6]
  wire  _T_794; // @[Monitor.scala 543:29:freechips.rocketchip.system.DefaultRV32Config.fir@101024.6]
  wire  _T_796; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@101026.6]
  wire  _T_797; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@101027.6]
  wire  _T_798; // @[Monitor.scala 544:29:freechips.rocketchip.system.DefaultRV32Config.fir@101032.6]
  wire  _T_800; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@101034.6]
  wire  _T_801; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@101035.6]
  wire  _T_803; // @[Monitor.scala 546:20:freechips.rocketchip.system.DefaultRV32Config.fir@101042.4]
  reg  inflight; // @[Monitor.scala 608:27:freechips.rocketchip.system.DefaultRV32Config.fir@101051.4]
  reg [3:0] inflight_opcodes; // @[Monitor.scala 610:35:freechips.rocketchip.system.DefaultRV32Config.fir@101052.4]
  reg [3:0] inflight_sizes; // @[Monitor.scala 612:33:freechips.rocketchip.system.DefaultRV32Config.fir@101053.4]
  reg  _T_813; // @[Edges.scala 230:27:freechips.rocketchip.system.DefaultRV32Config.fir@101063.4]
  wire  _T_815; // @[Edges.scala 231:28:freechips.rocketchip.system.DefaultRV32Config.fir@101065.4]
  wire  a_first; // @[Edges.scala 232:25:freechips.rocketchip.system.DefaultRV32Config.fir@101066.4]
  reg  _T_831; // @[Edges.scala 230:27:freechips.rocketchip.system.DefaultRV32Config.fir@101085.4]
  wire  _T_833; // @[Edges.scala 231:28:freechips.rocketchip.system.DefaultRV32Config.fir@101087.4]
  wire  d_first; // @[Edges.scala 232:25:freechips.rocketchip.system.DefaultRV32Config.fir@101088.4]
  wire [2:0] _GEN_56; // @[Monitor.scala 629:69:freechips.rocketchip.system.DefaultRV32Config.fir@101107.4]
  wire [3:0] _T_841; // @[Monitor.scala 629:69:freechips.rocketchip.system.DefaultRV32Config.fir@101107.4]
  wire [3:0] _T_842; // @[Monitor.scala 629:44:freechips.rocketchip.system.DefaultRV32Config.fir@101108.4]
  wire [15:0] _T_846; // @[Monitor.scala 606:57:freechips.rocketchip.system.DefaultRV32Config.fir@101112.4]
  wire [15:0] _GEN_57; // @[Monitor.scala 629:97:freechips.rocketchip.system.DefaultRV32Config.fir@101113.4]
  wire [15:0] _T_847; // @[Monitor.scala 629:97:freechips.rocketchip.system.DefaultRV32Config.fir@101113.4]
  wire [15:0] _T_848; // @[Monitor.scala 629:152:freechips.rocketchip.system.DefaultRV32Config.fir@101114.4]
  wire [3:0] _T_850; // @[Monitor.scala 633:40:freechips.rocketchip.system.DefaultRV32Config.fir@101119.4]
  wire [15:0] _GEN_60; // @[Monitor.scala 633:91:freechips.rocketchip.system.DefaultRV32Config.fir@101124.4]
  wire [15:0] _T_855; // @[Monitor.scala 633:91:freechips.rocketchip.system.DefaultRV32Config.fir@101124.4]
  wire [15:0] _T_856; // @[Monitor.scala 633:144:freechips.rocketchip.system.DefaultRV32Config.fir@101125.4]
  wire  _T_860; // @[Monitor.scala 643:27:freechips.rocketchip.system.DefaultRV32Config.fir@101150.4]
  wire [3:0] _T_863; // @[Monitor.scala 645:53:freechips.rocketchip.system.DefaultRV32Config.fir@101155.6]
  wire [3:0] _T_864; // @[Monitor.scala 645:61:freechips.rocketchip.system.DefaultRV32Config.fir@101156.6]
  wire [3:0] a_opcodes_set_interm; // @[Monitor.scala 643:72:freechips.rocketchip.system.DefaultRV32Config.fir@101152.4]
  wire [18:0] _T_868; // @[Monitor.scala 647:47:freechips.rocketchip.system.DefaultRV32Config.fir@101162.6]
  wire [2:0] a_sizes_set_interm; // @[Monitor.scala 643:72:freechips.rocketchip.system.DefaultRV32Config.fir@101152.4]
  wire [17:0] _T_870; // @[Monitor.scala 648:43:freechips.rocketchip.system.DefaultRV32Config.fir@101165.6]
  wire  _T_873; // @[Monitor.scala 649:17:freechips.rocketchip.system.DefaultRV32Config.fir@101169.6]
  wire  _T_875; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@101171.6]
  wire  _T_876; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@101172.6]
  wire [1:0] _GEN_15; // @[Monitor.scala 643:72:freechips.rocketchip.system.DefaultRV32Config.fir@101152.4]
  wire [18:0] _GEN_18; // @[Monitor.scala 643:72:freechips.rocketchip.system.DefaultRV32Config.fir@101152.4]
  wire [17:0] _GEN_19; // @[Monitor.scala 643:72:freechips.rocketchip.system.DefaultRV32Config.fir@101152.4]
  wire  _T_879; // @[Monitor.scala 660:27:freechips.rocketchip.system.DefaultRV32Config.fir@101186.4]
  wire  _T_881; // @[Monitor.scala 660:75:freechips.rocketchip.system.DefaultRV32Config.fir@101188.4]
  wire  _T_882; // @[Monitor.scala 660:72:freechips.rocketchip.system.DefaultRV32Config.fir@101189.4]
  wire [1:0] _T_883; // @[OneHot.scala 58:35:freechips.rocketchip.system.DefaultRV32Config.fir@101191.6]
  wire [30:0] _GEN_63; // @[Monitor.scala 662:76:freechips.rocketchip.system.DefaultRV32Config.fir@101198.6]
  wire [30:0] _T_889; // @[Monitor.scala 662:76:freechips.rocketchip.system.DefaultRV32Config.fir@101198.6]
  wire [1:0] _GEN_20; // @[Monitor.scala 660:91:freechips.rocketchip.system.DefaultRV32Config.fir@101190.4]
  wire [30:0] _GEN_21; // @[Monitor.scala 660:91:freechips.rocketchip.system.DefaultRV32Config.fir@101190.4]
  wire  _T_896; // @[Monitor.scala 665:26:freechips.rocketchip.system.DefaultRV32Config.fir@101208.4]
  wire  _T_899; // @[Monitor.scala 665:71:freechips.rocketchip.system.DefaultRV32Config.fir@101211.4]
  wire  _T_900; // @[Monitor.scala 666:25:freechips.rocketchip.system.DefaultRV32Config.fir@101213.6]
  wire  _T_903; // @[Monitor.scala 666:68:freechips.rocketchip.system.DefaultRV32Config.fir@101216.6]
  wire  _T_904; // @[Monitor.scala 666:142:freechips.rocketchip.system.DefaultRV32Config.fir@101217.6]
  wire  _T_905; // @[Monitor.scala 666:119:freechips.rocketchip.system.DefaultRV32Config.fir@101218.6]
  wire  _T_906; // @[Monitor.scala 666:166:freechips.rocketchip.system.DefaultRV32Config.fir@101219.6]
  wire  _T_907; // @[Monitor.scala 666:49:freechips.rocketchip.system.DefaultRV32Config.fir@101220.6]
  wire  _T_909; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@101222.6]
  wire  _T_910; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@101223.6]
  wire [3:0] a_opcode_lookup; // @[:freechips.rocketchip.system.DefaultRV32Config.fir@101105.4 :freechips.rocketchip.system.DefaultRV32Config.fir@101106.4 Monitor.scala 629:21:freechips.rocketchip.system.DefaultRV32Config.fir@101115.4]
  wire [2:0] _GEN_25; // @[Monitor.scala 667:37:freechips.rocketchip.system.DefaultRV32Config.fir@101229.6]
  wire [2:0] _GEN_26; // @[Monitor.scala 667:37:freechips.rocketchip.system.DefaultRV32Config.fir@101229.6]
  wire [2:0] _GEN_27; // @[Monitor.scala 667:37:freechips.rocketchip.system.DefaultRV32Config.fir@101229.6]
  wire [2:0] _GEN_28; // @[Monitor.scala 667:37:freechips.rocketchip.system.DefaultRV32Config.fir@101229.6]
  wire [2:0] _GEN_29; // @[Monitor.scala 667:37:freechips.rocketchip.system.DefaultRV32Config.fir@101229.6]
  wire [2:0] _GEN_30; // @[Monitor.scala 667:37:freechips.rocketchip.system.DefaultRV32Config.fir@101229.6]
  wire  _T_912; // @[Monitor.scala 667:37:freechips.rocketchip.system.DefaultRV32Config.fir@101229.6]
  wire [2:0] _GEN_37; // @[Monitor.scala 667:96:freechips.rocketchip.system.DefaultRV32Config.fir@101231.6]
  wire [2:0] _GEN_38; // @[Monitor.scala 667:96:freechips.rocketchip.system.DefaultRV32Config.fir@101231.6]
  wire  _T_914; // @[Monitor.scala 667:96:freechips.rocketchip.system.DefaultRV32Config.fir@101231.6]
  wire  _T_915; // @[Monitor.scala 667:71:freechips.rocketchip.system.DefaultRV32Config.fir@101232.6]
  wire [2:0] _GEN_41; // @[Monitor.scala 668:60:freechips.rocketchip.system.DefaultRV32Config.fir@101233.6]
  wire [2:0] _GEN_42; // @[Monitor.scala 668:60:freechips.rocketchip.system.DefaultRV32Config.fir@101233.6]
  wire [2:0] _GEN_43; // @[Monitor.scala 668:60:freechips.rocketchip.system.DefaultRV32Config.fir@101233.6]
  wire [2:0] _GEN_44; // @[Monitor.scala 668:60:freechips.rocketchip.system.DefaultRV32Config.fir@101233.6]
  wire [2:0] _GEN_45; // @[Monitor.scala 668:60:freechips.rocketchip.system.DefaultRV32Config.fir@101233.6]
  wire [2:0] _GEN_46; // @[Monitor.scala 668:60:freechips.rocketchip.system.DefaultRV32Config.fir@101233.6]
  wire  _T_916; // @[Monitor.scala 668:60:freechips.rocketchip.system.DefaultRV32Config.fir@101233.6]
  wire [2:0] _GEN_53; // @[Monitor.scala 668:124:freechips.rocketchip.system.DefaultRV32Config.fir@101234.6]
  wire [2:0] _GEN_54; // @[Monitor.scala 668:124:freechips.rocketchip.system.DefaultRV32Config.fir@101234.6]
  wire  _T_917; // @[Monitor.scala 668:124:freechips.rocketchip.system.DefaultRV32Config.fir@101234.6]
  wire  _T_918; // @[Monitor.scala 668:99:freechips.rocketchip.system.DefaultRV32Config.fir@101235.6]
  wire  _T_919; // @[Monitor.scala 668:34:freechips.rocketchip.system.DefaultRV32Config.fir@101236.6]
  wire  _T_920; // @[Monitor.scala 668:15:freechips.rocketchip.system.DefaultRV32Config.fir@101237.6]
  wire  _T_922; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@101239.6]
  wire  _T_923; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@101240.6]
  wire [3:0] a_size_lookup; // @[:freechips.rocketchip.system.DefaultRV32Config.fir@101116.4 :freechips.rocketchip.system.DefaultRV32Config.fir@101117.4 Monitor.scala 633:19:freechips.rocketchip.system.DefaultRV32Config.fir@101126.4]
  wire [3:0] _GEN_66; // @[Monitor.scala 670:34:freechips.rocketchip.system.DefaultRV32Config.fir@101245.6]
  wire  _T_924; // @[Monitor.scala 670:34:freechips.rocketchip.system.DefaultRV32Config.fir@101245.6]
  wire  _T_926; // @[Monitor.scala 670:72:freechips.rocketchip.system.DefaultRV32Config.fir@101247.6]
  wire  _T_927; // @[Monitor.scala 670:53:freechips.rocketchip.system.DefaultRV32Config.fir@101248.6]
  wire  _T_929; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@101250.6]
  wire  _T_930; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@101251.6]
  wire  _T_932; // @[Monitor.scala 672:36:freechips.rocketchip.system.DefaultRV32Config.fir@101258.4]
  wire  _T_933; // @[Monitor.scala 672:47:freechips.rocketchip.system.DefaultRV32Config.fir@101259.4]
  wire  _T_935; // @[Monitor.scala 672:65:freechips.rocketchip.system.DefaultRV32Config.fir@101261.4]
  wire  _T_937; // @[Monitor.scala 672:116:freechips.rocketchip.system.DefaultRV32Config.fir@101263.4]
  wire  _T_938; // @[Monitor.scala 673:15:freechips.rocketchip.system.DefaultRV32Config.fir@101265.6]
  wire  _T_939; // @[Monitor.scala 673:32:freechips.rocketchip.system.DefaultRV32Config.fir@101266.6]
  wire  _T_941; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@101268.6]
  wire  _T_942; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@101269.6]
  wire  a_set; // @[:freechips.rocketchip.system.DefaultRV32Config.fir@101099.4 :freechips.rocketchip.system.DefaultRV32Config.fir@101100.4 Monitor.scala 644:13:freechips.rocketchip.system.DefaultRV32Config.fir@101154.6]
  wire  _T_943; // @[Monitor.scala 680:27:freechips.rocketchip.system.DefaultRV32Config.fir@101275.4]
  wire  d_clr; // @[:freechips.rocketchip.system.DefaultRV32Config.fir@101178.4 :freechips.rocketchip.system.DefaultRV32Config.fir@101179.4 Monitor.scala 661:13:freechips.rocketchip.system.DefaultRV32Config.fir@101192.6]
  wire  _T_944; // @[Monitor.scala 680:38:freechips.rocketchip.system.DefaultRV32Config.fir@101276.4]
  wire  _T_945; // @[Monitor.scala 680:36:freechips.rocketchip.system.DefaultRV32Config.fir@101277.4]
  wire [3:0] a_opcodes_set; // @[:freechips.rocketchip.system.DefaultRV32Config.fir@101101.4 :freechips.rocketchip.system.DefaultRV32Config.fir@101102.4 Monitor.scala 647:21:freechips.rocketchip.system.DefaultRV32Config.fir@101163.6]
  wire [3:0] _T_946; // @[Monitor.scala 681:43:freechips.rocketchip.system.DefaultRV32Config.fir@101279.4]
  wire [3:0] d_opcodes_clr; // @[:freechips.rocketchip.system.DefaultRV32Config.fir@101180.4 :freechips.rocketchip.system.DefaultRV32Config.fir@101181.4 Monitor.scala 662:21:freechips.rocketchip.system.DefaultRV32Config.fir@101199.6]
  wire [3:0] _T_947; // @[Monitor.scala 681:62:freechips.rocketchip.system.DefaultRV32Config.fir@101280.4]
  wire [3:0] _T_948; // @[Monitor.scala 681:60:freechips.rocketchip.system.DefaultRV32Config.fir@101281.4]
  wire [3:0] a_sizes_set; // @[:freechips.rocketchip.system.DefaultRV32Config.fir@101103.4 :freechips.rocketchip.system.DefaultRV32Config.fir@101104.4 Monitor.scala 648:19:freechips.rocketchip.system.DefaultRV32Config.fir@101166.6]
  wire [3:0] _T_949; // @[Monitor.scala 682:39:freechips.rocketchip.system.DefaultRV32Config.fir@101283.4]
  wire [3:0] _T_951; // @[Monitor.scala 682:54:freechips.rocketchip.system.DefaultRV32Config.fir@101285.4]
  reg [31:0] _T_952; // @[Monitor.scala 684:27:freechips.rocketchip.system.DefaultRV32Config.fir@101287.4]
  wire  _T_953; // @[Monitor.scala 687:26:freechips.rocketchip.system.DefaultRV32Config.fir@101290.4]
  wire  _T_954; // @[Monitor.scala 687:16:freechips.rocketchip.system.DefaultRV32Config.fir@101291.4]
  wire  _T_955; // @[Monitor.scala 687:39:freechips.rocketchip.system.DefaultRV32Config.fir@101292.4]
  wire  _T_956; // @[Monitor.scala 687:30:freechips.rocketchip.system.DefaultRV32Config.fir@101293.4]
  wire  _T_957; // @[Monitor.scala 687:59:freechips.rocketchip.system.DefaultRV32Config.fir@101294.4]
  wire  _T_958; // @[Monitor.scala 687:47:freechips.rocketchip.system.DefaultRV32Config.fir@101295.4]
  wire  _T_960; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@101297.4]
  wire  _T_961; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@101298.4]
  wire [31:0] _T_963; // @[Monitor.scala 689:26:freechips.rocketchip.system.DefaultRV32Config.fir@101304.4]
  wire  _T_966; // @[Monitor.scala 690:27:freechips.rocketchip.system.DefaultRV32Config.fir@101308.4]
  wire  _GEN_67; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@99906.10]
  wire  _GEN_75; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@100008.10]
  wire  _GEN_85; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@100121.10]
  wire  _GEN_91; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@100210.10]
  wire  _GEN_97; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@100291.10]
  wire  _GEN_101; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@100371.10]
  wire  _GEN_107; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@100449.10]
  wire  _GEN_113; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@100527.10]
  wire  _GEN_119; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@100590.10]
  wire  _GEN_129; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@100632.10]
  wire  _GEN_141; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@100690.10]
  wire  _GEN_153; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@100749.10]
  wire  _GEN_159; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@100784.10]
  wire  _GEN_165; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@100820.10]
  plusarg_reader #(.FORMAT("tilelink_timeout=%d"), .DEFAULT(0), .WIDTH(32)) plusarg_reader ( // @[PlusArg.scala 80:11:freechips.rocketchip.system.DefaultRV32Config.fir@101288.4]
    .out(plusarg_reader_out)
  );
  assign _T_10 = io_in_a_bits_address & 9'h3; // @[Edges.scala 22:16:freechips.rocketchip.system.DefaultRV32Config.fir@99812.6]
  assign _T_11 = _T_10 == 9'h0; // @[Edges.scala 22:24:freechips.rocketchip.system.DefaultRV32Config.fir@99813.6]
  assign _T_48 = {1'b0,$signed(io_in_a_bits_address)}; // @[Parameters.scala 137:49:freechips.rocketchip.system.DefaultRV32Config.fir@99850.6]
  assign _T_56 = io_in_a_bits_opcode == 3'h6; // @[Monitor.scala 79:25:freechips.rocketchip.system.DefaultRV32Config.fir@99862.6]
  assign _T_61 = $signed(_T_48) & -10'sh40; // @[Parameters.scala 137:52:freechips.rocketchip.system.DefaultRV32Config.fir@99868.8]
  assign _T_62 = $signed(_T_61) == 10'sh0; // @[Parameters.scala 137:67:freechips.rocketchip.system.DefaultRV32Config.fir@99869.8]
  assign _T_63 = io_in_a_bits_address ^ 9'h44; // @[Parameters.scala 137:31:freechips.rocketchip.system.DefaultRV32Config.fir@99870.8]
  assign _T_64 = {1'b0,$signed(_T_63)}; // @[Parameters.scala 137:49:freechips.rocketchip.system.DefaultRV32Config.fir@99871.8]
  assign _T_66 = $signed(_T_64) & -10'sh4; // @[Parameters.scala 137:52:freechips.rocketchip.system.DefaultRV32Config.fir@99873.8]
  assign _T_67 = $signed(_T_66) == 10'sh0; // @[Parameters.scala 137:67:freechips.rocketchip.system.DefaultRV32Config.fir@99874.8]
  assign _T_68 = io_in_a_bits_address ^ 9'h48; // @[Parameters.scala 137:31:freechips.rocketchip.system.DefaultRV32Config.fir@99875.8]
  assign _T_69 = {1'b0,$signed(_T_68)}; // @[Parameters.scala 137:49:freechips.rocketchip.system.DefaultRV32Config.fir@99876.8]
  assign _T_71 = $signed(_T_69) & -10'sh18; // @[Parameters.scala 137:52:freechips.rocketchip.system.DefaultRV32Config.fir@99878.8]
  assign _T_72 = $signed(_T_71) == 10'sh0; // @[Parameters.scala 137:67:freechips.rocketchip.system.DefaultRV32Config.fir@99879.8]
  assign _T_73 = io_in_a_bits_address ^ 9'h60; // @[Parameters.scala 137:31:freechips.rocketchip.system.DefaultRV32Config.fir@99880.8]
  assign _T_74 = {1'b0,$signed(_T_73)}; // @[Parameters.scala 137:49:freechips.rocketchip.system.DefaultRV32Config.fir@99881.8]
  assign _T_76 = $signed(_T_74) & -10'sh20; // @[Parameters.scala 137:52:freechips.rocketchip.system.DefaultRV32Config.fir@99883.8]
  assign _T_77 = $signed(_T_76) == 10'sh0; // @[Parameters.scala 137:67:freechips.rocketchip.system.DefaultRV32Config.fir@99884.8]
  assign _T_78 = io_in_a_bits_address ^ 9'h80; // @[Parameters.scala 137:31:freechips.rocketchip.system.DefaultRV32Config.fir@99885.8]
  assign _T_79 = {1'b0,$signed(_T_78)}; // @[Parameters.scala 137:49:freechips.rocketchip.system.DefaultRV32Config.fir@99886.8]
  assign _T_81 = $signed(_T_79) & -10'sh80; // @[Parameters.scala 137:52:freechips.rocketchip.system.DefaultRV32Config.fir@99888.8]
  assign _T_82 = $signed(_T_81) == 10'sh0; // @[Parameters.scala 137:67:freechips.rocketchip.system.DefaultRV32Config.fir@99889.8]
  assign _T_83 = io_in_a_bits_address ^ 9'h100; // @[Parameters.scala 137:31:freechips.rocketchip.system.DefaultRV32Config.fir@99890.8]
  assign _T_84 = {1'b0,$signed(_T_83)}; // @[Parameters.scala 137:49:freechips.rocketchip.system.DefaultRV32Config.fir@99891.8]
  assign _T_86 = $signed(_T_84) & -10'sh100; // @[Parameters.scala 137:52:freechips.rocketchip.system.DefaultRV32Config.fir@99893.8]
  assign _T_87 = $signed(_T_86) == 10'sh0; // @[Parameters.scala 137:67:freechips.rocketchip.system.DefaultRV32Config.fir@99894.8]
  assign _T_88 = _T_62 | _T_67; // @[Parameters.scala 552:42:freechips.rocketchip.system.DefaultRV32Config.fir@99895.8]
  assign _T_89 = _T_88 | _T_72; // @[Parameters.scala 552:42:freechips.rocketchip.system.DefaultRV32Config.fir@99896.8]
  assign _T_90 = _T_89 | _T_77; // @[Parameters.scala 552:42:freechips.rocketchip.system.DefaultRV32Config.fir@99897.8]
  assign _T_91 = _T_90 | _T_82; // @[Parameters.scala 552:42:freechips.rocketchip.system.DefaultRV32Config.fir@99898.8]
  assign _T_92 = _T_91 | _T_87; // @[Parameters.scala 552:42:freechips.rocketchip.system.DefaultRV32Config.fir@99899.8]
  assign _T_97 = ~reset; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@99904.8]
  assign _T_109 = _T_11 | reset; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@99932.8]
  assign _T_110 = ~_T_109; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@99933.8]
  assign _T_115 = ~io_in_a_bits_mask; // @[Monitor.scala 86:18:freechips.rocketchip.system.DefaultRV32Config.fir@99946.8]
  assign _T_116 = _T_115 == 4'h0; // @[Monitor.scala 86:31:freechips.rocketchip.system.DefaultRV32Config.fir@99947.8]
  assign _T_118 = _T_116 | reset; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@99949.8]
  assign _T_119 = ~_T_118; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@99950.8]
  assign _T_124 = io_in_a_bits_opcode == 3'h7; // @[Monitor.scala 90:25:freechips.rocketchip.system.DefaultRV32Config.fir@99964.6]
  assign _T_196 = io_in_a_bits_opcode == 3'h4; // @[Monitor.scala 102:25:freechips.rocketchip.system.DefaultRV32Config.fir@100074.6]
  assign _T_239 = _T_92 | reset; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@100118.8]
  assign _T_240 = ~_T_239; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@100119.8]
  assign _T_251 = io_in_a_bits_mask == 4'hf; // @[Monitor.scala 107:30:freechips.rocketchip.system.DefaultRV32Config.fir@100146.8]
  assign _T_253 = _T_251 | reset; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@100148.8]
  assign _T_254 = ~_T_253; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@100149.8]
  assign _T_259 = io_in_a_bits_opcode == 3'h0; // @[Monitor.scala 111:25:freechips.rocketchip.system.DefaultRV32Config.fir@100163.6]
  assign _T_318 = io_in_a_bits_opcode == 3'h1; // @[Monitor.scala 119:25:freechips.rocketchip.system.DefaultRV32Config.fir@100244.6]
  assign _T_379 = io_in_a_bits_opcode == 3'h2; // @[Monitor.scala 127:25:freechips.rocketchip.system.DefaultRV32Config.fir@100327.6]
  assign _T_435 = io_in_a_bits_opcode == 3'h3; // @[Monitor.scala 135:25:freechips.rocketchip.system.DefaultRV32Config.fir@100405.6]
  assign _T_491 = io_in_a_bits_opcode == 3'h5; // @[Monitor.scala 143:25:freechips.rocketchip.system.DefaultRV32Config.fir@100483.6]
  assign _T_551 = io_in_d_bits_opcode <= 3'h6; // @[Bundles.scala 44:24:freechips.rocketchip.system.DefaultRV32Config.fir@100571.6]
  assign _T_553 = _T_551 | reset; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@100573.6]
  assign _T_554 = ~_T_553; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@100574.6]
  assign _T_555 = ~io_in_d_bits_source; // @[Parameters.scala 47:9:freechips.rocketchip.system.DefaultRV32Config.fir@100579.6]
  assign _T_558 = io_in_d_bits_opcode == 3'h6; // @[Monitor.scala 307:25:freechips.rocketchip.system.DefaultRV32Config.fir@100584.6]
  assign _T_560 = _T_555 | reset; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@100587.8]
  assign _T_561 = ~_T_560; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@100588.8]
  assign _T_562 = io_in_d_bits_size >= 2'h2; // @[Monitor.scala 309:27:freechips.rocketchip.system.DefaultRV32Config.fir@100593.8]
  assign _T_564 = _T_562 | reset; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@100595.8]
  assign _T_565 = ~_T_564; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@100596.8]
  assign _T_566 = io_in_d_bits_param == 2'h0; // @[Monitor.scala 310:28:freechips.rocketchip.system.DefaultRV32Config.fir@100601.8]
  assign _T_568 = _T_566 | reset; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@100603.8]
  assign _T_569 = ~_T_568; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@100604.8]
  assign _T_570 = ~io_in_d_bits_corrupt; // @[Monitor.scala 311:15:freechips.rocketchip.system.DefaultRV32Config.fir@100609.8]
  assign _T_572 = _T_570 | reset; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@100611.8]
  assign _T_573 = ~_T_572; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@100612.8]
  assign _T_574 = ~io_in_d_bits_denied; // @[Monitor.scala 312:15:freechips.rocketchip.system.DefaultRV32Config.fir@100617.8]
  assign _T_576 = _T_574 | reset; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@100619.8]
  assign _T_577 = ~_T_576; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@100620.8]
  assign _T_578 = io_in_d_bits_opcode == 3'h4; // @[Monitor.scala 315:25:freechips.rocketchip.system.DefaultRV32Config.fir@100626.6]
  assign _T_589 = io_in_d_bits_param <= 2'h2; // @[Bundles.scala 104:26:freechips.rocketchip.system.DefaultRV32Config.fir@100650.8]
  assign _T_591 = _T_589 | reset; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@100652.8]
  assign _T_592 = ~_T_591; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@100653.8]
  assign _T_593 = io_in_d_bits_param != 2'h2; // @[Monitor.scala 320:28:freechips.rocketchip.system.DefaultRV32Config.fir@100658.8]
  assign _T_595 = _T_593 | reset; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@100660.8]
  assign _T_596 = ~_T_595; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@100661.8]
  assign _T_606 = io_in_d_bits_opcode == 3'h5; // @[Monitor.scala 325:25:freechips.rocketchip.system.DefaultRV32Config.fir@100684.6]
  assign _T_626 = _T_574 | io_in_d_bits_corrupt; // @[Monitor.scala 331:30:freechips.rocketchip.system.DefaultRV32Config.fir@100725.8]
  assign _T_628 = _T_626 | reset; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@100727.8]
  assign _T_629 = ~_T_628; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@100728.8]
  assign _T_635 = io_in_d_bits_opcode == 3'h0; // @[Monitor.scala 335:25:freechips.rocketchip.system.DefaultRV32Config.fir@100743.6]
  assign _T_652 = io_in_d_bits_opcode == 3'h1; // @[Monitor.scala 343:25:freechips.rocketchip.system.DefaultRV32Config.fir@100778.6]
  assign _T_670 = io_in_d_bits_opcode == 3'h2; // @[Monitor.scala 351:25:freechips.rocketchip.system.DefaultRV32Config.fir@100814.6]
  assign _T_702 = io_in_a_ready & io_in_a_valid; // @[Decoupled.scala 40:37:freechips.rocketchip.system.DefaultRV32Config.fir@100880.4]
  assign _T_713 = _T_711 - 1'h1; // @[Edges.scala 231:28:freechips.rocketchip.system.DefaultRV32Config.fir@100891.4]
  assign _T_714 = ~_T_711; // @[Edges.scala 232:25:freechips.rocketchip.system.DefaultRV32Config.fir@100892.4]
  assign _T_727 = ~_T_714; // @[Monitor.scala 386:22:freechips.rocketchip.system.DefaultRV32Config.fir@100908.4]
  assign _T_728 = io_in_a_valid & _T_727; // @[Monitor.scala 386:19:freechips.rocketchip.system.DefaultRV32Config.fir@100909.4]
  assign _T_729 = io_in_a_bits_opcode == _T_722; // @[Monitor.scala 387:32:freechips.rocketchip.system.DefaultRV32Config.fir@100911.6]
  assign _T_731 = _T_729 | reset; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@100913.6]
  assign _T_732 = ~_T_731; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@100914.6]
  assign _T_745 = io_in_a_bits_address == _T_726; // @[Monitor.scala 391:32:freechips.rocketchip.system.DefaultRV32Config.fir@100943.6]
  assign _T_747 = _T_745 | reset; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@100945.6]
  assign _T_748 = ~_T_747; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@100946.6]
  assign _T_750 = _T_702 & _T_714; // @[Monitor.scala 393:20:freechips.rocketchip.system.DefaultRV32Config.fir@100953.4]
  assign _T_751 = io_in_d_ready & io_in_d_valid; // @[Decoupled.scala 40:37:freechips.rocketchip.system.DefaultRV32Config.fir@100961.4]
  assign _T_761 = _T_759 - 1'h1; // @[Edges.scala 231:28:freechips.rocketchip.system.DefaultRV32Config.fir@100971.4]
  assign _T_762 = ~_T_759; // @[Edges.scala 232:25:freechips.rocketchip.system.DefaultRV32Config.fir@100972.4]
  assign _T_776 = ~_T_762; // @[Monitor.scala 538:22:freechips.rocketchip.system.DefaultRV32Config.fir@100989.4]
  assign _T_777 = io_in_d_valid & _T_776; // @[Monitor.scala 538:19:freechips.rocketchip.system.DefaultRV32Config.fir@100990.4]
  assign _T_778 = io_in_d_bits_opcode == _T_770; // @[Monitor.scala 539:29:freechips.rocketchip.system.DefaultRV32Config.fir@100992.6]
  assign _T_780 = _T_778 | reset; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@100994.6]
  assign _T_781 = ~_T_780; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@100995.6]
  assign _T_782 = io_in_d_bits_param == _T_771; // @[Monitor.scala 540:29:freechips.rocketchip.system.DefaultRV32Config.fir@101000.6]
  assign _T_784 = _T_782 | reset; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@101002.6]
  assign _T_785 = ~_T_784; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@101003.6]
  assign _T_786 = io_in_d_bits_size == _T_772; // @[Monitor.scala 541:29:freechips.rocketchip.system.DefaultRV32Config.fir@101008.6]
  assign _T_788 = _T_786 | reset; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@101010.6]
  assign _T_789 = ~_T_788; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@101011.6]
  assign _T_790 = io_in_d_bits_source == _T_773; // @[Monitor.scala 542:29:freechips.rocketchip.system.DefaultRV32Config.fir@101016.6]
  assign _T_792 = _T_790 | reset; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@101018.6]
  assign _T_793 = ~_T_792; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@101019.6]
  assign _T_794 = io_in_d_bits_sink == _T_774; // @[Monitor.scala 543:29:freechips.rocketchip.system.DefaultRV32Config.fir@101024.6]
  assign _T_796 = _T_794 | reset; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@101026.6]
  assign _T_797 = ~_T_796; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@101027.6]
  assign _T_798 = io_in_d_bits_denied == _T_775; // @[Monitor.scala 544:29:freechips.rocketchip.system.DefaultRV32Config.fir@101032.6]
  assign _T_800 = _T_798 | reset; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@101034.6]
  assign _T_801 = ~_T_800; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@101035.6]
  assign _T_803 = _T_751 & _T_762; // @[Monitor.scala 546:20:freechips.rocketchip.system.DefaultRV32Config.fir@101042.4]
  assign _T_815 = _T_813 - 1'h1; // @[Edges.scala 231:28:freechips.rocketchip.system.DefaultRV32Config.fir@101065.4]
  assign a_first = ~_T_813; // @[Edges.scala 232:25:freechips.rocketchip.system.DefaultRV32Config.fir@101066.4]
  assign _T_833 = _T_831 - 1'h1; // @[Edges.scala 231:28:freechips.rocketchip.system.DefaultRV32Config.fir@101087.4]
  assign d_first = ~_T_831; // @[Edges.scala 232:25:freechips.rocketchip.system.DefaultRV32Config.fir@101088.4]
  assign _GEN_56 = {io_in_d_bits_source, 2'h0}; // @[Monitor.scala 629:69:freechips.rocketchip.system.DefaultRV32Config.fir@101107.4]
  assign _T_841 = {{1'd0}, _GEN_56}; // @[Monitor.scala 629:69:freechips.rocketchip.system.DefaultRV32Config.fir@101107.4]
  assign _T_842 = inflight_opcodes >> _T_841; // @[Monitor.scala 629:44:freechips.rocketchip.system.DefaultRV32Config.fir@101108.4]
  assign _T_846 = 16'h10 - 16'h1; // @[Monitor.scala 606:57:freechips.rocketchip.system.DefaultRV32Config.fir@101112.4]
  assign _GEN_57 = {{12'd0}, _T_842}; // @[Monitor.scala 629:97:freechips.rocketchip.system.DefaultRV32Config.fir@101113.4]
  assign _T_847 = _GEN_57 & _T_846; // @[Monitor.scala 629:97:freechips.rocketchip.system.DefaultRV32Config.fir@101113.4]
  assign _T_848 = {{1'd0}, _T_847[15:1]}; // @[Monitor.scala 629:152:freechips.rocketchip.system.DefaultRV32Config.fir@101114.4]
  assign _T_850 = inflight_sizes >> _T_841; // @[Monitor.scala 633:40:freechips.rocketchip.system.DefaultRV32Config.fir@101119.4]
  assign _GEN_60 = {{12'd0}, _T_850}; // @[Monitor.scala 633:91:freechips.rocketchip.system.DefaultRV32Config.fir@101124.4]
  assign _T_855 = _GEN_60 & _T_846; // @[Monitor.scala 633:91:freechips.rocketchip.system.DefaultRV32Config.fir@101124.4]
  assign _T_856 = {{1'd0}, _T_855[15:1]}; // @[Monitor.scala 633:144:freechips.rocketchip.system.DefaultRV32Config.fir@101125.4]
  assign _T_860 = _T_702 & a_first; // @[Monitor.scala 643:27:freechips.rocketchip.system.DefaultRV32Config.fir@101150.4]
  assign _T_863 = {io_in_a_bits_opcode, 1'h0}; // @[Monitor.scala 645:53:freechips.rocketchip.system.DefaultRV32Config.fir@101155.6]
  assign _T_864 = _T_863 | 4'h1; // @[Monitor.scala 645:61:freechips.rocketchip.system.DefaultRV32Config.fir@101156.6]
  assign a_opcodes_set_interm = _T_860 ? _T_864 : 4'h0; // @[Monitor.scala 643:72:freechips.rocketchip.system.DefaultRV32Config.fir@101152.4]
  assign _T_868 = {{15'd0}, a_opcodes_set_interm}; // @[Monitor.scala 647:47:freechips.rocketchip.system.DefaultRV32Config.fir@101162.6]
  assign a_sizes_set_interm = _T_860 ? 3'h5 : 3'h0; // @[Monitor.scala 643:72:freechips.rocketchip.system.DefaultRV32Config.fir@101152.4]
  assign _T_870 = {{15'd0}, a_sizes_set_interm}; // @[Monitor.scala 648:43:freechips.rocketchip.system.DefaultRV32Config.fir@101165.6]
  assign _T_873 = ~inflight; // @[Monitor.scala 649:17:freechips.rocketchip.system.DefaultRV32Config.fir@101169.6]
  assign _T_875 = _T_873 | reset; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@101171.6]
  assign _T_876 = ~_T_875; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@101172.6]
  assign _GEN_15 = _T_860 ? 2'h1 : 2'h0; // @[Monitor.scala 643:72:freechips.rocketchip.system.DefaultRV32Config.fir@101152.4]
  assign _GEN_18 = _T_860 ? _T_868 : 19'h0; // @[Monitor.scala 643:72:freechips.rocketchip.system.DefaultRV32Config.fir@101152.4]
  assign _GEN_19 = _T_860 ? _T_870 : 18'h0; // @[Monitor.scala 643:72:freechips.rocketchip.system.DefaultRV32Config.fir@101152.4]
  assign _T_879 = _T_751 & d_first; // @[Monitor.scala 660:27:freechips.rocketchip.system.DefaultRV32Config.fir@101186.4]
  assign _T_881 = ~_T_558; // @[Monitor.scala 660:75:freechips.rocketchip.system.DefaultRV32Config.fir@101188.4]
  assign _T_882 = _T_879 & _T_881; // @[Monitor.scala 660:72:freechips.rocketchip.system.DefaultRV32Config.fir@101189.4]
  assign _T_883 = 2'h1 << io_in_d_bits_source; // @[OneHot.scala 58:35:freechips.rocketchip.system.DefaultRV32Config.fir@101191.6]
  assign _GEN_63 = {{15'd0}, _T_846}; // @[Monitor.scala 662:76:freechips.rocketchip.system.DefaultRV32Config.fir@101198.6]
  assign _T_889 = _GEN_63 << _T_841; // @[Monitor.scala 662:76:freechips.rocketchip.system.DefaultRV32Config.fir@101198.6]
  assign _GEN_20 = _T_882 ? _T_883 : 2'h0; // @[Monitor.scala 660:91:freechips.rocketchip.system.DefaultRV32Config.fir@101190.4]
  assign _GEN_21 = _T_882 ? _T_889 : 31'h0; // @[Monitor.scala 660:91:freechips.rocketchip.system.DefaultRV32Config.fir@101190.4]
  assign _T_896 = io_in_d_valid & d_first; // @[Monitor.scala 665:26:freechips.rocketchip.system.DefaultRV32Config.fir@101208.4]
  assign _T_899 = _T_896 & _T_881; // @[Monitor.scala 665:71:freechips.rocketchip.system.DefaultRV32Config.fir@101211.4]
  assign _T_900 = inflight >> io_in_d_bits_source; // @[Monitor.scala 666:25:freechips.rocketchip.system.DefaultRV32Config.fir@101213.6]
  assign _T_903 = io_in_a_valid & _T_555; // @[Monitor.scala 666:68:freechips.rocketchip.system.DefaultRV32Config.fir@101216.6]
  assign _T_904 = 2'h2 == io_in_d_bits_size; // @[Monitor.scala 666:142:freechips.rocketchip.system.DefaultRV32Config.fir@101217.6]
  assign _T_905 = _T_903 & _T_904; // @[Monitor.scala 666:119:freechips.rocketchip.system.DefaultRV32Config.fir@101218.6]
  assign _T_906 = _T_905 & a_first; // @[Monitor.scala 666:166:freechips.rocketchip.system.DefaultRV32Config.fir@101219.6]
  assign _T_907 = _T_900 | _T_906; // @[Monitor.scala 666:49:freechips.rocketchip.system.DefaultRV32Config.fir@101220.6]
  assign _T_909 = _T_907 | reset; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@101222.6]
  assign _T_910 = ~_T_909; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@101223.6]
  assign a_opcode_lookup = _T_848[3:0]; // @[:freechips.rocketchip.system.DefaultRV32Config.fir@101105.4 :freechips.rocketchip.system.DefaultRV32Config.fir@101106.4 Monitor.scala 629:21:freechips.rocketchip.system.DefaultRV32Config.fir@101115.4]
  assign _GEN_25 = 3'h2 == a_opcode_lookup[2:0] ? 3'h1 : 3'h0; // @[Monitor.scala 667:37:freechips.rocketchip.system.DefaultRV32Config.fir@101229.6]
  assign _GEN_26 = 3'h3 == a_opcode_lookup[2:0] ? 3'h1 : _GEN_25; // @[Monitor.scala 667:37:freechips.rocketchip.system.DefaultRV32Config.fir@101229.6]
  assign _GEN_27 = 3'h4 == a_opcode_lookup[2:0] ? 3'h1 : _GEN_26; // @[Monitor.scala 667:37:freechips.rocketchip.system.DefaultRV32Config.fir@101229.6]
  assign _GEN_28 = 3'h5 == a_opcode_lookup[2:0] ? 3'h2 : _GEN_27; // @[Monitor.scala 667:37:freechips.rocketchip.system.DefaultRV32Config.fir@101229.6]
  assign _GEN_29 = 3'h6 == a_opcode_lookup[2:0] ? 3'h4 : _GEN_28; // @[Monitor.scala 667:37:freechips.rocketchip.system.DefaultRV32Config.fir@101229.6]
  assign _GEN_30 = 3'h7 == a_opcode_lookup[2:0] ? 3'h4 : _GEN_29; // @[Monitor.scala 667:37:freechips.rocketchip.system.DefaultRV32Config.fir@101229.6]
  assign _T_912 = io_in_d_bits_opcode == _GEN_30; // @[Monitor.scala 667:37:freechips.rocketchip.system.DefaultRV32Config.fir@101229.6]
  assign _GEN_37 = 3'h6 == a_opcode_lookup[2:0] ? 3'h5 : _GEN_28; // @[Monitor.scala 667:96:freechips.rocketchip.system.DefaultRV32Config.fir@101231.6]
  assign _GEN_38 = 3'h7 == a_opcode_lookup[2:0] ? 3'h4 : _GEN_37; // @[Monitor.scala 667:96:freechips.rocketchip.system.DefaultRV32Config.fir@101231.6]
  assign _T_914 = io_in_d_bits_opcode == _GEN_38; // @[Monitor.scala 667:96:freechips.rocketchip.system.DefaultRV32Config.fir@101231.6]
  assign _T_915 = _T_912 | _T_914; // @[Monitor.scala 667:71:freechips.rocketchip.system.DefaultRV32Config.fir@101232.6]
  assign _GEN_41 = 3'h2 == io_in_a_bits_opcode ? 3'h1 : 3'h0; // @[Monitor.scala 668:60:freechips.rocketchip.system.DefaultRV32Config.fir@101233.6]
  assign _GEN_42 = 3'h3 == io_in_a_bits_opcode ? 3'h1 : _GEN_41; // @[Monitor.scala 668:60:freechips.rocketchip.system.DefaultRV32Config.fir@101233.6]
  assign _GEN_43 = 3'h4 == io_in_a_bits_opcode ? 3'h1 : _GEN_42; // @[Monitor.scala 668:60:freechips.rocketchip.system.DefaultRV32Config.fir@101233.6]
  assign _GEN_44 = 3'h5 == io_in_a_bits_opcode ? 3'h2 : _GEN_43; // @[Monitor.scala 668:60:freechips.rocketchip.system.DefaultRV32Config.fir@101233.6]
  assign _GEN_45 = 3'h6 == io_in_a_bits_opcode ? 3'h4 : _GEN_44; // @[Monitor.scala 668:60:freechips.rocketchip.system.DefaultRV32Config.fir@101233.6]
  assign _GEN_46 = 3'h7 == io_in_a_bits_opcode ? 3'h4 : _GEN_45; // @[Monitor.scala 668:60:freechips.rocketchip.system.DefaultRV32Config.fir@101233.6]
  assign _T_916 = io_in_d_bits_opcode == _GEN_46; // @[Monitor.scala 668:60:freechips.rocketchip.system.DefaultRV32Config.fir@101233.6]
  assign _GEN_53 = 3'h6 == io_in_a_bits_opcode ? 3'h5 : _GEN_44; // @[Monitor.scala 668:124:freechips.rocketchip.system.DefaultRV32Config.fir@101234.6]
  assign _GEN_54 = 3'h7 == io_in_a_bits_opcode ? 3'h4 : _GEN_53; // @[Monitor.scala 668:124:freechips.rocketchip.system.DefaultRV32Config.fir@101234.6]
  assign _T_917 = io_in_d_bits_opcode == _GEN_54; // @[Monitor.scala 668:124:freechips.rocketchip.system.DefaultRV32Config.fir@101234.6]
  assign _T_918 = _T_916 | _T_917; // @[Monitor.scala 668:99:freechips.rocketchip.system.DefaultRV32Config.fir@101235.6]
  assign _T_919 = io_in_a_valid & _T_918; // @[Monitor.scala 668:34:freechips.rocketchip.system.DefaultRV32Config.fir@101236.6]
  assign _T_920 = _T_915 | _T_919; // @[Monitor.scala 668:15:freechips.rocketchip.system.DefaultRV32Config.fir@101237.6]
  assign _T_922 = _T_920 | reset; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@101239.6]
  assign _T_923 = ~_T_922; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@101240.6]
  assign a_size_lookup = _T_856[3:0]; // @[:freechips.rocketchip.system.DefaultRV32Config.fir@101116.4 :freechips.rocketchip.system.DefaultRV32Config.fir@101117.4 Monitor.scala 633:19:freechips.rocketchip.system.DefaultRV32Config.fir@101126.4]
  assign _GEN_66 = {{2'd0}, io_in_d_bits_size}; // @[Monitor.scala 670:34:freechips.rocketchip.system.DefaultRV32Config.fir@101245.6]
  assign _T_924 = _GEN_66 == a_size_lookup; // @[Monitor.scala 670:34:freechips.rocketchip.system.DefaultRV32Config.fir@101245.6]
  assign _T_926 = io_in_a_valid & _T_904; // @[Monitor.scala 670:72:freechips.rocketchip.system.DefaultRV32Config.fir@101247.6]
  assign _T_927 = _T_924 | _T_926; // @[Monitor.scala 670:53:freechips.rocketchip.system.DefaultRV32Config.fir@101248.6]
  assign _T_929 = _T_927 | reset; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@101250.6]
  assign _T_930 = ~_T_929; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@101251.6]
  assign _T_932 = _T_896 & a_first; // @[Monitor.scala 672:36:freechips.rocketchip.system.DefaultRV32Config.fir@101258.4]
  assign _T_933 = _T_932 & io_in_a_valid; // @[Monitor.scala 672:47:freechips.rocketchip.system.DefaultRV32Config.fir@101259.4]
  assign _T_935 = _T_933 & _T_555; // @[Monitor.scala 672:65:freechips.rocketchip.system.DefaultRV32Config.fir@101261.4]
  assign _T_937 = _T_935 & _T_881; // @[Monitor.scala 672:116:freechips.rocketchip.system.DefaultRV32Config.fir@101263.4]
  assign _T_938 = ~io_in_d_ready; // @[Monitor.scala 673:15:freechips.rocketchip.system.DefaultRV32Config.fir@101265.6]
  assign _T_939 = _T_938 | io_in_a_ready; // @[Monitor.scala 673:32:freechips.rocketchip.system.DefaultRV32Config.fir@101266.6]
  assign _T_941 = _T_939 | reset; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@101268.6]
  assign _T_942 = ~_T_941; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@101269.6]
  assign a_set = _GEN_15[0]; // @[:freechips.rocketchip.system.DefaultRV32Config.fir@101099.4 :freechips.rocketchip.system.DefaultRV32Config.fir@101100.4 Monitor.scala 644:13:freechips.rocketchip.system.DefaultRV32Config.fir@101154.6]
  assign _T_943 = inflight | a_set; // @[Monitor.scala 680:27:freechips.rocketchip.system.DefaultRV32Config.fir@101275.4]
  assign d_clr = _GEN_20[0]; // @[:freechips.rocketchip.system.DefaultRV32Config.fir@101178.4 :freechips.rocketchip.system.DefaultRV32Config.fir@101179.4 Monitor.scala 661:13:freechips.rocketchip.system.DefaultRV32Config.fir@101192.6]
  assign _T_944 = ~d_clr; // @[Monitor.scala 680:38:freechips.rocketchip.system.DefaultRV32Config.fir@101276.4]
  assign _T_945 = _T_943 & _T_944; // @[Monitor.scala 680:36:freechips.rocketchip.system.DefaultRV32Config.fir@101277.4]
  assign a_opcodes_set = _GEN_18[3:0]; // @[:freechips.rocketchip.system.DefaultRV32Config.fir@101101.4 :freechips.rocketchip.system.DefaultRV32Config.fir@101102.4 Monitor.scala 647:21:freechips.rocketchip.system.DefaultRV32Config.fir@101163.6]
  assign _T_946 = inflight_opcodes | a_opcodes_set; // @[Monitor.scala 681:43:freechips.rocketchip.system.DefaultRV32Config.fir@101279.4]
  assign d_opcodes_clr = _GEN_21[3:0]; // @[:freechips.rocketchip.system.DefaultRV32Config.fir@101180.4 :freechips.rocketchip.system.DefaultRV32Config.fir@101181.4 Monitor.scala 662:21:freechips.rocketchip.system.DefaultRV32Config.fir@101199.6]
  assign _T_947 = ~d_opcodes_clr; // @[Monitor.scala 681:62:freechips.rocketchip.system.DefaultRV32Config.fir@101280.4]
  assign _T_948 = _T_946 & _T_947; // @[Monitor.scala 681:60:freechips.rocketchip.system.DefaultRV32Config.fir@101281.4]
  assign a_sizes_set = _GEN_19[3:0]; // @[:freechips.rocketchip.system.DefaultRV32Config.fir@101103.4 :freechips.rocketchip.system.DefaultRV32Config.fir@101104.4 Monitor.scala 648:19:freechips.rocketchip.system.DefaultRV32Config.fir@101166.6]
  assign _T_949 = inflight_sizes | a_sizes_set; // @[Monitor.scala 682:39:freechips.rocketchip.system.DefaultRV32Config.fir@101283.4]
  assign _T_951 = _T_949 & _T_947; // @[Monitor.scala 682:54:freechips.rocketchip.system.DefaultRV32Config.fir@101285.4]
  assign _T_953 = |inflight; // @[Monitor.scala 687:26:freechips.rocketchip.system.DefaultRV32Config.fir@101290.4]
  assign _T_954 = ~_T_953; // @[Monitor.scala 687:16:freechips.rocketchip.system.DefaultRV32Config.fir@101291.4]
  assign _T_955 = plusarg_reader_out == 32'h0; // @[Monitor.scala 687:39:freechips.rocketchip.system.DefaultRV32Config.fir@101292.4]
  assign _T_956 = _T_954 | _T_955; // @[Monitor.scala 687:30:freechips.rocketchip.system.DefaultRV32Config.fir@101293.4]
  assign _T_957 = _T_952 < plusarg_reader_out; // @[Monitor.scala 687:59:freechips.rocketchip.system.DefaultRV32Config.fir@101294.4]
  assign _T_958 = _T_956 | _T_957; // @[Monitor.scala 687:47:freechips.rocketchip.system.DefaultRV32Config.fir@101295.4]
  assign _T_960 = _T_958 | reset; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@101297.4]
  assign _T_961 = ~_T_960; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@101298.4]
  assign _T_963 = _T_952 + 32'h1; // @[Monitor.scala 689:26:freechips.rocketchip.system.DefaultRV32Config.fir@101304.4]
  assign _T_966 = _T_702 | _T_751; // @[Monitor.scala 690:27:freechips.rocketchip.system.DefaultRV32Config.fir@101308.4]
  assign _GEN_67 = io_in_a_valid & _T_56; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@99906.10]
  assign _GEN_75 = io_in_a_valid & _T_124; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@100008.10]
  assign _GEN_85 = io_in_a_valid & _T_196; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@100121.10]
  assign _GEN_91 = io_in_a_valid & _T_259; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@100210.10]
  assign _GEN_97 = io_in_a_valid & _T_318; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@100291.10]
  assign _GEN_101 = io_in_a_valid & _T_379; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@100371.10]
  assign _GEN_107 = io_in_a_valid & _T_435; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@100449.10]
  assign _GEN_113 = io_in_a_valid & _T_491; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@100527.10]
  assign _GEN_119 = io_in_d_valid & _T_558; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@100590.10]
  assign _GEN_129 = io_in_d_valid & _T_578; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@100632.10]
  assign _GEN_141 = io_in_d_valid & _T_606; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@100690.10]
  assign _GEN_153 = io_in_d_valid & _T_635; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@100749.10]
  assign _GEN_159 = io_in_d_valid & _T_652; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@100784.10]
  assign _GEN_165 = io_in_d_valid & _T_670; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@100820.10]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_711 = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  _T_722 = _RAND_1[2:0];
  _RAND_2 = {1{`RANDOM}};
  _T_726 = _RAND_2[8:0];
  _RAND_3 = {1{`RANDOM}};
  _T_759 = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  _T_770 = _RAND_4[2:0];
  _RAND_5 = {1{`RANDOM}};
  _T_771 = _RAND_5[1:0];
  _RAND_6 = {1{`RANDOM}};
  _T_772 = _RAND_6[1:0];
  _RAND_7 = {1{`RANDOM}};
  _T_773 = _RAND_7[0:0];
  _RAND_8 = {1{`RANDOM}};
  _T_774 = _RAND_8[0:0];
  _RAND_9 = {1{`RANDOM}};
  _T_775 = _RAND_9[0:0];
  _RAND_10 = {1{`RANDOM}};
  inflight = _RAND_10[0:0];
  _RAND_11 = {1{`RANDOM}};
  inflight_opcodes = _RAND_11[3:0];
  _RAND_12 = {1{`RANDOM}};
  inflight_sizes = _RAND_12[3:0];
  _RAND_13 = {1{`RANDOM}};
  _T_813 = _RAND_13[0:0];
  _RAND_14 = {1{`RANDOM}};
  _T_831 = _RAND_14[0:0];
  _RAND_15 = {1{`RANDOM}};
  _T_952 = _RAND_15[31:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      _T_711 <= 1'h0;
    end else if (_T_702) begin
      if (_T_714) begin
        _T_711 <= 1'h0;
      end else begin
        _T_711 <= _T_713;
      end
    end
    if (_T_750) begin
      _T_722 <= io_in_a_bits_opcode;
    end
    if (_T_750) begin
      _T_726 <= io_in_a_bits_address;
    end
    if (reset) begin
      _T_759 <= 1'h0;
    end else if (_T_751) begin
      if (_T_762) begin
        _T_759 <= 1'h0;
      end else begin
        _T_759 <= _T_761;
      end
    end
    if (_T_803) begin
      _T_770 <= io_in_d_bits_opcode;
    end
    if (_T_803) begin
      _T_771 <= io_in_d_bits_param;
    end
    if (_T_803) begin
      _T_772 <= io_in_d_bits_size;
    end
    if (_T_803) begin
      _T_773 <= io_in_d_bits_source;
    end
    if (_T_803) begin
      _T_774 <= io_in_d_bits_sink;
    end
    if (_T_803) begin
      _T_775 <= io_in_d_bits_denied;
    end
    if (reset) begin
      inflight <= 1'h0;
    end else begin
      inflight <= _T_945;
    end
    if (reset) begin
      inflight_opcodes <= 4'h0;
    end else begin
      inflight_opcodes <= _T_948;
    end
    if (reset) begin
      inflight_sizes <= 4'h0;
    end else begin
      inflight_sizes <= _T_951;
    end
    if (reset) begin
      _T_813 <= 1'h0;
    end else if (_T_702) begin
      if (a_first) begin
        _T_813 <= 1'h0;
      end else begin
        _T_813 <= _T_815;
      end
    end
    if (reset) begin
      _T_831 <= 1'h0;
    end else if (_T_751) begin
      if (d_first) begin
        _T_831 <= 1'h0;
      end else begin
        _T_831 <= _T_833;
      end
    end
    if (reset) begin
      _T_952 <= 32'h0;
    end else if (_T_966) begin
      _T_952 <= 32'h0;
    end else begin
      _T_952 <= _T_963;
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_67 & _T_97) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel carries AcquireBlock type unsupported by manager (connected at BusBypass.scala:35:12)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@99906.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_67 & _T_97) begin
          $fatal; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@99907.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_67 & _T_97) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel carries AcquireBlock from a client which does not support Probe (connected at BusBypass.scala:35:12)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@99913.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_67 & _T_97) begin
          $fatal; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@99914.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_67 & _T_110) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel AcquireBlock address not aligned to size (connected at BusBypass.scala:35:12)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@99935.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_67 & _T_110) begin
          $fatal; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@99936.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_67 & _T_119) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel AcquireBlock contains invalid mask (connected at BusBypass.scala:35:12)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@99952.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_67 & _T_119) begin
          $fatal; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@99953.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_75 & _T_97) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel carries AcquirePerm type unsupported by manager (connected at BusBypass.scala:35:12)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@100008.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_75 & _T_97) begin
          $fatal; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@100009.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_75 & _T_97) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel carries AcquirePerm from a client which does not support Probe (connected at BusBypass.scala:35:12)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@100015.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_75 & _T_97) begin
          $fatal; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@100016.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_75 & _T_110) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel AcquirePerm address not aligned to size (connected at BusBypass.scala:35:12)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@100037.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_75 & _T_110) begin
          $fatal; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@100038.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_75 & _T_97) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel AcquirePerm requests NtoB (connected at BusBypass.scala:35:12)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@100053.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_75 & _T_97) begin
          $fatal; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@100054.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_75 & _T_119) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel AcquirePerm contains invalid mask (connected at BusBypass.scala:35:12)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@100062.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_75 & _T_119) begin
          $fatal; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@100063.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_85 & _T_240) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel carries Get type unsupported by manager (connected at BusBypass.scala:35:12)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@100121.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_85 & _T_240) begin
          $fatal; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@100122.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_85 & _T_110) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel Get address not aligned to size (connected at BusBypass.scala:35:12)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@100135.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_85 & _T_110) begin
          $fatal; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@100136.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_85 & _T_254) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel Get contains invalid mask (connected at BusBypass.scala:35:12)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@100151.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_85 & _T_254) begin
          $fatal; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@100152.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_91 & _T_240) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel carries PutFull type unsupported by manager (connected at BusBypass.scala:35:12)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@100210.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_91 & _T_240) begin
          $fatal; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@100211.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_91 & _T_110) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel PutFull address not aligned to size (connected at BusBypass.scala:35:12)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@100224.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_91 & _T_110) begin
          $fatal; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@100225.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_91 & _T_254) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel PutFull contains invalid mask (connected at BusBypass.scala:35:12)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@100240.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_91 & _T_254) begin
          $fatal; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@100241.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_97 & _T_240) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel carries PutPartial type unsupported by manager (connected at BusBypass.scala:35:12)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@100291.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_97 & _T_240) begin
          $fatal; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@100292.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_97 & _T_110) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel PutPartial address not aligned to size (connected at BusBypass.scala:35:12)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@100305.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_97 & _T_110) begin
          $fatal; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@100306.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_101 & _T_97) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel carries Arithmetic type unsupported by manager (connected at BusBypass.scala:35:12)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@100371.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_101 & _T_97) begin
          $fatal; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@100372.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_101 & _T_110) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel Arithmetic address not aligned to size (connected at BusBypass.scala:35:12)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@100385.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_101 & _T_110) begin
          $fatal; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@100386.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_101 & _T_254) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel Arithmetic contains invalid mask (connected at BusBypass.scala:35:12)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@100401.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_101 & _T_254) begin
          $fatal; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@100402.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_107 & _T_97) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel carries Logical type unsupported by manager (connected at BusBypass.scala:35:12)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@100449.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_107 & _T_97) begin
          $fatal; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@100450.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_107 & _T_110) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel Logical address not aligned to size (connected at BusBypass.scala:35:12)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@100463.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_107 & _T_110) begin
          $fatal; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@100464.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_107 & _T_254) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel Logical contains invalid mask (connected at BusBypass.scala:35:12)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@100479.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_107 & _T_254) begin
          $fatal; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@100480.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_113 & _T_97) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel carries Hint type unsupported by manager (connected at BusBypass.scala:35:12)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@100527.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_113 & _T_97) begin
          $fatal; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@100528.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_113 & _T_110) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel Hint address not aligned to size (connected at BusBypass.scala:35:12)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@100541.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_113 & _T_110) begin
          $fatal; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@100542.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_113 & _T_254) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel Hint contains invalid mask (connected at BusBypass.scala:35:12)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@100557.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_113 & _T_254) begin
          $fatal; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@100558.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_d_valid & _T_554) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel has invalid opcode (connected at BusBypass.scala:35:12)\n    at Monitor.scala:51 assert(cond, message)\n"); // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@100576.8]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_d_valid & _T_554) begin
          $fatal; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@100577.8]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_119 & _T_561) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel ReleaseAck carries invalid source ID (connected at BusBypass.scala:35:12)\n    at Monitor.scala:51 assert(cond, message)\n"); // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@100590.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_119 & _T_561) begin
          $fatal; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@100591.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_119 & _T_565) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel ReleaseAck smaller than a beat (connected at BusBypass.scala:35:12)\n    at Monitor.scala:51 assert(cond, message)\n"); // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@100598.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_119 & _T_565) begin
          $fatal; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@100599.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_119 & _T_569) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel ReleaseeAck carries invalid param (connected at BusBypass.scala:35:12)\n    at Monitor.scala:51 assert(cond, message)\n"); // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@100606.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_119 & _T_569) begin
          $fatal; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@100607.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_119 & _T_573) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel ReleaseAck is corrupt (connected at BusBypass.scala:35:12)\n    at Monitor.scala:51 assert(cond, message)\n"); // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@100614.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_119 & _T_573) begin
          $fatal; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@100615.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_119 & _T_577) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel ReleaseAck is denied (connected at BusBypass.scala:35:12)\n    at Monitor.scala:51 assert(cond, message)\n"); // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@100622.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_119 & _T_577) begin
          $fatal; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@100623.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_129 & _T_561) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel Grant carries invalid source ID (connected at BusBypass.scala:35:12)\n    at Monitor.scala:51 assert(cond, message)\n"); // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@100632.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_129 & _T_561) begin
          $fatal; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@100633.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_129 & _T_97) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel Grant carries invalid sink ID (connected at BusBypass.scala:35:12)\n    at Monitor.scala:51 assert(cond, message)\n"); // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@100639.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_129 & _T_97) begin
          $fatal; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@100640.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_129 & _T_565) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel Grant smaller than a beat (connected at BusBypass.scala:35:12)\n    at Monitor.scala:51 assert(cond, message)\n"); // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@100647.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_129 & _T_565) begin
          $fatal; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@100648.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_129 & _T_592) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel Grant carries invalid cap param (connected at BusBypass.scala:35:12)\n    at Monitor.scala:51 assert(cond, message)\n"); // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@100655.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_129 & _T_592) begin
          $fatal; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@100656.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_129 & _T_596) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel Grant carries toN param (connected at BusBypass.scala:35:12)\n    at Monitor.scala:51 assert(cond, message)\n"); // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@100663.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_129 & _T_596) begin
          $fatal; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@100664.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_129 & _T_573) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel Grant is corrupt (connected at BusBypass.scala:35:12)\n    at Monitor.scala:51 assert(cond, message)\n"); // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@100671.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_129 & _T_573) begin
          $fatal; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@100672.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_141 & _T_561) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel GrantData carries invalid source ID (connected at BusBypass.scala:35:12)\n    at Monitor.scala:51 assert(cond, message)\n"); // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@100690.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_141 & _T_561) begin
          $fatal; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@100691.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_141 & _T_97) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel GrantData carries invalid sink ID (connected at BusBypass.scala:35:12)\n    at Monitor.scala:51 assert(cond, message)\n"); // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@100697.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_141 & _T_97) begin
          $fatal; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@100698.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_141 & _T_565) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel GrantData smaller than a beat (connected at BusBypass.scala:35:12)\n    at Monitor.scala:51 assert(cond, message)\n"); // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@100705.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_141 & _T_565) begin
          $fatal; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@100706.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_141 & _T_592) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel GrantData carries invalid cap param (connected at BusBypass.scala:35:12)\n    at Monitor.scala:51 assert(cond, message)\n"); // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@100713.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_141 & _T_592) begin
          $fatal; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@100714.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_141 & _T_596) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel GrantData carries toN param (connected at BusBypass.scala:35:12)\n    at Monitor.scala:51 assert(cond, message)\n"); // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@100721.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_141 & _T_596) begin
          $fatal; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@100722.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_141 & _T_629) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel GrantData is denied but not corrupt (connected at BusBypass.scala:35:12)\n    at Monitor.scala:51 assert(cond, message)\n"); // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@100730.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_141 & _T_629) begin
          $fatal; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@100731.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_153 & _T_561) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel AccessAck carries invalid source ID (connected at BusBypass.scala:35:12)\n    at Monitor.scala:51 assert(cond, message)\n"); // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@100749.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_153 & _T_561) begin
          $fatal; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@100750.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_153 & _T_569) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel AccessAck carries invalid param (connected at BusBypass.scala:35:12)\n    at Monitor.scala:51 assert(cond, message)\n"); // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@100757.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_153 & _T_569) begin
          $fatal; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@100758.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_153 & _T_573) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel AccessAck is corrupt (connected at BusBypass.scala:35:12)\n    at Monitor.scala:51 assert(cond, message)\n"); // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@100765.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_153 & _T_573) begin
          $fatal; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@100766.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_159 & _T_561) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel AccessAckData carries invalid source ID (connected at BusBypass.scala:35:12)\n    at Monitor.scala:51 assert(cond, message)\n"); // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@100784.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_159 & _T_561) begin
          $fatal; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@100785.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_159 & _T_569) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel AccessAckData carries invalid param (connected at BusBypass.scala:35:12)\n    at Monitor.scala:51 assert(cond, message)\n"); // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@100792.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_159 & _T_569) begin
          $fatal; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@100793.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_159 & _T_629) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel AccessAckData is denied but not corrupt (connected at BusBypass.scala:35:12)\n    at Monitor.scala:51 assert(cond, message)\n"); // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@100801.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_159 & _T_629) begin
          $fatal; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@100802.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_165 & _T_561) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel HintAck carries invalid source ID (connected at BusBypass.scala:35:12)\n    at Monitor.scala:51 assert(cond, message)\n"); // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@100820.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_165 & _T_561) begin
          $fatal; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@100821.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_165 & _T_569) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel HintAck carries invalid param (connected at BusBypass.scala:35:12)\n    at Monitor.scala:51 assert(cond, message)\n"); // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@100828.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_165 & _T_569) begin
          $fatal; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@100829.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_165 & _T_573) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel HintAck is corrupt (connected at BusBypass.scala:35:12)\n    at Monitor.scala:51 assert(cond, message)\n"); // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@100836.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_165 & _T_573) begin
          $fatal; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@100837.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_728 & _T_732) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel opcode changed within multibeat operation (connected at BusBypass.scala:35:12)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@100916.8]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_728 & _T_732) begin
          $fatal; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@100917.8]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_728 & _T_748) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel address changed with multibeat operation (connected at BusBypass.scala:35:12)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@100948.8]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_728 & _T_748) begin
          $fatal; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@100949.8]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_777 & _T_781) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel opcode changed within multibeat operation (connected at BusBypass.scala:35:12)\n    at Monitor.scala:51 assert(cond, message)\n"); // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@100997.8]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_777 & _T_781) begin
          $fatal; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@100998.8]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_777 & _T_785) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel param changed within multibeat operation (connected at BusBypass.scala:35:12)\n    at Monitor.scala:51 assert(cond, message)\n"); // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@101005.8]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_777 & _T_785) begin
          $fatal; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@101006.8]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_777 & _T_789) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel size changed within multibeat operation (connected at BusBypass.scala:35:12)\n    at Monitor.scala:51 assert(cond, message)\n"); // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@101013.8]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_777 & _T_789) begin
          $fatal; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@101014.8]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_777 & _T_793) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel source changed within multibeat operation (connected at BusBypass.scala:35:12)\n    at Monitor.scala:51 assert(cond, message)\n"); // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@101021.8]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_777 & _T_793) begin
          $fatal; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@101022.8]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_777 & _T_797) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel sink changed with multibeat operation (connected at BusBypass.scala:35:12)\n    at Monitor.scala:51 assert(cond, message)\n"); // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@101029.8]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_777 & _T_797) begin
          $fatal; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@101030.8]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_777 & _T_801) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel denied changed with multibeat operation (connected at BusBypass.scala:35:12)\n    at Monitor.scala:51 assert(cond, message)\n"); // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@101037.8]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_777 & _T_801) begin
          $fatal; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@101038.8]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_860 & _T_876) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel re-used a source ID (connected at BusBypass.scala:35:12)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@101174.8]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_860 & _T_876) begin
          $fatal; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@101175.8]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_899 & _T_910) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel acknowledged for nothing inflight (connected at BusBypass.scala:35:12)\n    at Monitor.scala:51 assert(cond, message)\n"); // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@101225.8]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_899 & _T_910) begin
          $fatal; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@101226.8]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_899 & _T_923) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel contains improper opcode response (connected at BusBypass.scala:35:12)\n    at Monitor.scala:51 assert(cond, message)\n"); // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@101242.8]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_899 & _T_923) begin
          $fatal; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@101243.8]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_899 & _T_930) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel contains improper response size (connected at BusBypass.scala:35:12)\n    at Monitor.scala:51 assert(cond, message)\n"); // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@101253.8]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_899 & _T_930) begin
          $fatal; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@101254.8]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_937 & _T_942) begin
          $fwrite(32'h80000002,"Assertion failed: ready check\n    at Monitor.scala:51 assert(cond, message)\n"); // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@101271.8]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_937 & _T_942) begin
          $fatal; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@101272.8]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_961) begin
          $fwrite(32'h80000002,"Assertion failed: TileLink timeout expired (connected at BusBypass.scala:35:12)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@101300.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_961) begin
          $fatal; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@101301.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
  end
endmodule
