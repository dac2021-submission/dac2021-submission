module ClockGroupAggregator_1( // @[:freechips.rocketchip.system.DefaultRV32Config.fir@29037.2]
  input   auto_in_member_0_clock, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@29038.4]
  input   auto_in_member_0_reset, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@29038.4]
  output  auto_out_member_0_clock, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@29038.4]
  output  auto_out_member_0_reset // @[:freechips.rocketchip.system.DefaultRV32Config.fir@29038.4]
);
  assign auto_out_member_0_clock = auto_in_member_0_clock; // @[LazyModule.scala 305:12:freechips.rocketchip.system.DefaultRV32Config.fir@29052.4]
  assign auto_out_member_0_reset = auto_in_member_0_reset; // @[LazyModule.scala 305:12:freechips.rocketchip.system.DefaultRV32Config.fir@29052.4]
endmodule
