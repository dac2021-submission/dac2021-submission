module TLMonitor_48( // @[:freechips.rocketchip.system.DefaultRV32Config.fir@207093.2]
  input         clock, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@207094.4]
  input         reset, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@207095.4]
  input         io_in_a_ready, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@207096.4]
  input         io_in_a_valid, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@207096.4]
  input  [2:0]  io_in_a_bits_opcode, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@207096.4]
  input  [2:0]  io_in_a_bits_param, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@207096.4]
  input  [3:0]  io_in_a_bits_size, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@207096.4]
  input  [1:0]  io_in_a_bits_source, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@207096.4]
  input  [31:0] io_in_a_bits_address, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@207096.4]
  input  [3:0]  io_in_a_bits_mask, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@207096.4]
  input         io_in_a_bits_corrupt, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@207096.4]
  input         io_in_b_ready, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@207096.4]
  input         io_in_b_valid, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@207096.4]
  input  [2:0]  io_in_b_bits_opcode, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@207096.4]
  input  [1:0]  io_in_b_bits_param, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@207096.4]
  input  [3:0]  io_in_b_bits_size, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@207096.4]
  input  [1:0]  io_in_b_bits_source, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@207096.4]
  input  [31:0] io_in_b_bits_address, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@207096.4]
  input  [3:0]  io_in_b_bits_mask, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@207096.4]
  input         io_in_b_bits_corrupt, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@207096.4]
  input         io_in_c_ready, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@207096.4]
  input         io_in_c_valid, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@207096.4]
  input  [2:0]  io_in_c_bits_opcode, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@207096.4]
  input  [2:0]  io_in_c_bits_param, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@207096.4]
  input  [3:0]  io_in_c_bits_size, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@207096.4]
  input  [1:0]  io_in_c_bits_source, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@207096.4]
  input  [31:0] io_in_c_bits_address, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@207096.4]
  input         io_in_d_ready, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@207096.4]
  input         io_in_d_valid, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@207096.4]
  input  [2:0]  io_in_d_bits_opcode, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@207096.4]
  input  [1:0]  io_in_d_bits_param, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@207096.4]
  input  [3:0]  io_in_d_bits_size, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@207096.4]
  input  [1:0]  io_in_d_bits_source, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@207096.4]
  input  [1:0]  io_in_d_bits_sink, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@207096.4]
  input         io_in_d_bits_denied, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@207096.4]
  input         io_in_d_bits_corrupt, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@207096.4]
  input         io_in_e_ready, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@207096.4]
  input         io_in_e_valid, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@207096.4]
  input  [1:0]  io_in_e_bits_sink // @[:freechips.rocketchip.system.DefaultRV32Config.fir@207096.4]
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
`endif // RANDOMIZE_REG_INIT
  wire [31:0] plusarg_reader_out; // @[PlusArg.scala 80:11:freechips.rocketchip.system.DefaultRV32Config.fir@209959.4]
  wire  _T_4; // @[Parameters.scala 47:9:freechips.rocketchip.system.DefaultRV32Config.fir@207107.6]
  wire  _T_5; // @[Parameters.scala 47:9:freechips.rocketchip.system.DefaultRV32Config.fir@207108.6]
  wire  _T_6; // @[Parameters.scala 47:9:freechips.rocketchip.system.DefaultRV32Config.fir@207109.6]
  wire  _T_8; // @[Parameters.scala 924:46:freechips.rocketchip.system.DefaultRV32Config.fir@207115.6]
  wire  _T_9; // @[Parameters.scala 924:46:freechips.rocketchip.system.DefaultRV32Config.fir@207116.6]
  wire [26:0] _T_11; // @[package.scala 207:77:freechips.rocketchip.system.DefaultRV32Config.fir@207118.6]
  wire [11:0] _T_13; // @[package.scala 207:46:freechips.rocketchip.system.DefaultRV32Config.fir@207120.6]
  wire [31:0] _GEN_71; // @[Edges.scala 22:16:freechips.rocketchip.system.DefaultRV32Config.fir@207121.6]
  wire [31:0] _T_14; // @[Edges.scala 22:16:freechips.rocketchip.system.DefaultRV32Config.fir@207121.6]
  wire  _T_15; // @[Edges.scala 22:24:freechips.rocketchip.system.DefaultRV32Config.fir@207122.6]
  wire [1:0] _T_18; // @[OneHot.scala 65:12:freechips.rocketchip.system.DefaultRV32Config.fir@207125.6]
  wire [1:0] _T_20; // @[Misc.scala 201:81:freechips.rocketchip.system.DefaultRV32Config.fir@207127.6]
  wire  _T_21; // @[Misc.scala 205:21:freechips.rocketchip.system.DefaultRV32Config.fir@207128.6]
  wire  _T_24; // @[Misc.scala 210:20:freechips.rocketchip.system.DefaultRV32Config.fir@207131.6]
  wire  _T_26; // @[Misc.scala 214:38:freechips.rocketchip.system.DefaultRV32Config.fir@207133.6]
  wire  _T_27; // @[Misc.scala 214:29:freechips.rocketchip.system.DefaultRV32Config.fir@207134.6]
  wire  _T_29; // @[Misc.scala 214:38:freechips.rocketchip.system.DefaultRV32Config.fir@207136.6]
  wire  _T_30; // @[Misc.scala 214:29:freechips.rocketchip.system.DefaultRV32Config.fir@207137.6]
  wire  _T_33; // @[Misc.scala 210:20:freechips.rocketchip.system.DefaultRV32Config.fir@207140.6]
  wire  _T_34; // @[Misc.scala 213:27:freechips.rocketchip.system.DefaultRV32Config.fir@207141.6]
  wire  _T_35; // @[Misc.scala 214:38:freechips.rocketchip.system.DefaultRV32Config.fir@207142.6]
  wire  _T_36; // @[Misc.scala 214:29:freechips.rocketchip.system.DefaultRV32Config.fir@207143.6]
  wire  _T_37; // @[Misc.scala 213:27:freechips.rocketchip.system.DefaultRV32Config.fir@207144.6]
  wire  _T_38; // @[Misc.scala 214:38:freechips.rocketchip.system.DefaultRV32Config.fir@207145.6]
  wire  _T_39; // @[Misc.scala 214:29:freechips.rocketchip.system.DefaultRV32Config.fir@207146.6]
  wire  _T_40; // @[Misc.scala 213:27:freechips.rocketchip.system.DefaultRV32Config.fir@207147.6]
  wire  _T_41; // @[Misc.scala 214:38:freechips.rocketchip.system.DefaultRV32Config.fir@207148.6]
  wire  _T_42; // @[Misc.scala 214:29:freechips.rocketchip.system.DefaultRV32Config.fir@207149.6]
  wire  _T_43; // @[Misc.scala 213:27:freechips.rocketchip.system.DefaultRV32Config.fir@207150.6]
  wire  _T_44; // @[Misc.scala 214:38:freechips.rocketchip.system.DefaultRV32Config.fir@207151.6]
  wire  _T_45; // @[Misc.scala 214:29:freechips.rocketchip.system.DefaultRV32Config.fir@207152.6]
  wire [3:0] _T_48; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@207155.6]
  wire [32:0] _T_52; // @[Parameters.scala 137:49:freechips.rocketchip.system.DefaultRV32Config.fir@207159.6]
  wire  _T_78; // @[Monitor.scala 79:25:freechips.rocketchip.system.DefaultRV32Config.fir@207189.6]
  wire [32:0] _T_83; // @[Parameters.scala 137:52:freechips.rocketchip.system.DefaultRV32Config.fir@207195.8]
  wire  _T_84; // @[Parameters.scala 137:67:freechips.rocketchip.system.DefaultRV32Config.fir@207196.8]
  wire [31:0] _T_85; // @[Parameters.scala 137:31:freechips.rocketchip.system.DefaultRV32Config.fir@207197.8]
  wire [32:0] _T_86; // @[Parameters.scala 137:49:freechips.rocketchip.system.DefaultRV32Config.fir@207198.8]
  wire [32:0] _T_88; // @[Parameters.scala 137:52:freechips.rocketchip.system.DefaultRV32Config.fir@207200.8]
  wire  _T_89; // @[Parameters.scala 137:67:freechips.rocketchip.system.DefaultRV32Config.fir@207201.8]
  wire [31:0] _T_90; // @[Parameters.scala 137:31:freechips.rocketchip.system.DefaultRV32Config.fir@207202.8]
  wire [32:0] _T_91; // @[Parameters.scala 137:49:freechips.rocketchip.system.DefaultRV32Config.fir@207203.8]
  wire [32:0] _T_93; // @[Parameters.scala 137:52:freechips.rocketchip.system.DefaultRV32Config.fir@207205.8]
  wire  _T_94; // @[Parameters.scala 137:67:freechips.rocketchip.system.DefaultRV32Config.fir@207206.8]
  wire [31:0] _T_95; // @[Parameters.scala 137:31:freechips.rocketchip.system.DefaultRV32Config.fir@207207.8]
  wire [32:0] _T_96; // @[Parameters.scala 137:49:freechips.rocketchip.system.DefaultRV32Config.fir@207208.8]
  wire [32:0] _T_98; // @[Parameters.scala 137:52:freechips.rocketchip.system.DefaultRV32Config.fir@207210.8]
  wire  _T_99; // @[Parameters.scala 137:67:freechips.rocketchip.system.DefaultRV32Config.fir@207211.8]
  wire [31:0] _T_100; // @[Parameters.scala 137:31:freechips.rocketchip.system.DefaultRV32Config.fir@207212.8]
  wire [32:0] _T_101; // @[Parameters.scala 137:49:freechips.rocketchip.system.DefaultRV32Config.fir@207213.8]
  wire [32:0] _T_103; // @[Parameters.scala 137:52:freechips.rocketchip.system.DefaultRV32Config.fir@207215.8]
  wire  _T_104; // @[Parameters.scala 137:67:freechips.rocketchip.system.DefaultRV32Config.fir@207216.8]
  wire [31:0] _T_105; // @[Parameters.scala 137:31:freechips.rocketchip.system.DefaultRV32Config.fir@207217.8]
  wire [32:0] _T_106; // @[Parameters.scala 137:49:freechips.rocketchip.system.DefaultRV32Config.fir@207218.8]
  wire [32:0] _T_108; // @[Parameters.scala 137:52:freechips.rocketchip.system.DefaultRV32Config.fir@207220.8]
  wire  _T_109; // @[Parameters.scala 137:67:freechips.rocketchip.system.DefaultRV32Config.fir@207221.8]
  wire  _T_110; // @[Parameters.scala 552:42:freechips.rocketchip.system.DefaultRV32Config.fir@207222.8]
  wire  _T_117; // @[Parameters.scala 93:42:freechips.rocketchip.system.DefaultRV32Config.fir@207229.8]
  wire [31:0] _T_120; // @[Parameters.scala 137:31:freechips.rocketchip.system.DefaultRV32Config.fir@207232.8]
  wire [32:0] _T_121; // @[Parameters.scala 137:49:freechips.rocketchip.system.DefaultRV32Config.fir@207233.8]
  wire [32:0] _T_123; // @[Parameters.scala 137:52:freechips.rocketchip.system.DefaultRV32Config.fir@207235.8]
  wire  _T_124; // @[Parameters.scala 137:67:freechips.rocketchip.system.DefaultRV32Config.fir@207236.8]
  wire  _T_125; // @[Parameters.scala 551:56:freechips.rocketchip.system.DefaultRV32Config.fir@207237.8]
  wire  _T_129; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@207241.8]
  wire  _T_130; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@207242.8]
  wire  _T_135; // @[Parameters.scala 92:48:freechips.rocketchip.system.DefaultRV32Config.fir@207255.8]
  wire  _T_136; // @[Mux.scala 27:72:freechips.rocketchip.system.DefaultRV32Config.fir@207256.8]
  wire  _T_143; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@207264.8]
  wire  _T_144; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@207265.8]
  wire  _T_146; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@207271.8]
  wire  _T_147; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@207272.8]
  wire  _T_150; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@207279.8]
  wire  _T_151; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@207280.8]
  wire  _T_153; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@207286.8]
  wire  _T_154; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@207287.8]
  wire  _T_155; // @[Bundles.scala 110:27:freechips.rocketchip.system.DefaultRV32Config.fir@207292.8]
  wire  _T_157; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@207294.8]
  wire  _T_158; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@207295.8]
  wire [3:0] _T_159; // @[Monitor.scala 86:18:freechips.rocketchip.system.DefaultRV32Config.fir@207300.8]
  wire  _T_160; // @[Monitor.scala 86:31:freechips.rocketchip.system.DefaultRV32Config.fir@207301.8]
  wire  _T_162; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@207303.8]
  wire  _T_163; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@207304.8]
  wire  _T_164; // @[Monitor.scala 87:18:freechips.rocketchip.system.DefaultRV32Config.fir@207309.8]
  wire  _T_166; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@207311.8]
  wire  _T_167; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@207312.8]
  wire  _T_168; // @[Monitor.scala 90:25:freechips.rocketchip.system.DefaultRV32Config.fir@207318.6]
  wire  _T_249; // @[Monitor.scala 97:31:freechips.rocketchip.system.DefaultRV32Config.fir@207429.8]
  wire  _T_251; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@207431.8]
  wire  _T_252; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@207432.8]
  wire  _T_262; // @[Monitor.scala 102:25:freechips.rocketchip.system.DefaultRV32Config.fir@207455.6]
  wire  _T_264; // @[Parameters.scala 93:42:freechips.rocketchip.system.DefaultRV32Config.fir@207458.8]
  wire  _T_272; // @[Parameters.scala 551:56:freechips.rocketchip.system.DefaultRV32Config.fir@207466.8]
  wire  _T_307; // @[Parameters.scala 552:42:freechips.rocketchip.system.DefaultRV32Config.fir@207501.8]
  wire  _T_308; // @[Parameters.scala 552:42:freechips.rocketchip.system.DefaultRV32Config.fir@207502.8]
  wire  _T_309; // @[Parameters.scala 552:42:freechips.rocketchip.system.DefaultRV32Config.fir@207503.8]
  wire  _T_310; // @[Parameters.scala 552:42:freechips.rocketchip.system.DefaultRV32Config.fir@207504.8]
  wire  _T_311; // @[Parameters.scala 552:42:freechips.rocketchip.system.DefaultRV32Config.fir@207505.8]
  wire  _T_312; // @[Parameters.scala 551:56:freechips.rocketchip.system.DefaultRV32Config.fir@207506.8]
  wire  _T_314; // @[Parameters.scala 553:30:freechips.rocketchip.system.DefaultRV32Config.fir@207508.8]
  wire  _T_316; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@207510.8]
  wire  _T_317; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@207511.8]
  wire  _T_324; // @[Monitor.scala 106:31:freechips.rocketchip.system.DefaultRV32Config.fir@207530.8]
  wire  _T_326; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@207532.8]
  wire  _T_327; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@207533.8]
  wire  _T_328; // @[Monitor.scala 107:30:freechips.rocketchip.system.DefaultRV32Config.fir@207538.8]
  wire  _T_330; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@207540.8]
  wire  _T_331; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@207541.8]
  wire  _T_336; // @[Monitor.scala 111:25:freechips.rocketchip.system.DefaultRV32Config.fir@207555.6]
  wire  _T_371; // @[Parameters.scala 552:42:freechips.rocketchip.system.DefaultRV32Config.fir@207591.8]
  wire  _T_372; // @[Parameters.scala 552:42:freechips.rocketchip.system.DefaultRV32Config.fir@207592.8]
  wire  _T_373; // @[Parameters.scala 552:42:freechips.rocketchip.system.DefaultRV32Config.fir@207593.8]
  wire  _T_374; // @[Parameters.scala 551:56:freechips.rocketchip.system.DefaultRV32Config.fir@207594.8]
  wire  _T_383; // @[Parameters.scala 93:42:freechips.rocketchip.system.DefaultRV32Config.fir@207603.8]
  wire  _T_391; // @[Parameters.scala 551:56:freechips.rocketchip.system.DefaultRV32Config.fir@207611.8]
  wire  _T_393; // @[Parameters.scala 553:30:freechips.rocketchip.system.DefaultRV32Config.fir@207613.8]
  wire  _T_395; // @[Parameters.scala 553:30:freechips.rocketchip.system.DefaultRV32Config.fir@207615.8]
  wire  _T_397; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@207617.8]
  wire  _T_398; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@207618.8]
  wire  _T_413; // @[Monitor.scala 119:25:freechips.rocketchip.system.DefaultRV32Config.fir@207654.6]
  wire [3:0] _T_486; // @[Monitor.scala 124:33:freechips.rocketchip.system.DefaultRV32Config.fir@207744.8]
  wire [3:0] _T_487; // @[Monitor.scala 124:31:freechips.rocketchip.system.DefaultRV32Config.fir@207745.8]
  wire  _T_488; // @[Monitor.scala 124:40:freechips.rocketchip.system.DefaultRV32Config.fir@207746.8]
  wire  _T_490; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@207748.8]
  wire  _T_491; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@207749.8]
  wire  _T_492; // @[Monitor.scala 127:25:freechips.rocketchip.system.DefaultRV32Config.fir@207755.6]
  wire  _T_494; // @[Parameters.scala 93:42:freechips.rocketchip.system.DefaultRV32Config.fir@207758.8]
  wire  _T_518; // @[Parameters.scala 552:42:freechips.rocketchip.system.DefaultRV32Config.fir@207782.8]
  wire  _T_519; // @[Parameters.scala 552:42:freechips.rocketchip.system.DefaultRV32Config.fir@207783.8]
  wire  _T_520; // @[Parameters.scala 551:56:freechips.rocketchip.system.DefaultRV32Config.fir@207784.8]
  wire  _T_543; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@207807.8]
  wire  _T_544; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@207808.8]
  wire  _T_551; // @[Bundles.scala 140:33:freechips.rocketchip.system.DefaultRV32Config.fir@207827.8]
  wire  _T_553; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@207829.8]
  wire  _T_554; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@207830.8]
  wire  _T_559; // @[Monitor.scala 135:25:freechips.rocketchip.system.DefaultRV32Config.fir@207844.6]
  wire  _T_618; // @[Bundles.scala 147:30:freechips.rocketchip.system.DefaultRV32Config.fir@207916.8]
  wire  _T_620; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@207918.8]
  wire  _T_621; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@207919.8]
  wire  _T_626; // @[Monitor.scala 143:25:freechips.rocketchip.system.DefaultRV32Config.fir@207933.6]
  wire  _T_677; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@207985.8]
  wire  _T_678; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@207986.8]
  wire  _T_685; // @[Bundles.scala 160:28:freechips.rocketchip.system.DefaultRV32Config.fir@208005.8]
  wire  _T_687; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@208007.8]
  wire  _T_688; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@208008.8]
  wire  _T_697; // @[Bundles.scala 44:24:freechips.rocketchip.system.DefaultRV32Config.fir@208032.6]
  wire  _T_699; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@208034.6]
  wire  _T_700; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@208035.6]
  wire  _T_701; // @[Parameters.scala 47:9:freechips.rocketchip.system.DefaultRV32Config.fir@208040.6]
  wire  _T_702; // @[Parameters.scala 47:9:freechips.rocketchip.system.DefaultRV32Config.fir@208041.6]
  wire  _T_703; // @[Parameters.scala 47:9:freechips.rocketchip.system.DefaultRV32Config.fir@208042.6]
  wire  _T_705; // @[Parameters.scala 924:46:freechips.rocketchip.system.DefaultRV32Config.fir@208048.6]
  wire  _T_706; // @[Parameters.scala 924:46:freechips.rocketchip.system.DefaultRV32Config.fir@208049.6]
  wire  _T_708; // @[Monitor.scala 307:25:freechips.rocketchip.system.DefaultRV32Config.fir@208051.6]
  wire  _T_710; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@208054.8]
  wire  _T_711; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@208055.8]
  wire  _T_712; // @[Monitor.scala 309:27:freechips.rocketchip.system.DefaultRV32Config.fir@208060.8]
  wire  _T_714; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@208062.8]
  wire  _T_715; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@208063.8]
  wire  _T_716; // @[Monitor.scala 310:28:freechips.rocketchip.system.DefaultRV32Config.fir@208068.8]
  wire  _T_718; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@208070.8]
  wire  _T_719; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@208071.8]
  wire  _T_720; // @[Monitor.scala 311:15:freechips.rocketchip.system.DefaultRV32Config.fir@208076.8]
  wire  _T_722; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@208078.8]
  wire  _T_723; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@208079.8]
  wire  _T_724; // @[Monitor.scala 312:15:freechips.rocketchip.system.DefaultRV32Config.fir@208084.8]
  wire  _T_726; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@208086.8]
  wire  _T_727; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@208087.8]
  wire  _T_728; // @[Monitor.scala 315:25:freechips.rocketchip.system.DefaultRV32Config.fir@208093.6]
  wire  _T_739; // @[Bundles.scala 104:26:freechips.rocketchip.system.DefaultRV32Config.fir@208117.8]
  wire  _T_741; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@208119.8]
  wire  _T_742; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@208120.8]
  wire  _T_743; // @[Monitor.scala 320:28:freechips.rocketchip.system.DefaultRV32Config.fir@208125.8]
  wire  _T_745; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@208127.8]
  wire  _T_746; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@208128.8]
  wire  _T_756; // @[Monitor.scala 325:25:freechips.rocketchip.system.DefaultRV32Config.fir@208151.6]
  wire  _T_776; // @[Monitor.scala 331:30:freechips.rocketchip.system.DefaultRV32Config.fir@208192.8]
  wire  _T_778; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@208194.8]
  wire  _T_779; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@208195.8]
  wire  _T_785; // @[Monitor.scala 335:25:freechips.rocketchip.system.DefaultRV32Config.fir@208210.6]
  wire  _T_802; // @[Monitor.scala 343:25:freechips.rocketchip.system.DefaultRV32Config.fir@208245.6]
  wire  _T_820; // @[Monitor.scala 351:25:freechips.rocketchip.system.DefaultRV32Config.fir@208281.6]
  wire  _T_837; // @[Bundles.scala 42:24:freechips.rocketchip.system.DefaultRV32Config.fir@208318.6]
  wire  _T_839; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@208320.6]
  wire  _T_840; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@208321.6]
  wire  _T_841; // @[Parameters.scala 47:9:freechips.rocketchip.system.DefaultRV32Config.fir@208326.6]
  wire [32:0] _T_844; // @[Parameters.scala 137:49:freechips.rocketchip.system.DefaultRV32Config.fir@208329.6]
  wire  _T_849; // @[Parameters.scala 47:9:freechips.rocketchip.system.DefaultRV32Config.fir@208334.6]
  wire  _T_857; // @[Parameters.scala 47:9:freechips.rocketchip.system.DefaultRV32Config.fir@208342.6]
  wire [31:0] _T_870; // @[Parameters.scala 137:31:freechips.rocketchip.system.DefaultRV32Config.fir@208359.6]
  wire [32:0] _T_871; // @[Parameters.scala 137:49:freechips.rocketchip.system.DefaultRV32Config.fir@208360.6]
  wire [32:0] _T_873; // @[Parameters.scala 137:52:freechips.rocketchip.system.DefaultRV32Config.fir@208362.6]
  wire  _T_874; // @[Parameters.scala 137:67:freechips.rocketchip.system.DefaultRV32Config.fir@208363.6]
  wire [31:0] _T_875; // @[Parameters.scala 137:31:freechips.rocketchip.system.DefaultRV32Config.fir@208364.6]
  wire [32:0] _T_876; // @[Parameters.scala 137:49:freechips.rocketchip.system.DefaultRV32Config.fir@208365.6]
  wire [32:0] _T_878; // @[Parameters.scala 137:52:freechips.rocketchip.system.DefaultRV32Config.fir@208367.6]
  wire  _T_879; // @[Parameters.scala 137:67:freechips.rocketchip.system.DefaultRV32Config.fir@208368.6]
  wire [31:0] _T_880; // @[Parameters.scala 137:31:freechips.rocketchip.system.DefaultRV32Config.fir@208369.6]
  wire [32:0] _T_881; // @[Parameters.scala 137:49:freechips.rocketchip.system.DefaultRV32Config.fir@208370.6]
  wire [32:0] _T_883; // @[Parameters.scala 137:52:freechips.rocketchip.system.DefaultRV32Config.fir@208372.6]
  wire  _T_884; // @[Parameters.scala 137:67:freechips.rocketchip.system.DefaultRV32Config.fir@208373.6]
  wire [32:0] _T_888; // @[Parameters.scala 137:52:freechips.rocketchip.system.DefaultRV32Config.fir@208377.6]
  wire  _T_889; // @[Parameters.scala 137:67:freechips.rocketchip.system.DefaultRV32Config.fir@208378.6]
  wire [31:0] _T_890; // @[Parameters.scala 137:31:freechips.rocketchip.system.DefaultRV32Config.fir@208379.6]
  wire [32:0] _T_891; // @[Parameters.scala 137:49:freechips.rocketchip.system.DefaultRV32Config.fir@208380.6]
  wire [32:0] _T_893; // @[Parameters.scala 137:52:freechips.rocketchip.system.DefaultRV32Config.fir@208382.6]
  wire  _T_894; // @[Parameters.scala 137:67:freechips.rocketchip.system.DefaultRV32Config.fir@208383.6]
  wire [31:0] _T_895; // @[Parameters.scala 137:31:freechips.rocketchip.system.DefaultRV32Config.fir@208384.6]
  wire [32:0] _T_896; // @[Parameters.scala 137:49:freechips.rocketchip.system.DefaultRV32Config.fir@208385.6]
  wire [32:0] _T_898; // @[Parameters.scala 137:52:freechips.rocketchip.system.DefaultRV32Config.fir@208387.6]
  wire  _T_899; // @[Parameters.scala 137:67:freechips.rocketchip.system.DefaultRV32Config.fir@208388.6]
  wire [31:0] _T_900; // @[Parameters.scala 137:31:freechips.rocketchip.system.DefaultRV32Config.fir@208389.6]
  wire [32:0] _T_901; // @[Parameters.scala 137:49:freechips.rocketchip.system.DefaultRV32Config.fir@208390.6]
  wire [32:0] _T_903; // @[Parameters.scala 137:52:freechips.rocketchip.system.DefaultRV32Config.fir@208392.6]
  wire  _T_904; // @[Parameters.scala 137:67:freechips.rocketchip.system.DefaultRV32Config.fir@208393.6]
  wire  _T_906; // @[Parameters.scala 535:64:freechips.rocketchip.system.DefaultRV32Config.fir@208403.6]
  wire  _T_907; // @[Parameters.scala 535:64:freechips.rocketchip.system.DefaultRV32Config.fir@208404.6]
  wire  _T_908; // @[Parameters.scala 535:64:freechips.rocketchip.system.DefaultRV32Config.fir@208405.6]
  wire  _T_909; // @[Parameters.scala 535:64:freechips.rocketchip.system.DefaultRV32Config.fir@208406.6]
  wire  _T_910; // @[Parameters.scala 535:64:freechips.rocketchip.system.DefaultRV32Config.fir@208407.6]
  wire  _T_911; // @[Parameters.scala 535:64:freechips.rocketchip.system.DefaultRV32Config.fir@208408.6]
  wire [26:0] _T_913; // @[package.scala 207:77:freechips.rocketchip.system.DefaultRV32Config.fir@208410.6]
  wire [11:0] _T_915; // @[package.scala 207:46:freechips.rocketchip.system.DefaultRV32Config.fir@208412.6]
  wire [31:0] _GEN_72; // @[Edges.scala 22:16:freechips.rocketchip.system.DefaultRV32Config.fir@208413.6]
  wire [31:0] _T_916; // @[Edges.scala 22:16:freechips.rocketchip.system.DefaultRV32Config.fir@208413.6]
  wire  _T_917; // @[Edges.scala 22:24:freechips.rocketchip.system.DefaultRV32Config.fir@208414.6]
  wire [1:0] _T_920; // @[OneHot.scala 65:12:freechips.rocketchip.system.DefaultRV32Config.fir@208417.6]
  wire [1:0] _T_922; // @[Misc.scala 201:81:freechips.rocketchip.system.DefaultRV32Config.fir@208419.6]
  wire  _T_923; // @[Misc.scala 205:21:freechips.rocketchip.system.DefaultRV32Config.fir@208420.6]
  wire  _T_926; // @[Misc.scala 210:20:freechips.rocketchip.system.DefaultRV32Config.fir@208423.6]
  wire  _T_928; // @[Misc.scala 214:38:freechips.rocketchip.system.DefaultRV32Config.fir@208425.6]
  wire  _T_929; // @[Misc.scala 214:29:freechips.rocketchip.system.DefaultRV32Config.fir@208426.6]
  wire  _T_931; // @[Misc.scala 214:38:freechips.rocketchip.system.DefaultRV32Config.fir@208428.6]
  wire  _T_932; // @[Misc.scala 214:29:freechips.rocketchip.system.DefaultRV32Config.fir@208429.6]
  wire  _T_935; // @[Misc.scala 210:20:freechips.rocketchip.system.DefaultRV32Config.fir@208432.6]
  wire  _T_936; // @[Misc.scala 213:27:freechips.rocketchip.system.DefaultRV32Config.fir@208433.6]
  wire  _T_937; // @[Misc.scala 214:38:freechips.rocketchip.system.DefaultRV32Config.fir@208434.6]
  wire  _T_938; // @[Misc.scala 214:29:freechips.rocketchip.system.DefaultRV32Config.fir@208435.6]
  wire  _T_939; // @[Misc.scala 213:27:freechips.rocketchip.system.DefaultRV32Config.fir@208436.6]
  wire  _T_940; // @[Misc.scala 214:38:freechips.rocketchip.system.DefaultRV32Config.fir@208437.6]
  wire  _T_941; // @[Misc.scala 214:29:freechips.rocketchip.system.DefaultRV32Config.fir@208438.6]
  wire  _T_942; // @[Misc.scala 213:27:freechips.rocketchip.system.DefaultRV32Config.fir@208439.6]
  wire  _T_943; // @[Misc.scala 214:38:freechips.rocketchip.system.DefaultRV32Config.fir@208440.6]
  wire  _T_944; // @[Misc.scala 214:29:freechips.rocketchip.system.DefaultRV32Config.fir@208441.6]
  wire  _T_945; // @[Misc.scala 213:27:freechips.rocketchip.system.DefaultRV32Config.fir@208442.6]
  wire  _T_946; // @[Misc.scala 214:38:freechips.rocketchip.system.DefaultRV32Config.fir@208443.6]
  wire  _T_947; // @[Misc.scala 214:29:freechips.rocketchip.system.DefaultRV32Config.fir@208444.6]
  wire [3:0] _T_950; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@208447.6]
  wire [1:0] _T_957; // @[Mux.scala 27:72:freechips.rocketchip.system.DefaultRV32Config.fir@208458.6]
  wire [1:0] _GEN_73; // @[Mux.scala 27:72:freechips.rocketchip.system.DefaultRV32Config.fir@208460.6]
  wire [1:0] _T_959; // @[Mux.scala 27:72:freechips.rocketchip.system.DefaultRV32Config.fir@208460.6]
  wire  _T_961; // @[Monitor.scala 162:113:freechips.rocketchip.system.DefaultRV32Config.fir@208463.6]
  wire  _T_962; // @[Monitor.scala 164:25:freechips.rocketchip.system.DefaultRV32Config.fir@208464.6]
  wire  _T_967; // @[Parameters.scala 92:48:freechips.rocketchip.system.DefaultRV32Config.fir@208474.8]
  wire  _T_968; // @[Mux.scala 27:72:freechips.rocketchip.system.DefaultRV32Config.fir@208475.8]
  wire  _T_975; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@208483.8]
  wire  _T_976; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@208484.8]
  wire  _T_978; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@208490.8]
  wire  _T_979; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@208491.8]
  wire  _T_981; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@208497.8]
  wire  _T_982; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@208498.8]
  wire  _T_984; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@208504.8]
  wire  _T_985; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@208505.8]
  wire  _T_986; // @[Bundles.scala 104:26:freechips.rocketchip.system.DefaultRV32Config.fir@208510.8]
  wire  _T_988; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@208512.8]
  wire  _T_989; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@208513.8]
  wire  _T_990; // @[Monitor.scala 170:30:freechips.rocketchip.system.DefaultRV32Config.fir@208518.8]
  wire  _T_992; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@208520.8]
  wire  _T_993; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@208521.8]
  wire  _T_994; // @[Monitor.scala 171:18:freechips.rocketchip.system.DefaultRV32Config.fir@208526.8]
  wire  _T_996; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@208528.8]
  wire  _T_997; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@208529.8]
  wire  _T_998; // @[Monitor.scala 174:25:freechips.rocketchip.system.DefaultRV32Config.fir@208535.6]
  wire  _T_1001; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@208539.8]
  wire  _T_1011; // @[Monitor.scala 179:31:freechips.rocketchip.system.DefaultRV32Config.fir@208565.8]
  wire  _T_1013; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@208567.8]
  wire  _T_1014; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@208568.8]
  wire  _T_1023; // @[Monitor.scala 184:25:freechips.rocketchip.system.DefaultRV32Config.fir@208590.6]
  wire  _T_1044; // @[Monitor.scala 193:25:freechips.rocketchip.system.DefaultRV32Config.fir@208637.6]
  wire [3:0] _T_1061; // @[Monitor.scala 199:33:freechips.rocketchip.system.DefaultRV32Config.fir@208675.8]
  wire [3:0] _T_1062; // @[Monitor.scala 199:31:freechips.rocketchip.system.DefaultRV32Config.fir@208676.8]
  wire  _T_1063; // @[Monitor.scala 199:40:freechips.rocketchip.system.DefaultRV32Config.fir@208677.8]
  wire  _T_1065; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@208679.8]
  wire  _T_1066; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@208680.8]
  wire  _T_1067; // @[Monitor.scala 202:25:freechips.rocketchip.system.DefaultRV32Config.fir@208686.6]
  wire  _T_1088; // @[Monitor.scala 211:25:freechips.rocketchip.system.DefaultRV32Config.fir@208733.6]
  wire  _T_1109; // @[Monitor.scala 220:25:freechips.rocketchip.system.DefaultRV32Config.fir@208780.6]
  wire  _T_1134; // @[Parameters.scala 47:9:freechips.rocketchip.system.DefaultRV32Config.fir@208837.6]
  wire  _T_1135; // @[Parameters.scala 47:9:freechips.rocketchip.system.DefaultRV32Config.fir@208838.6]
  wire  _T_1136; // @[Parameters.scala 47:9:freechips.rocketchip.system.DefaultRV32Config.fir@208839.6]
  wire  _T_1138; // @[Parameters.scala 924:46:freechips.rocketchip.system.DefaultRV32Config.fir@208845.6]
  wire  _T_1139; // @[Parameters.scala 924:46:freechips.rocketchip.system.DefaultRV32Config.fir@208846.6]
  wire [26:0] _T_1141; // @[package.scala 207:77:freechips.rocketchip.system.DefaultRV32Config.fir@208848.6]
  wire [11:0] _T_1143; // @[package.scala 207:46:freechips.rocketchip.system.DefaultRV32Config.fir@208850.6]
  wire [31:0] _GEN_74; // @[Edges.scala 22:16:freechips.rocketchip.system.DefaultRV32Config.fir@208851.6]
  wire [31:0] _T_1144; // @[Edges.scala 22:16:freechips.rocketchip.system.DefaultRV32Config.fir@208851.6]
  wire  _T_1145; // @[Edges.scala 22:24:freechips.rocketchip.system.DefaultRV32Config.fir@208852.6]
  wire [31:0] _T_1146; // @[Parameters.scala 137:31:freechips.rocketchip.system.DefaultRV32Config.fir@208853.6]
  wire [32:0] _T_1147; // @[Parameters.scala 137:49:freechips.rocketchip.system.DefaultRV32Config.fir@208854.6]
  wire [32:0] _T_1149; // @[Parameters.scala 137:52:freechips.rocketchip.system.DefaultRV32Config.fir@208856.6]
  wire  _T_1150; // @[Parameters.scala 137:67:freechips.rocketchip.system.DefaultRV32Config.fir@208857.6]
  wire [31:0] _T_1151; // @[Parameters.scala 137:31:freechips.rocketchip.system.DefaultRV32Config.fir@208858.6]
  wire [32:0] _T_1152; // @[Parameters.scala 137:49:freechips.rocketchip.system.DefaultRV32Config.fir@208859.6]
  wire [32:0] _T_1154; // @[Parameters.scala 137:52:freechips.rocketchip.system.DefaultRV32Config.fir@208861.6]
  wire  _T_1155; // @[Parameters.scala 137:67:freechips.rocketchip.system.DefaultRV32Config.fir@208862.6]
  wire [31:0] _T_1156; // @[Parameters.scala 137:31:freechips.rocketchip.system.DefaultRV32Config.fir@208863.6]
  wire [32:0] _T_1157; // @[Parameters.scala 137:49:freechips.rocketchip.system.DefaultRV32Config.fir@208864.6]
  wire [32:0] _T_1159; // @[Parameters.scala 137:52:freechips.rocketchip.system.DefaultRV32Config.fir@208866.6]
  wire  _T_1160; // @[Parameters.scala 137:67:freechips.rocketchip.system.DefaultRV32Config.fir@208867.6]
  wire [32:0] _T_1162; // @[Parameters.scala 137:49:freechips.rocketchip.system.DefaultRV32Config.fir@208869.6]
  wire [32:0] _T_1164; // @[Parameters.scala 137:52:freechips.rocketchip.system.DefaultRV32Config.fir@208871.6]
  wire  _T_1165; // @[Parameters.scala 137:67:freechips.rocketchip.system.DefaultRV32Config.fir@208872.6]
  wire [31:0] _T_1166; // @[Parameters.scala 137:31:freechips.rocketchip.system.DefaultRV32Config.fir@208873.6]
  wire [32:0] _T_1167; // @[Parameters.scala 137:49:freechips.rocketchip.system.DefaultRV32Config.fir@208874.6]
  wire [32:0] _T_1169; // @[Parameters.scala 137:52:freechips.rocketchip.system.DefaultRV32Config.fir@208876.6]
  wire  _T_1170; // @[Parameters.scala 137:67:freechips.rocketchip.system.DefaultRV32Config.fir@208877.6]
  wire [31:0] _T_1171; // @[Parameters.scala 137:31:freechips.rocketchip.system.DefaultRV32Config.fir@208878.6]
  wire [32:0] _T_1172; // @[Parameters.scala 137:49:freechips.rocketchip.system.DefaultRV32Config.fir@208879.6]
  wire [32:0] _T_1174; // @[Parameters.scala 137:52:freechips.rocketchip.system.DefaultRV32Config.fir@208881.6]
  wire  _T_1175; // @[Parameters.scala 137:67:freechips.rocketchip.system.DefaultRV32Config.fir@208882.6]
  wire [31:0] _T_1176; // @[Parameters.scala 137:31:freechips.rocketchip.system.DefaultRV32Config.fir@208883.6]
  wire [32:0] _T_1177; // @[Parameters.scala 137:49:freechips.rocketchip.system.DefaultRV32Config.fir@208884.6]
  wire [32:0] _T_1179; // @[Parameters.scala 137:52:freechips.rocketchip.system.DefaultRV32Config.fir@208886.6]
  wire  _T_1180; // @[Parameters.scala 137:67:freechips.rocketchip.system.DefaultRV32Config.fir@208887.6]
  wire  _T_1182; // @[Parameters.scala 535:64:freechips.rocketchip.system.DefaultRV32Config.fir@208897.6]
  wire  _T_1183; // @[Parameters.scala 535:64:freechips.rocketchip.system.DefaultRV32Config.fir@208898.6]
  wire  _T_1184; // @[Parameters.scala 535:64:freechips.rocketchip.system.DefaultRV32Config.fir@208899.6]
  wire  _T_1185; // @[Parameters.scala 535:64:freechips.rocketchip.system.DefaultRV32Config.fir@208900.6]
  wire  _T_1186; // @[Parameters.scala 535:64:freechips.rocketchip.system.DefaultRV32Config.fir@208901.6]
  wire  _T_1187; // @[Parameters.scala 535:64:freechips.rocketchip.system.DefaultRV32Config.fir@208902.6]
  wire  _T_1217; // @[Monitor.scala 239:25:freechips.rocketchip.system.DefaultRV32Config.fir@208936.6]
  wire  _T_1219; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@208939.8]
  wire  _T_1220; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@208940.8]
  wire  _T_1222; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@208946.8]
  wire  _T_1223; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@208947.8]
  wire  _T_1224; // @[Monitor.scala 242:30:freechips.rocketchip.system.DefaultRV32Config.fir@208952.8]
  wire  _T_1226; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@208954.8]
  wire  _T_1227; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@208955.8]
  wire  _T_1229; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@208961.8]
  wire  _T_1230; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@208962.8]
  wire  _T_1231; // @[Bundles.scala 122:29:freechips.rocketchip.system.DefaultRV32Config.fir@208967.8]
  wire  _T_1233; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@208969.8]
  wire  _T_1234; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@208970.8]
  wire  _T_1239; // @[Monitor.scala 248:25:freechips.rocketchip.system.DefaultRV32Config.fir@208984.6]
  wire  _T_1257; // @[Monitor.scala 256:25:freechips.rocketchip.system.DefaultRV32Config.fir@209024.6]
  wire  _T_1296; // @[Parameters.scala 93:42:freechips.rocketchip.system.DefaultRV32Config.fir@209064.8]
  wire  _T_1304; // @[Parameters.scala 551:56:freechips.rocketchip.system.DefaultRV32Config.fir@209072.8]
  wire  _T_1308; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@209076.8]
  wire  _T_1309; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@209077.8]
  wire  _T_1314; // @[Parameters.scala 92:48:freechips.rocketchip.system.DefaultRV32Config.fir@209090.8]
  wire  _T_1315; // @[Mux.scala 27:72:freechips.rocketchip.system.DefaultRV32Config.fir@209091.8]
  wire  _T_1322; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@209099.8]
  wire  _T_1323; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@209100.8]
  wire  _T_1334; // @[Bundles.scala 116:29:freechips.rocketchip.system.DefaultRV32Config.fir@209127.8]
  wire  _T_1336; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@209129.8]
  wire  _T_1337; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@209130.8]
  wire  _T_1342; // @[Monitor.scala 266:25:freechips.rocketchip.system.DefaultRV32Config.fir@209144.6]
  wire  _T_1423; // @[Monitor.scala 275:25:freechips.rocketchip.system.DefaultRV32Config.fir@209256.6]
  wire  _T_1433; // @[Monitor.scala 279:31:freechips.rocketchip.system.DefaultRV32Config.fir@209279.8]
  wire  _T_1435; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@209281.8]
  wire  _T_1436; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@209282.8]
  wire  _T_1441; // @[Monitor.scala 283:25:freechips.rocketchip.system.DefaultRV32Config.fir@209296.6]
  wire  _T_1455; // @[Monitor.scala 290:25:freechips.rocketchip.system.DefaultRV32Config.fir@209328.6]
  wire  _T_1477; // @[Decoupled.scala 40:37:freechips.rocketchip.system.DefaultRV32Config.fir@209379.4]
  wire  _T_1484; // @[Edges.scala 93:28:freechips.rocketchip.system.DefaultRV32Config.fir@209386.4]
  reg [9:0] _T_1486; // @[Edges.scala 230:27:freechips.rocketchip.system.DefaultRV32Config.fir@209388.4]
  wire [9:0] _T_1488; // @[Edges.scala 231:28:freechips.rocketchip.system.DefaultRV32Config.fir@209390.4]
  wire  _T_1489; // @[Edges.scala 232:25:freechips.rocketchip.system.DefaultRV32Config.fir@209391.4]
  reg [2:0] _T_1497; // @[Monitor.scala 381:22:freechips.rocketchip.system.DefaultRV32Config.fir@209402.4]
  reg [2:0] _T_1498; // @[Monitor.scala 382:22:freechips.rocketchip.system.DefaultRV32Config.fir@209403.4]
  reg [3:0] _T_1499; // @[Monitor.scala 383:22:freechips.rocketchip.system.DefaultRV32Config.fir@209404.4]
  reg [1:0] _T_1500; // @[Monitor.scala 384:22:freechips.rocketchip.system.DefaultRV32Config.fir@209405.4]
  reg [31:0] _T_1501; // @[Monitor.scala 385:22:freechips.rocketchip.system.DefaultRV32Config.fir@209406.4]
  wire  _T_1502; // @[Monitor.scala 386:22:freechips.rocketchip.system.DefaultRV32Config.fir@209407.4]
  wire  _T_1503; // @[Monitor.scala 386:19:freechips.rocketchip.system.DefaultRV32Config.fir@209408.4]
  wire  _T_1504; // @[Monitor.scala 387:32:freechips.rocketchip.system.DefaultRV32Config.fir@209410.6]
  wire  _T_1506; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@209412.6]
  wire  _T_1507; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@209413.6]
  wire  _T_1508; // @[Monitor.scala 388:32:freechips.rocketchip.system.DefaultRV32Config.fir@209418.6]
  wire  _T_1510; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@209420.6]
  wire  _T_1511; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@209421.6]
  wire  _T_1512; // @[Monitor.scala 389:32:freechips.rocketchip.system.DefaultRV32Config.fir@209426.6]
  wire  _T_1514; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@209428.6]
  wire  _T_1515; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@209429.6]
  wire  _T_1516; // @[Monitor.scala 390:32:freechips.rocketchip.system.DefaultRV32Config.fir@209434.6]
  wire  _T_1518; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@209436.6]
  wire  _T_1519; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@209437.6]
  wire  _T_1520; // @[Monitor.scala 391:32:freechips.rocketchip.system.DefaultRV32Config.fir@209442.6]
  wire  _T_1522; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@209444.6]
  wire  _T_1523; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@209445.6]
  wire  _T_1525; // @[Monitor.scala 393:20:freechips.rocketchip.system.DefaultRV32Config.fir@209452.4]
  wire  _T_1526; // @[Decoupled.scala 40:37:freechips.rocketchip.system.DefaultRV32Config.fir@209460.4]
  wire [26:0] _T_1528; // @[package.scala 207:77:freechips.rocketchip.system.DefaultRV32Config.fir@209462.4]
  wire [11:0] _T_1530; // @[package.scala 207:46:freechips.rocketchip.system.DefaultRV32Config.fir@209464.4]
  reg [9:0] _T_1534; // @[Edges.scala 230:27:freechips.rocketchip.system.DefaultRV32Config.fir@209468.4]
  wire [9:0] _T_1536; // @[Edges.scala 231:28:freechips.rocketchip.system.DefaultRV32Config.fir@209470.4]
  wire  _T_1537; // @[Edges.scala 232:25:freechips.rocketchip.system.DefaultRV32Config.fir@209471.4]
  reg [2:0] _T_1545; // @[Monitor.scala 532:22:freechips.rocketchip.system.DefaultRV32Config.fir@209482.4]
  reg [1:0] _T_1546; // @[Monitor.scala 533:22:freechips.rocketchip.system.DefaultRV32Config.fir@209483.4]
  reg [3:0] _T_1547; // @[Monitor.scala 534:22:freechips.rocketchip.system.DefaultRV32Config.fir@209484.4]
  reg [1:0] _T_1548; // @[Monitor.scala 535:22:freechips.rocketchip.system.DefaultRV32Config.fir@209485.4]
  reg [1:0] _T_1549; // @[Monitor.scala 536:22:freechips.rocketchip.system.DefaultRV32Config.fir@209486.4]
  reg  _T_1550; // @[Monitor.scala 537:22:freechips.rocketchip.system.DefaultRV32Config.fir@209487.4]
  wire  _T_1551; // @[Monitor.scala 538:22:freechips.rocketchip.system.DefaultRV32Config.fir@209488.4]
  wire  _T_1552; // @[Monitor.scala 538:19:freechips.rocketchip.system.DefaultRV32Config.fir@209489.4]
  wire  _T_1553; // @[Monitor.scala 539:29:freechips.rocketchip.system.DefaultRV32Config.fir@209491.6]
  wire  _T_1555; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@209493.6]
  wire  _T_1556; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@209494.6]
  wire  _T_1557; // @[Monitor.scala 540:29:freechips.rocketchip.system.DefaultRV32Config.fir@209499.6]
  wire  _T_1559; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@209501.6]
  wire  _T_1560; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@209502.6]
  wire  _T_1561; // @[Monitor.scala 541:29:freechips.rocketchip.system.DefaultRV32Config.fir@209507.6]
  wire  _T_1563; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@209509.6]
  wire  _T_1564; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@209510.6]
  wire  _T_1565; // @[Monitor.scala 542:29:freechips.rocketchip.system.DefaultRV32Config.fir@209515.6]
  wire  _T_1567; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@209517.6]
  wire  _T_1568; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@209518.6]
  wire  _T_1569; // @[Monitor.scala 543:29:freechips.rocketchip.system.DefaultRV32Config.fir@209523.6]
  wire  _T_1571; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@209525.6]
  wire  _T_1572; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@209526.6]
  wire  _T_1573; // @[Monitor.scala 544:29:freechips.rocketchip.system.DefaultRV32Config.fir@209531.6]
  wire  _T_1575; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@209533.6]
  wire  _T_1576; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@209534.6]
  wire  _T_1578; // @[Monitor.scala 546:20:freechips.rocketchip.system.DefaultRV32Config.fir@209541.4]
  wire  _T_1579; // @[Decoupled.scala 40:37:freechips.rocketchip.system.DefaultRV32Config.fir@209550.4]
  reg [9:0] _T_1588; // @[Edges.scala 230:27:freechips.rocketchip.system.DefaultRV32Config.fir@209559.4]
  wire [9:0] _T_1590; // @[Edges.scala 231:28:freechips.rocketchip.system.DefaultRV32Config.fir@209561.4]
  wire  _T_1591; // @[Edges.scala 232:25:freechips.rocketchip.system.DefaultRV32Config.fir@209562.4]
  reg [2:0] _T_1599; // @[Monitor.scala 404:22:freechips.rocketchip.system.DefaultRV32Config.fir@209573.4]
  reg [1:0] _T_1600; // @[Monitor.scala 405:22:freechips.rocketchip.system.DefaultRV32Config.fir@209574.4]
  reg [3:0] _T_1601; // @[Monitor.scala 406:22:freechips.rocketchip.system.DefaultRV32Config.fir@209575.4]
  reg [1:0] _T_1602; // @[Monitor.scala 407:22:freechips.rocketchip.system.DefaultRV32Config.fir@209576.4]
  reg [31:0] _T_1603; // @[Monitor.scala 408:22:freechips.rocketchip.system.DefaultRV32Config.fir@209577.4]
  wire  _T_1604; // @[Monitor.scala 409:22:freechips.rocketchip.system.DefaultRV32Config.fir@209578.4]
  wire  _T_1605; // @[Monitor.scala 409:19:freechips.rocketchip.system.DefaultRV32Config.fir@209579.4]
  wire  _T_1606; // @[Monitor.scala 410:32:freechips.rocketchip.system.DefaultRV32Config.fir@209581.6]
  wire  _T_1608; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@209583.6]
  wire  _T_1609; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@209584.6]
  wire  _T_1610; // @[Monitor.scala 411:32:freechips.rocketchip.system.DefaultRV32Config.fir@209589.6]
  wire  _T_1612; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@209591.6]
  wire  _T_1613; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@209592.6]
  wire  _T_1614; // @[Monitor.scala 412:32:freechips.rocketchip.system.DefaultRV32Config.fir@209597.6]
  wire  _T_1616; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@209599.6]
  wire  _T_1617; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@209600.6]
  wire  _T_1618; // @[Monitor.scala 413:32:freechips.rocketchip.system.DefaultRV32Config.fir@209605.6]
  wire  _T_1620; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@209607.6]
  wire  _T_1621; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@209608.6]
  wire  _T_1622; // @[Monitor.scala 414:32:freechips.rocketchip.system.DefaultRV32Config.fir@209613.6]
  wire  _T_1624; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@209615.6]
  wire  _T_1625; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@209616.6]
  wire  _T_1627; // @[Monitor.scala 416:20:freechips.rocketchip.system.DefaultRV32Config.fir@209623.4]
  wire  _T_1628; // @[Decoupled.scala 40:37:freechips.rocketchip.system.DefaultRV32Config.fir@209631.4]
  reg [9:0] _T_1636; // @[Edges.scala 230:27:freechips.rocketchip.system.DefaultRV32Config.fir@209639.4]
  wire [9:0] _T_1638; // @[Edges.scala 231:28:freechips.rocketchip.system.DefaultRV32Config.fir@209641.4]
  wire  _T_1639; // @[Edges.scala 232:25:freechips.rocketchip.system.DefaultRV32Config.fir@209642.4]
  reg [2:0] _T_1647; // @[Monitor.scala 509:22:freechips.rocketchip.system.DefaultRV32Config.fir@209653.4]
  reg [2:0] _T_1648; // @[Monitor.scala 510:22:freechips.rocketchip.system.DefaultRV32Config.fir@209654.4]
  reg [3:0] _T_1649; // @[Monitor.scala 511:22:freechips.rocketchip.system.DefaultRV32Config.fir@209655.4]
  reg [1:0] _T_1650; // @[Monitor.scala 512:22:freechips.rocketchip.system.DefaultRV32Config.fir@209656.4]
  reg [31:0] _T_1651; // @[Monitor.scala 513:22:freechips.rocketchip.system.DefaultRV32Config.fir@209657.4]
  wire  _T_1652; // @[Monitor.scala 514:22:freechips.rocketchip.system.DefaultRV32Config.fir@209658.4]
  wire  _T_1653; // @[Monitor.scala 514:19:freechips.rocketchip.system.DefaultRV32Config.fir@209659.4]
  wire  _T_1654; // @[Monitor.scala 515:32:freechips.rocketchip.system.DefaultRV32Config.fir@209661.6]
  wire  _T_1656; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@209663.6]
  wire  _T_1657; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@209664.6]
  wire  _T_1658; // @[Monitor.scala 516:32:freechips.rocketchip.system.DefaultRV32Config.fir@209669.6]
  wire  _T_1660; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@209671.6]
  wire  _T_1661; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@209672.6]
  wire  _T_1662; // @[Monitor.scala 517:32:freechips.rocketchip.system.DefaultRV32Config.fir@209677.6]
  wire  _T_1664; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@209679.6]
  wire  _T_1665; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@209680.6]
  wire  _T_1666; // @[Monitor.scala 518:32:freechips.rocketchip.system.DefaultRV32Config.fir@209685.6]
  wire  _T_1668; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@209687.6]
  wire  _T_1669; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@209688.6]
  wire  _T_1670; // @[Monitor.scala 519:32:freechips.rocketchip.system.DefaultRV32Config.fir@209693.6]
  wire  _T_1672; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@209695.6]
  wire  _T_1673; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@209696.6]
  wire  _T_1675; // @[Monitor.scala 521:20:freechips.rocketchip.system.DefaultRV32Config.fir@209703.4]
  reg [2:0] inflight; // @[Monitor.scala 608:27:freechips.rocketchip.system.DefaultRV32Config.fir@209711.4]
  reg [11:0] inflight_opcodes; // @[Monitor.scala 610:35:freechips.rocketchip.system.DefaultRV32Config.fir@209712.4]
  reg [23:0] inflight_sizes; // @[Monitor.scala 612:33:freechips.rocketchip.system.DefaultRV32Config.fir@209713.4]
  reg [9:0] _T_1685; // @[Edges.scala 230:27:freechips.rocketchip.system.DefaultRV32Config.fir@209723.4]
  wire [9:0] _T_1687; // @[Edges.scala 231:28:freechips.rocketchip.system.DefaultRV32Config.fir@209725.4]
  wire  a_first; // @[Edges.scala 232:25:freechips.rocketchip.system.DefaultRV32Config.fir@209726.4]
  reg [9:0] _T_1703; // @[Edges.scala 230:27:freechips.rocketchip.system.DefaultRV32Config.fir@209745.4]
  wire [9:0] _T_1705; // @[Edges.scala 231:28:freechips.rocketchip.system.DefaultRV32Config.fir@209747.4]
  wire  d_first; // @[Edges.scala 232:25:freechips.rocketchip.system.DefaultRV32Config.fir@209748.4]
  wire [3:0] _GEN_75; // @[Monitor.scala 629:69:freechips.rocketchip.system.DefaultRV32Config.fir@209767.4]
  wire [4:0] _T_1713; // @[Monitor.scala 629:69:freechips.rocketchip.system.DefaultRV32Config.fir@209767.4]
  wire [11:0] _T_1714; // @[Monitor.scala 629:44:freechips.rocketchip.system.DefaultRV32Config.fir@209768.4]
  wire [15:0] _T_1718; // @[Monitor.scala 606:57:freechips.rocketchip.system.DefaultRV32Config.fir@209772.4]
  wire [15:0] _GEN_76; // @[Monitor.scala 629:97:freechips.rocketchip.system.DefaultRV32Config.fir@209773.4]
  wire [15:0] _T_1719; // @[Monitor.scala 629:97:freechips.rocketchip.system.DefaultRV32Config.fir@209773.4]
  wire [15:0] _T_1720; // @[Monitor.scala 629:152:freechips.rocketchip.system.DefaultRV32Config.fir@209774.4]
  wire [4:0] _T_1721; // @[Monitor.scala 633:65:freechips.rocketchip.system.DefaultRV32Config.fir@209778.4]
  wire [23:0] _T_1722; // @[Monitor.scala 633:40:freechips.rocketchip.system.DefaultRV32Config.fir@209779.4]
  wire [15:0] _T_1726; // @[Monitor.scala 606:57:freechips.rocketchip.system.DefaultRV32Config.fir@209783.4]
  wire [23:0] _GEN_78; // @[Monitor.scala 633:91:freechips.rocketchip.system.DefaultRV32Config.fir@209784.4]
  wire [23:0] _T_1727; // @[Monitor.scala 633:91:freechips.rocketchip.system.DefaultRV32Config.fir@209784.4]
  wire [23:0] _T_1728; // @[Monitor.scala 633:144:freechips.rocketchip.system.DefaultRV32Config.fir@209785.4]
  wire  _T_1732; // @[Monitor.scala 643:27:freechips.rocketchip.system.DefaultRV32Config.fir@209810.4]
  wire [3:0] _T_1734; // @[OneHot.scala 58:35:freechips.rocketchip.system.DefaultRV32Config.fir@209813.6]
  wire [3:0] _T_1735; // @[Monitor.scala 645:53:freechips.rocketchip.system.DefaultRV32Config.fir@209815.6]
  wire [3:0] _T_1736; // @[Monitor.scala 645:61:freechips.rocketchip.system.DefaultRV32Config.fir@209816.6]
  wire [4:0] _T_1737; // @[Monitor.scala 646:49:freechips.rocketchip.system.DefaultRV32Config.fir@209818.6]
  wire [4:0] _T_1738; // @[Monitor.scala 646:57:freechips.rocketchip.system.DefaultRV32Config.fir@209819.6]
  wire [3:0] _GEN_80; // @[Monitor.scala 647:72:freechips.rocketchip.system.DefaultRV32Config.fir@209821.6]
  wire [4:0] _T_1739; // @[Monitor.scala 647:72:freechips.rocketchip.system.DefaultRV32Config.fir@209821.6]
  wire [3:0] a_opcodes_set_interm; // @[Monitor.scala 643:72:freechips.rocketchip.system.DefaultRV32Config.fir@209812.4]
  wire [34:0] _GEN_81; // @[Monitor.scala 647:47:freechips.rocketchip.system.DefaultRV32Config.fir@209822.6]
  wire [34:0] _T_1740; // @[Monitor.scala 647:47:freechips.rocketchip.system.DefaultRV32Config.fir@209822.6]
  wire [4:0] _T_1741; // @[Monitor.scala 648:68:freechips.rocketchip.system.DefaultRV32Config.fir@209824.6]
  wire [4:0] a_sizes_set_interm; // @[Monitor.scala 643:72:freechips.rocketchip.system.DefaultRV32Config.fir@209812.4]
  wire [35:0] _GEN_82; // @[Monitor.scala 648:43:freechips.rocketchip.system.DefaultRV32Config.fir@209825.6]
  wire [35:0] _T_1742; // @[Monitor.scala 648:43:freechips.rocketchip.system.DefaultRV32Config.fir@209825.6]
  wire [2:0] _T_1743; // @[Monitor.scala 649:26:freechips.rocketchip.system.DefaultRV32Config.fir@209827.6]
  wire  _T_1745; // @[Monitor.scala 649:17:freechips.rocketchip.system.DefaultRV32Config.fir@209829.6]
  wire  _T_1747; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@209831.6]
  wire  _T_1748; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@209832.6]
  wire [3:0] _GEN_27; // @[Monitor.scala 643:72:freechips.rocketchip.system.DefaultRV32Config.fir@209812.4]
  wire [34:0] _GEN_30; // @[Monitor.scala 643:72:freechips.rocketchip.system.DefaultRV32Config.fir@209812.4]
  wire [35:0] _GEN_31; // @[Monitor.scala 643:72:freechips.rocketchip.system.DefaultRV32Config.fir@209812.4]
  wire  _T_1751; // @[Monitor.scala 660:27:freechips.rocketchip.system.DefaultRV32Config.fir@209846.4]
  wire  _T_1753; // @[Monitor.scala 660:75:freechips.rocketchip.system.DefaultRV32Config.fir@209848.4]
  wire  _T_1754; // @[Monitor.scala 660:72:freechips.rocketchip.system.DefaultRV32Config.fir@209849.4]
  wire [3:0] _T_1755; // @[OneHot.scala 58:35:freechips.rocketchip.system.DefaultRV32Config.fir@209851.6]
  wire [46:0] _GEN_84; // @[Monitor.scala 662:76:freechips.rocketchip.system.DefaultRV32Config.fir@209858.6]
  wire [46:0] _T_1761; // @[Monitor.scala 662:76:freechips.rocketchip.system.DefaultRV32Config.fir@209858.6]
  wire [46:0] _GEN_85; // @[Monitor.scala 663:72:freechips.rocketchip.system.DefaultRV32Config.fir@209865.6]
  wire [46:0] _T_1767; // @[Monitor.scala 663:72:freechips.rocketchip.system.DefaultRV32Config.fir@209865.6]
  wire [3:0] _GEN_32; // @[Monitor.scala 660:91:freechips.rocketchip.system.DefaultRV32Config.fir@209850.4]
  wire [46:0] _GEN_33; // @[Monitor.scala 660:91:freechips.rocketchip.system.DefaultRV32Config.fir@209850.4]
  wire [46:0] _GEN_34; // @[Monitor.scala 660:91:freechips.rocketchip.system.DefaultRV32Config.fir@209850.4]
  wire  _T_1768; // @[Monitor.scala 665:26:freechips.rocketchip.system.DefaultRV32Config.fir@209868.4]
  wire  _T_1771; // @[Monitor.scala 665:71:freechips.rocketchip.system.DefaultRV32Config.fir@209871.4]
  wire [2:0] _T_1772; // @[Monitor.scala 666:25:freechips.rocketchip.system.DefaultRV32Config.fir@209873.6]
  wire  _T_1774; // @[Monitor.scala 666:93:freechips.rocketchip.system.DefaultRV32Config.fir@209875.6]
  wire  _T_1775; // @[Monitor.scala 666:68:freechips.rocketchip.system.DefaultRV32Config.fir@209876.6]
  wire  _T_1776; // @[Monitor.scala 666:142:freechips.rocketchip.system.DefaultRV32Config.fir@209877.6]
  wire  _T_1777; // @[Monitor.scala 666:119:freechips.rocketchip.system.DefaultRV32Config.fir@209878.6]
  wire  _T_1778; // @[Monitor.scala 666:166:freechips.rocketchip.system.DefaultRV32Config.fir@209879.6]
  wire  _T_1779; // @[Monitor.scala 666:49:freechips.rocketchip.system.DefaultRV32Config.fir@209880.6]
  wire  _T_1781; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@209882.6]
  wire  _T_1782; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@209883.6]
  wire [3:0] a_opcode_lookup; // @[:freechips.rocketchip.system.DefaultRV32Config.fir@209765.4 :freechips.rocketchip.system.DefaultRV32Config.fir@209766.4 Monitor.scala 629:21:freechips.rocketchip.system.DefaultRV32Config.fir@209775.4]
  wire [2:0] _GEN_37; // @[Monitor.scala 667:37:freechips.rocketchip.system.DefaultRV32Config.fir@209889.6]
  wire [2:0] _GEN_38; // @[Monitor.scala 667:37:freechips.rocketchip.system.DefaultRV32Config.fir@209889.6]
  wire [2:0] _GEN_39; // @[Monitor.scala 667:37:freechips.rocketchip.system.DefaultRV32Config.fir@209889.6]
  wire [2:0] _GEN_40; // @[Monitor.scala 667:37:freechips.rocketchip.system.DefaultRV32Config.fir@209889.6]
  wire [2:0] _GEN_41; // @[Monitor.scala 667:37:freechips.rocketchip.system.DefaultRV32Config.fir@209889.6]
  wire [2:0] _GEN_42; // @[Monitor.scala 667:37:freechips.rocketchip.system.DefaultRV32Config.fir@209889.6]
  wire  _T_1784; // @[Monitor.scala 667:37:freechips.rocketchip.system.DefaultRV32Config.fir@209889.6]
  wire [2:0] _GEN_49; // @[Monitor.scala 667:96:freechips.rocketchip.system.DefaultRV32Config.fir@209891.6]
  wire [2:0] _GEN_50; // @[Monitor.scala 667:96:freechips.rocketchip.system.DefaultRV32Config.fir@209891.6]
  wire  _T_1786; // @[Monitor.scala 667:96:freechips.rocketchip.system.DefaultRV32Config.fir@209891.6]
  wire  _T_1787; // @[Monitor.scala 667:71:freechips.rocketchip.system.DefaultRV32Config.fir@209892.6]
  wire [2:0] _GEN_53; // @[Monitor.scala 668:60:freechips.rocketchip.system.DefaultRV32Config.fir@209893.6]
  wire [2:0] _GEN_54; // @[Monitor.scala 668:60:freechips.rocketchip.system.DefaultRV32Config.fir@209893.6]
  wire [2:0] _GEN_55; // @[Monitor.scala 668:60:freechips.rocketchip.system.DefaultRV32Config.fir@209893.6]
  wire [2:0] _GEN_56; // @[Monitor.scala 668:60:freechips.rocketchip.system.DefaultRV32Config.fir@209893.6]
  wire [2:0] _GEN_57; // @[Monitor.scala 668:60:freechips.rocketchip.system.DefaultRV32Config.fir@209893.6]
  wire [2:0] _GEN_58; // @[Monitor.scala 668:60:freechips.rocketchip.system.DefaultRV32Config.fir@209893.6]
  wire  _T_1788; // @[Monitor.scala 668:60:freechips.rocketchip.system.DefaultRV32Config.fir@209893.6]
  wire [2:0] _GEN_65; // @[Monitor.scala 668:124:freechips.rocketchip.system.DefaultRV32Config.fir@209894.6]
  wire [2:0] _GEN_66; // @[Monitor.scala 668:124:freechips.rocketchip.system.DefaultRV32Config.fir@209894.6]
  wire  _T_1789; // @[Monitor.scala 668:124:freechips.rocketchip.system.DefaultRV32Config.fir@209894.6]
  wire  _T_1790; // @[Monitor.scala 668:99:freechips.rocketchip.system.DefaultRV32Config.fir@209895.6]
  wire  _T_1791; // @[Monitor.scala 668:34:freechips.rocketchip.system.DefaultRV32Config.fir@209896.6]
  wire  _T_1792; // @[Monitor.scala 668:15:freechips.rocketchip.system.DefaultRV32Config.fir@209897.6]
  wire  _T_1794; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@209899.6]
  wire  _T_1795; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@209900.6]
  wire [7:0] a_size_lookup; // @[:freechips.rocketchip.system.DefaultRV32Config.fir@209776.4 :freechips.rocketchip.system.DefaultRV32Config.fir@209777.4 Monitor.scala 633:19:freechips.rocketchip.system.DefaultRV32Config.fir@209786.4]
  wire [7:0] _GEN_86; // @[Monitor.scala 670:34:freechips.rocketchip.system.DefaultRV32Config.fir@209905.6]
  wire  _T_1796; // @[Monitor.scala 670:34:freechips.rocketchip.system.DefaultRV32Config.fir@209905.6]
  wire  _T_1798; // @[Monitor.scala 670:72:freechips.rocketchip.system.DefaultRV32Config.fir@209907.6]
  wire  _T_1799; // @[Monitor.scala 670:53:freechips.rocketchip.system.DefaultRV32Config.fir@209908.6]
  wire  _T_1801; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@209910.6]
  wire  _T_1802; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@209911.6]
  wire  _T_1804; // @[Monitor.scala 672:36:freechips.rocketchip.system.DefaultRV32Config.fir@209918.4]
  wire  _T_1805; // @[Monitor.scala 672:47:freechips.rocketchip.system.DefaultRV32Config.fir@209919.4]
  wire  _T_1807; // @[Monitor.scala 672:65:freechips.rocketchip.system.DefaultRV32Config.fir@209921.4]
  wire  _T_1809; // @[Monitor.scala 672:116:freechips.rocketchip.system.DefaultRV32Config.fir@209923.4]
  wire  _T_1810; // @[Monitor.scala 673:15:freechips.rocketchip.system.DefaultRV32Config.fir@209925.6]
  wire  _T_1811; // @[Monitor.scala 673:32:freechips.rocketchip.system.DefaultRV32Config.fir@209926.6]
  wire  _T_1813; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@209928.6]
  wire  _T_1814; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@209929.6]
  wire [2:0] a_set; // @[:freechips.rocketchip.system.DefaultRV32Config.fir@209759.4 :freechips.rocketchip.system.DefaultRV32Config.fir@209760.4 Monitor.scala 644:13:freechips.rocketchip.system.DefaultRV32Config.fir@209814.6]
  wire [2:0] d_clr; // @[:freechips.rocketchip.system.DefaultRV32Config.fir@209838.4 :freechips.rocketchip.system.DefaultRV32Config.fir@209839.4 Monitor.scala 661:13:freechips.rocketchip.system.DefaultRV32Config.fir@209852.6]
  wire  _T_1815; // @[Monitor.scala 677:20:freechips.rocketchip.system.DefaultRV32Config.fir@209935.4]
  wire  _T_1816; // @[Monitor.scala 677:40:freechips.rocketchip.system.DefaultRV32Config.fir@209936.4]
  wire  _T_1817; // @[Monitor.scala 677:33:freechips.rocketchip.system.DefaultRV32Config.fir@209937.4]
  wire  _T_1818; // @[Monitor.scala 677:30:freechips.rocketchip.system.DefaultRV32Config.fir@209938.4]
  wire  _T_1820; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@209940.4]
  wire  _T_1821; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@209941.4]
  wire [2:0] _T_1822; // @[Monitor.scala 680:27:freechips.rocketchip.system.DefaultRV32Config.fir@209946.4]
  wire [2:0] _T_1823; // @[Monitor.scala 680:38:freechips.rocketchip.system.DefaultRV32Config.fir@209947.4]
  wire [2:0] _T_1824; // @[Monitor.scala 680:36:freechips.rocketchip.system.DefaultRV32Config.fir@209948.4]
  wire [11:0] a_opcodes_set; // @[:freechips.rocketchip.system.DefaultRV32Config.fir@209761.4 :freechips.rocketchip.system.DefaultRV32Config.fir@209762.4 Monitor.scala 647:21:freechips.rocketchip.system.DefaultRV32Config.fir@209823.6]
  wire [11:0] _T_1825; // @[Monitor.scala 681:43:freechips.rocketchip.system.DefaultRV32Config.fir@209950.4]
  wire [11:0] d_opcodes_clr; // @[:freechips.rocketchip.system.DefaultRV32Config.fir@209840.4 :freechips.rocketchip.system.DefaultRV32Config.fir@209841.4 Monitor.scala 662:21:freechips.rocketchip.system.DefaultRV32Config.fir@209859.6]
  wire [11:0] _T_1826; // @[Monitor.scala 681:62:freechips.rocketchip.system.DefaultRV32Config.fir@209951.4]
  wire [11:0] _T_1827; // @[Monitor.scala 681:60:freechips.rocketchip.system.DefaultRV32Config.fir@209952.4]
  wire [23:0] a_sizes_set; // @[:freechips.rocketchip.system.DefaultRV32Config.fir@209763.4 :freechips.rocketchip.system.DefaultRV32Config.fir@209764.4 Monitor.scala 648:19:freechips.rocketchip.system.DefaultRV32Config.fir@209826.6]
  wire [23:0] _T_1828; // @[Monitor.scala 682:39:freechips.rocketchip.system.DefaultRV32Config.fir@209954.4]
  wire [23:0] d_sizes_clr; // @[:freechips.rocketchip.system.DefaultRV32Config.fir@209842.4 :freechips.rocketchip.system.DefaultRV32Config.fir@209843.4 Monitor.scala 663:19:freechips.rocketchip.system.DefaultRV32Config.fir@209866.6]
  wire [23:0] _T_1829; // @[Monitor.scala 682:56:freechips.rocketchip.system.DefaultRV32Config.fir@209955.4]
  wire [23:0] _T_1830; // @[Monitor.scala 682:54:freechips.rocketchip.system.DefaultRV32Config.fir@209956.4]
  reg [31:0] _T_1831; // @[Monitor.scala 684:27:freechips.rocketchip.system.DefaultRV32Config.fir@209958.4]
  wire  _T_1832; // @[Monitor.scala 687:26:freechips.rocketchip.system.DefaultRV32Config.fir@209961.4]
  wire  _T_1833; // @[Monitor.scala 687:16:freechips.rocketchip.system.DefaultRV32Config.fir@209962.4]
  wire  _T_1834; // @[Monitor.scala 687:39:freechips.rocketchip.system.DefaultRV32Config.fir@209963.4]
  wire  _T_1835; // @[Monitor.scala 687:30:freechips.rocketchip.system.DefaultRV32Config.fir@209964.4]
  wire  _T_1836; // @[Monitor.scala 687:59:freechips.rocketchip.system.DefaultRV32Config.fir@209965.4]
  wire  _T_1837; // @[Monitor.scala 687:47:freechips.rocketchip.system.DefaultRV32Config.fir@209966.4]
  wire  _T_1839; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@209968.4]
  wire  _T_1840; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@209969.4]
  wire [31:0] _T_1842; // @[Monitor.scala 689:26:freechips.rocketchip.system.DefaultRV32Config.fir@209975.4]
  wire  _T_1845; // @[Monitor.scala 690:27:freechips.rocketchip.system.DefaultRV32Config.fir@209979.4]
  reg [3:0] _T_1846; // @[Monitor.scala 694:27:freechips.rocketchip.system.DefaultRV32Config.fir@209983.4]
  reg [9:0] _T_1855; // @[Edges.scala 230:27:freechips.rocketchip.system.DefaultRV32Config.fir@209992.4]
  wire [9:0] _T_1857; // @[Edges.scala 231:28:freechips.rocketchip.system.DefaultRV32Config.fir@209994.4]
  wire  _T_1858; // @[Edges.scala 232:25:freechips.rocketchip.system.DefaultRV32Config.fir@209995.4]
  wire  _T_1868; // @[Monitor.scala 700:27:freechips.rocketchip.system.DefaultRV32Config.fir@210009.4]
  wire  _T_1871; // @[Edges.scala 72:43:freechips.rocketchip.system.DefaultRV32Config.fir@210012.4]
  wire  _T_1872; // @[Edges.scala 72:40:freechips.rocketchip.system.DefaultRV32Config.fir@210013.4]
  wire  _T_1873; // @[Monitor.scala 700:38:freechips.rocketchip.system.DefaultRV32Config.fir@210014.4]
  wire [3:0] _T_1874; // @[OneHot.scala 58:35:freechips.rocketchip.system.DefaultRV32Config.fir@210016.6]
  wire [3:0] _T_1875; // @[Monitor.scala 702:23:freechips.rocketchip.system.DefaultRV32Config.fir@210018.6]
  wire  _T_1877; // @[Monitor.scala 702:14:freechips.rocketchip.system.DefaultRV32Config.fir@210020.6]
  wire  _T_1879; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@210022.6]
  wire  _T_1880; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@210023.6]
  wire [3:0] _GEN_69; // @[Monitor.scala 700:72:freechips.rocketchip.system.DefaultRV32Config.fir@210015.4]
  wire  _T_1882; // @[Decoupled.scala 40:37:freechips.rocketchip.system.DefaultRV32Config.fir@210031.4]
  wire [3:0] _T_1885; // @[OneHot.scala 58:35:freechips.rocketchip.system.DefaultRV32Config.fir@210035.6]
  wire [3:0] _T_1886; // @[Monitor.scala 708:24:freechips.rocketchip.system.DefaultRV32Config.fir@210037.6]
  wire [3:0] _T_1887; // @[Monitor.scala 708:35:freechips.rocketchip.system.DefaultRV32Config.fir@210038.6]
  wire  _T_1890; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@210041.6]
  wire  _T_1891; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@210042.6]
  wire [3:0] _GEN_70; // @[Monitor.scala 706:73:freechips.rocketchip.system.DefaultRV32Config.fir@210034.4]
  wire [3:0] _T_1892; // @[Monitor.scala 713:27:freechips.rocketchip.system.DefaultRV32Config.fir@210048.4]
  wire [3:0] _T_1893; // @[Monitor.scala 713:38:freechips.rocketchip.system.DefaultRV32Config.fir@210049.4]
  wire [3:0] _T_1894; // @[Monitor.scala 713:36:freechips.rocketchip.system.DefaultRV32Config.fir@210050.4]
  wire  _GEN_87; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@207244.10]
  wire  _GEN_103; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@207373.10]
  wire  _GEN_121; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@207513.10]
  wire  _GEN_133; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@207620.10]
  wire  _GEN_143; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@207719.10]
  wire  _GEN_153; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@207810.10]
  wire  _GEN_163; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@207899.10]
  wire  _GEN_173; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@207988.10]
  wire  _GEN_185; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@208057.10]
  wire  _GEN_195; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@208099.10]
  wire  _GEN_205; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@208157.10]
  wire  _GEN_215; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@208216.10]
  wire  _GEN_221; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@208251.10]
  wire  _GEN_227; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@208287.10]
  wire  _GEN_233; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@208486.10]
  wire  _GEN_247; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@208541.10]
  wire  _GEN_261; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@208596.10]
  wire  _GEN_273; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@208643.10]
  wire  _GEN_285; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@208692.10]
  wire  _GEN_295; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@208739.10]
  wire  _GEN_305; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@208786.10]
  wire  _GEN_317; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@208942.10]
  wire  _GEN_327; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@208990.10]
  wire  _GEN_337; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@209079.10]
  wire  _GEN_349; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@209199.10]
  wire  _GEN_361; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@209262.10]
  wire  _GEN_369; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@209302.10]
  wire  _GEN_377; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@209334.10]
  plusarg_reader #(.FORMAT("tilelink_timeout=%d"), .DEFAULT(0), .WIDTH(32)) plusarg_reader ( // @[PlusArg.scala 80:11:freechips.rocketchip.system.DefaultRV32Config.fir@209959.4]
    .out(plusarg_reader_out)
  );
  assign _T_4 = io_in_a_bits_source == 2'h0; // @[Parameters.scala 47:9:freechips.rocketchip.system.DefaultRV32Config.fir@207107.6]
  assign _T_5 = io_in_a_bits_source == 2'h1; // @[Parameters.scala 47:9:freechips.rocketchip.system.DefaultRV32Config.fir@207108.6]
  assign _T_6 = io_in_a_bits_source == 2'h2; // @[Parameters.scala 47:9:freechips.rocketchip.system.DefaultRV32Config.fir@207109.6]
  assign _T_8 = _T_4 | _T_5; // @[Parameters.scala 924:46:freechips.rocketchip.system.DefaultRV32Config.fir@207115.6]
  assign _T_9 = _T_8 | _T_6; // @[Parameters.scala 924:46:freechips.rocketchip.system.DefaultRV32Config.fir@207116.6]
  assign _T_11 = 27'hfff << io_in_a_bits_size; // @[package.scala 207:77:freechips.rocketchip.system.DefaultRV32Config.fir@207118.6]
  assign _T_13 = ~_T_11[11:0]; // @[package.scala 207:46:freechips.rocketchip.system.DefaultRV32Config.fir@207120.6]
  assign _GEN_71 = {{20'd0}, _T_13}; // @[Edges.scala 22:16:freechips.rocketchip.system.DefaultRV32Config.fir@207121.6]
  assign _T_14 = io_in_a_bits_address & _GEN_71; // @[Edges.scala 22:16:freechips.rocketchip.system.DefaultRV32Config.fir@207121.6]
  assign _T_15 = _T_14 == 32'h0; // @[Edges.scala 22:24:freechips.rocketchip.system.DefaultRV32Config.fir@207122.6]
  assign _T_18 = 2'h1 << io_in_a_bits_size[0]; // @[OneHot.scala 65:12:freechips.rocketchip.system.DefaultRV32Config.fir@207125.6]
  assign _T_20 = _T_18 | 2'h1; // @[Misc.scala 201:81:freechips.rocketchip.system.DefaultRV32Config.fir@207127.6]
  assign _T_21 = io_in_a_bits_size >= 4'h2; // @[Misc.scala 205:21:freechips.rocketchip.system.DefaultRV32Config.fir@207128.6]
  assign _T_24 = ~io_in_a_bits_address[1]; // @[Misc.scala 210:20:freechips.rocketchip.system.DefaultRV32Config.fir@207131.6]
  assign _T_26 = _T_20[1] & _T_24; // @[Misc.scala 214:38:freechips.rocketchip.system.DefaultRV32Config.fir@207133.6]
  assign _T_27 = _T_21 | _T_26; // @[Misc.scala 214:29:freechips.rocketchip.system.DefaultRV32Config.fir@207134.6]
  assign _T_29 = _T_20[1] & io_in_a_bits_address[1]; // @[Misc.scala 214:38:freechips.rocketchip.system.DefaultRV32Config.fir@207136.6]
  assign _T_30 = _T_21 | _T_29; // @[Misc.scala 214:29:freechips.rocketchip.system.DefaultRV32Config.fir@207137.6]
  assign _T_33 = ~io_in_a_bits_address[0]; // @[Misc.scala 210:20:freechips.rocketchip.system.DefaultRV32Config.fir@207140.6]
  assign _T_34 = _T_24 & _T_33; // @[Misc.scala 213:27:freechips.rocketchip.system.DefaultRV32Config.fir@207141.6]
  assign _T_35 = _T_20[0] & _T_34; // @[Misc.scala 214:38:freechips.rocketchip.system.DefaultRV32Config.fir@207142.6]
  assign _T_36 = _T_27 | _T_35; // @[Misc.scala 214:29:freechips.rocketchip.system.DefaultRV32Config.fir@207143.6]
  assign _T_37 = _T_24 & io_in_a_bits_address[0]; // @[Misc.scala 213:27:freechips.rocketchip.system.DefaultRV32Config.fir@207144.6]
  assign _T_38 = _T_20[0] & _T_37; // @[Misc.scala 214:38:freechips.rocketchip.system.DefaultRV32Config.fir@207145.6]
  assign _T_39 = _T_27 | _T_38; // @[Misc.scala 214:29:freechips.rocketchip.system.DefaultRV32Config.fir@207146.6]
  assign _T_40 = io_in_a_bits_address[1] & _T_33; // @[Misc.scala 213:27:freechips.rocketchip.system.DefaultRV32Config.fir@207147.6]
  assign _T_41 = _T_20[0] & _T_40; // @[Misc.scala 214:38:freechips.rocketchip.system.DefaultRV32Config.fir@207148.6]
  assign _T_42 = _T_30 | _T_41; // @[Misc.scala 214:29:freechips.rocketchip.system.DefaultRV32Config.fir@207149.6]
  assign _T_43 = io_in_a_bits_address[1] & io_in_a_bits_address[0]; // @[Misc.scala 213:27:freechips.rocketchip.system.DefaultRV32Config.fir@207150.6]
  assign _T_44 = _T_20[0] & _T_43; // @[Misc.scala 214:38:freechips.rocketchip.system.DefaultRV32Config.fir@207151.6]
  assign _T_45 = _T_30 | _T_44; // @[Misc.scala 214:29:freechips.rocketchip.system.DefaultRV32Config.fir@207152.6]
  assign _T_48 = {_T_45,_T_42,_T_39,_T_36}; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@207155.6]
  assign _T_52 = {1'b0,$signed(io_in_a_bits_address)}; // @[Parameters.scala 137:49:freechips.rocketchip.system.DefaultRV32Config.fir@207159.6]
  assign _T_78 = io_in_a_bits_opcode == 3'h6; // @[Monitor.scala 79:25:freechips.rocketchip.system.DefaultRV32Config.fir@207189.6]
  assign _T_83 = $signed(_T_52) & -33'sh1000; // @[Parameters.scala 137:52:freechips.rocketchip.system.DefaultRV32Config.fir@207195.8]
  assign _T_84 = $signed(_T_83) == 33'sh0; // @[Parameters.scala 137:67:freechips.rocketchip.system.DefaultRV32Config.fir@207196.8]
  assign _T_85 = io_in_a_bits_address ^ 32'h3000; // @[Parameters.scala 137:31:freechips.rocketchip.system.DefaultRV32Config.fir@207197.8]
  assign _T_86 = {1'b0,$signed(_T_85)}; // @[Parameters.scala 137:49:freechips.rocketchip.system.DefaultRV32Config.fir@207198.8]
  assign _T_88 = $signed(_T_86) & -33'sh1000; // @[Parameters.scala 137:52:freechips.rocketchip.system.DefaultRV32Config.fir@207200.8]
  assign _T_89 = $signed(_T_88) == 33'sh0; // @[Parameters.scala 137:67:freechips.rocketchip.system.DefaultRV32Config.fir@207201.8]
  assign _T_90 = io_in_a_bits_address ^ 32'h10000; // @[Parameters.scala 137:31:freechips.rocketchip.system.DefaultRV32Config.fir@207202.8]
  assign _T_91 = {1'b0,$signed(_T_90)}; // @[Parameters.scala 137:49:freechips.rocketchip.system.DefaultRV32Config.fir@207203.8]
  assign _T_93 = $signed(_T_91) & -33'sh10000; // @[Parameters.scala 137:52:freechips.rocketchip.system.DefaultRV32Config.fir@207205.8]
  assign _T_94 = $signed(_T_93) == 33'sh0; // @[Parameters.scala 137:67:freechips.rocketchip.system.DefaultRV32Config.fir@207206.8]
  assign _T_95 = io_in_a_bits_address ^ 32'h2000000; // @[Parameters.scala 137:31:freechips.rocketchip.system.DefaultRV32Config.fir@207207.8]
  assign _T_96 = {1'b0,$signed(_T_95)}; // @[Parameters.scala 137:49:freechips.rocketchip.system.DefaultRV32Config.fir@207208.8]
  assign _T_98 = $signed(_T_96) & -33'sh10000; // @[Parameters.scala 137:52:freechips.rocketchip.system.DefaultRV32Config.fir@207210.8]
  assign _T_99 = $signed(_T_98) == 33'sh0; // @[Parameters.scala 137:67:freechips.rocketchip.system.DefaultRV32Config.fir@207211.8]
  assign _T_100 = io_in_a_bits_address ^ 32'hc000000; // @[Parameters.scala 137:31:freechips.rocketchip.system.DefaultRV32Config.fir@207212.8]
  assign _T_101 = {1'b0,$signed(_T_100)}; // @[Parameters.scala 137:49:freechips.rocketchip.system.DefaultRV32Config.fir@207213.8]
  assign _T_103 = $signed(_T_101) & -33'sh4000000; // @[Parameters.scala 137:52:freechips.rocketchip.system.DefaultRV32Config.fir@207215.8]
  assign _T_104 = $signed(_T_103) == 33'sh0; // @[Parameters.scala 137:67:freechips.rocketchip.system.DefaultRV32Config.fir@207216.8]
  assign _T_105 = io_in_a_bits_address ^ 32'h60000000; // @[Parameters.scala 137:31:freechips.rocketchip.system.DefaultRV32Config.fir@207217.8]
  assign _T_106 = {1'b0,$signed(_T_105)}; // @[Parameters.scala 137:49:freechips.rocketchip.system.DefaultRV32Config.fir@207218.8]
  assign _T_108 = $signed(_T_106) & -33'sh20000000; // @[Parameters.scala 137:52:freechips.rocketchip.system.DefaultRV32Config.fir@207220.8]
  assign _T_109 = $signed(_T_108) == 33'sh0; // @[Parameters.scala 137:67:freechips.rocketchip.system.DefaultRV32Config.fir@207221.8]
  assign _T_110 = _T_84 | _T_89; // @[Parameters.scala 552:42:freechips.rocketchip.system.DefaultRV32Config.fir@207222.8]
  assign _T_117 = io_in_a_bits_size <= 4'h6; // @[Parameters.scala 93:42:freechips.rocketchip.system.DefaultRV32Config.fir@207229.8]
  assign _T_120 = io_in_a_bits_address ^ 32'h80000000; // @[Parameters.scala 137:31:freechips.rocketchip.system.DefaultRV32Config.fir@207232.8]
  assign _T_121 = {1'b0,$signed(_T_120)}; // @[Parameters.scala 137:49:freechips.rocketchip.system.DefaultRV32Config.fir@207233.8]
  assign _T_123 = $signed(_T_121) & -33'sh10000000; // @[Parameters.scala 137:52:freechips.rocketchip.system.DefaultRV32Config.fir@207235.8]
  assign _T_124 = $signed(_T_123) == 33'sh0; // @[Parameters.scala 137:67:freechips.rocketchip.system.DefaultRV32Config.fir@207236.8]
  assign _T_125 = _T_117 & _T_124; // @[Parameters.scala 551:56:freechips.rocketchip.system.DefaultRV32Config.fir@207237.8]
  assign _T_129 = _T_125 | reset; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@207241.8]
  assign _T_130 = ~_T_129; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@207242.8]
  assign _T_135 = 4'h6 == io_in_a_bits_size; // @[Parameters.scala 92:48:freechips.rocketchip.system.DefaultRV32Config.fir@207255.8]
  assign _T_136 = _T_4 & _T_135; // @[Mux.scala 27:72:freechips.rocketchip.system.DefaultRV32Config.fir@207256.8]
  assign _T_143 = _T_136 | reset; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@207264.8]
  assign _T_144 = ~_T_143; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@207265.8]
  assign _T_146 = _T_9 | reset; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@207271.8]
  assign _T_147 = ~_T_146; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@207272.8]
  assign _T_150 = _T_21 | reset; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@207279.8]
  assign _T_151 = ~_T_150; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@207280.8]
  assign _T_153 = _T_15 | reset; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@207286.8]
  assign _T_154 = ~_T_153; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@207287.8]
  assign _T_155 = io_in_a_bits_param <= 3'h2; // @[Bundles.scala 110:27:freechips.rocketchip.system.DefaultRV32Config.fir@207292.8]
  assign _T_157 = _T_155 | reset; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@207294.8]
  assign _T_158 = ~_T_157; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@207295.8]
  assign _T_159 = ~io_in_a_bits_mask; // @[Monitor.scala 86:18:freechips.rocketchip.system.DefaultRV32Config.fir@207300.8]
  assign _T_160 = _T_159 == 4'h0; // @[Monitor.scala 86:31:freechips.rocketchip.system.DefaultRV32Config.fir@207301.8]
  assign _T_162 = _T_160 | reset; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@207303.8]
  assign _T_163 = ~_T_162; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@207304.8]
  assign _T_164 = ~io_in_a_bits_corrupt; // @[Monitor.scala 87:18:freechips.rocketchip.system.DefaultRV32Config.fir@207309.8]
  assign _T_166 = _T_164 | reset; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@207311.8]
  assign _T_167 = ~_T_166; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@207312.8]
  assign _T_168 = io_in_a_bits_opcode == 3'h7; // @[Monitor.scala 90:25:freechips.rocketchip.system.DefaultRV32Config.fir@207318.6]
  assign _T_249 = io_in_a_bits_param != 3'h0; // @[Monitor.scala 97:31:freechips.rocketchip.system.DefaultRV32Config.fir@207429.8]
  assign _T_251 = _T_249 | reset; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@207431.8]
  assign _T_252 = ~_T_251; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@207432.8]
  assign _T_262 = io_in_a_bits_opcode == 3'h4; // @[Monitor.scala 102:25:freechips.rocketchip.system.DefaultRV32Config.fir@207455.6]
  assign _T_264 = io_in_a_bits_size <= 4'hc; // @[Parameters.scala 93:42:freechips.rocketchip.system.DefaultRV32Config.fir@207458.8]
  assign _T_272 = _T_264 & _T_89; // @[Parameters.scala 551:56:freechips.rocketchip.system.DefaultRV32Config.fir@207466.8]
  assign _T_307 = _T_84 | _T_94; // @[Parameters.scala 552:42:freechips.rocketchip.system.DefaultRV32Config.fir@207501.8]
  assign _T_308 = _T_307 | _T_99; // @[Parameters.scala 552:42:freechips.rocketchip.system.DefaultRV32Config.fir@207502.8]
  assign _T_309 = _T_308 | _T_104; // @[Parameters.scala 552:42:freechips.rocketchip.system.DefaultRV32Config.fir@207503.8]
  assign _T_310 = _T_309 | _T_109; // @[Parameters.scala 552:42:freechips.rocketchip.system.DefaultRV32Config.fir@207504.8]
  assign _T_311 = _T_310 | _T_124; // @[Parameters.scala 552:42:freechips.rocketchip.system.DefaultRV32Config.fir@207505.8]
  assign _T_312 = _T_117 & _T_311; // @[Parameters.scala 551:56:freechips.rocketchip.system.DefaultRV32Config.fir@207506.8]
  assign _T_314 = _T_272 | _T_312; // @[Parameters.scala 553:30:freechips.rocketchip.system.DefaultRV32Config.fir@207508.8]
  assign _T_316 = _T_314 | reset; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@207510.8]
  assign _T_317 = ~_T_316; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@207511.8]
  assign _T_324 = io_in_a_bits_param == 3'h0; // @[Monitor.scala 106:31:freechips.rocketchip.system.DefaultRV32Config.fir@207530.8]
  assign _T_326 = _T_324 | reset; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@207532.8]
  assign _T_327 = ~_T_326; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@207533.8]
  assign _T_328 = io_in_a_bits_mask == _T_48; // @[Monitor.scala 107:30:freechips.rocketchip.system.DefaultRV32Config.fir@207538.8]
  assign _T_330 = _T_328 | reset; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@207540.8]
  assign _T_331 = ~_T_330; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@207541.8]
  assign _T_336 = io_in_a_bits_opcode == 3'h0; // @[Monitor.scala 111:25:freechips.rocketchip.system.DefaultRV32Config.fir@207555.6]
  assign _T_371 = _T_84 | _T_99; // @[Parameters.scala 552:42:freechips.rocketchip.system.DefaultRV32Config.fir@207591.8]
  assign _T_372 = _T_371 | _T_104; // @[Parameters.scala 552:42:freechips.rocketchip.system.DefaultRV32Config.fir@207592.8]
  assign _T_373 = _T_372 | _T_124; // @[Parameters.scala 552:42:freechips.rocketchip.system.DefaultRV32Config.fir@207593.8]
  assign _T_374 = _T_117 & _T_373; // @[Parameters.scala 551:56:freechips.rocketchip.system.DefaultRV32Config.fir@207594.8]
  assign _T_383 = io_in_a_bits_size <= 4'h8; // @[Parameters.scala 93:42:freechips.rocketchip.system.DefaultRV32Config.fir@207603.8]
  assign _T_391 = _T_383 & _T_109; // @[Parameters.scala 551:56:freechips.rocketchip.system.DefaultRV32Config.fir@207611.8]
  assign _T_393 = _T_272 | _T_374; // @[Parameters.scala 553:30:freechips.rocketchip.system.DefaultRV32Config.fir@207613.8]
  assign _T_395 = _T_393 | _T_391; // @[Parameters.scala 553:30:freechips.rocketchip.system.DefaultRV32Config.fir@207615.8]
  assign _T_397 = _T_395 | reset; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@207617.8]
  assign _T_398 = ~_T_397; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@207618.8]
  assign _T_413 = io_in_a_bits_opcode == 3'h1; // @[Monitor.scala 119:25:freechips.rocketchip.system.DefaultRV32Config.fir@207654.6]
  assign _T_486 = ~_T_48; // @[Monitor.scala 124:33:freechips.rocketchip.system.DefaultRV32Config.fir@207744.8]
  assign _T_487 = io_in_a_bits_mask & _T_486; // @[Monitor.scala 124:31:freechips.rocketchip.system.DefaultRV32Config.fir@207745.8]
  assign _T_488 = _T_487 == 4'h0; // @[Monitor.scala 124:40:freechips.rocketchip.system.DefaultRV32Config.fir@207746.8]
  assign _T_490 = _T_488 | reset; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@207748.8]
  assign _T_491 = ~_T_490; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@207749.8]
  assign _T_492 = io_in_a_bits_opcode == 3'h2; // @[Monitor.scala 127:25:freechips.rocketchip.system.DefaultRV32Config.fir@207755.6]
  assign _T_494 = io_in_a_bits_size <= 4'h2; // @[Parameters.scala 93:42:freechips.rocketchip.system.DefaultRV32Config.fir@207758.8]
  assign _T_518 = _T_110 | _T_99; // @[Parameters.scala 552:42:freechips.rocketchip.system.DefaultRV32Config.fir@207782.8]
  assign _T_519 = _T_518 | _T_104; // @[Parameters.scala 552:42:freechips.rocketchip.system.DefaultRV32Config.fir@207783.8]
  assign _T_520 = _T_494 & _T_519; // @[Parameters.scala 551:56:freechips.rocketchip.system.DefaultRV32Config.fir@207784.8]
  assign _T_543 = _T_520 | reset; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@207807.8]
  assign _T_544 = ~_T_543; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@207808.8]
  assign _T_551 = io_in_a_bits_param <= 3'h4; // @[Bundles.scala 140:33:freechips.rocketchip.system.DefaultRV32Config.fir@207827.8]
  assign _T_553 = _T_551 | reset; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@207829.8]
  assign _T_554 = ~_T_553; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@207830.8]
  assign _T_559 = io_in_a_bits_opcode == 3'h3; // @[Monitor.scala 135:25:freechips.rocketchip.system.DefaultRV32Config.fir@207844.6]
  assign _T_618 = io_in_a_bits_param <= 3'h3; // @[Bundles.scala 147:30:freechips.rocketchip.system.DefaultRV32Config.fir@207916.8]
  assign _T_620 = _T_618 | reset; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@207918.8]
  assign _T_621 = ~_T_620; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@207919.8]
  assign _T_626 = io_in_a_bits_opcode == 3'h5; // @[Monitor.scala 143:25:freechips.rocketchip.system.DefaultRV32Config.fir@207933.6]
  assign _T_677 = _T_272 | reset; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@207985.8]
  assign _T_678 = ~_T_677; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@207986.8]
  assign _T_685 = io_in_a_bits_param <= 3'h1; // @[Bundles.scala 160:28:freechips.rocketchip.system.DefaultRV32Config.fir@208005.8]
  assign _T_687 = _T_685 | reset; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@208007.8]
  assign _T_688 = ~_T_687; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@208008.8]
  assign _T_697 = io_in_d_bits_opcode <= 3'h6; // @[Bundles.scala 44:24:freechips.rocketchip.system.DefaultRV32Config.fir@208032.6]
  assign _T_699 = _T_697 | reset; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@208034.6]
  assign _T_700 = ~_T_699; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@208035.6]
  assign _T_701 = io_in_d_bits_source == 2'h0; // @[Parameters.scala 47:9:freechips.rocketchip.system.DefaultRV32Config.fir@208040.6]
  assign _T_702 = io_in_d_bits_source == 2'h1; // @[Parameters.scala 47:9:freechips.rocketchip.system.DefaultRV32Config.fir@208041.6]
  assign _T_703 = io_in_d_bits_source == 2'h2; // @[Parameters.scala 47:9:freechips.rocketchip.system.DefaultRV32Config.fir@208042.6]
  assign _T_705 = _T_701 | _T_702; // @[Parameters.scala 924:46:freechips.rocketchip.system.DefaultRV32Config.fir@208048.6]
  assign _T_706 = _T_705 | _T_703; // @[Parameters.scala 924:46:freechips.rocketchip.system.DefaultRV32Config.fir@208049.6]
  assign _T_708 = io_in_d_bits_opcode == 3'h6; // @[Monitor.scala 307:25:freechips.rocketchip.system.DefaultRV32Config.fir@208051.6]
  assign _T_710 = _T_706 | reset; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@208054.8]
  assign _T_711 = ~_T_710; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@208055.8]
  assign _T_712 = io_in_d_bits_size >= 4'h2; // @[Monitor.scala 309:27:freechips.rocketchip.system.DefaultRV32Config.fir@208060.8]
  assign _T_714 = _T_712 | reset; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@208062.8]
  assign _T_715 = ~_T_714; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@208063.8]
  assign _T_716 = io_in_d_bits_param == 2'h0; // @[Monitor.scala 310:28:freechips.rocketchip.system.DefaultRV32Config.fir@208068.8]
  assign _T_718 = _T_716 | reset; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@208070.8]
  assign _T_719 = ~_T_718; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@208071.8]
  assign _T_720 = ~io_in_d_bits_corrupt; // @[Monitor.scala 311:15:freechips.rocketchip.system.DefaultRV32Config.fir@208076.8]
  assign _T_722 = _T_720 | reset; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@208078.8]
  assign _T_723 = ~_T_722; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@208079.8]
  assign _T_724 = ~io_in_d_bits_denied; // @[Monitor.scala 312:15:freechips.rocketchip.system.DefaultRV32Config.fir@208084.8]
  assign _T_726 = _T_724 | reset; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@208086.8]
  assign _T_727 = ~_T_726; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@208087.8]
  assign _T_728 = io_in_d_bits_opcode == 3'h4; // @[Monitor.scala 315:25:freechips.rocketchip.system.DefaultRV32Config.fir@208093.6]
  assign _T_739 = io_in_d_bits_param <= 2'h2; // @[Bundles.scala 104:26:freechips.rocketchip.system.DefaultRV32Config.fir@208117.8]
  assign _T_741 = _T_739 | reset; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@208119.8]
  assign _T_742 = ~_T_741; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@208120.8]
  assign _T_743 = io_in_d_bits_param != 2'h2; // @[Monitor.scala 320:28:freechips.rocketchip.system.DefaultRV32Config.fir@208125.8]
  assign _T_745 = _T_743 | reset; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@208127.8]
  assign _T_746 = ~_T_745; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@208128.8]
  assign _T_756 = io_in_d_bits_opcode == 3'h5; // @[Monitor.scala 325:25:freechips.rocketchip.system.DefaultRV32Config.fir@208151.6]
  assign _T_776 = _T_724 | io_in_d_bits_corrupt; // @[Monitor.scala 331:30:freechips.rocketchip.system.DefaultRV32Config.fir@208192.8]
  assign _T_778 = _T_776 | reset; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@208194.8]
  assign _T_779 = ~_T_778; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@208195.8]
  assign _T_785 = io_in_d_bits_opcode == 3'h0; // @[Monitor.scala 335:25:freechips.rocketchip.system.DefaultRV32Config.fir@208210.6]
  assign _T_802 = io_in_d_bits_opcode == 3'h1; // @[Monitor.scala 343:25:freechips.rocketchip.system.DefaultRV32Config.fir@208245.6]
  assign _T_820 = io_in_d_bits_opcode == 3'h2; // @[Monitor.scala 351:25:freechips.rocketchip.system.DefaultRV32Config.fir@208281.6]
  assign _T_837 = io_in_b_bits_opcode <= 3'h6; // @[Bundles.scala 42:24:freechips.rocketchip.system.DefaultRV32Config.fir@208318.6]
  assign _T_839 = _T_837 | reset; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@208320.6]
  assign _T_840 = ~_T_839; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@208321.6]
  assign _T_841 = io_in_b_bits_source == 2'h0; // @[Parameters.scala 47:9:freechips.rocketchip.system.DefaultRV32Config.fir@208326.6]
  assign _T_844 = {1'b0,$signed(io_in_b_bits_address)}; // @[Parameters.scala 137:49:freechips.rocketchip.system.DefaultRV32Config.fir@208329.6]
  assign _T_849 = io_in_b_bits_source == 2'h1; // @[Parameters.scala 47:9:freechips.rocketchip.system.DefaultRV32Config.fir@208334.6]
  assign _T_857 = io_in_b_bits_source == 2'h2; // @[Parameters.scala 47:9:freechips.rocketchip.system.DefaultRV32Config.fir@208342.6]
  assign _T_870 = io_in_b_bits_address ^ 32'h3000; // @[Parameters.scala 137:31:freechips.rocketchip.system.DefaultRV32Config.fir@208359.6]
  assign _T_871 = {1'b0,$signed(_T_870)}; // @[Parameters.scala 137:49:freechips.rocketchip.system.DefaultRV32Config.fir@208360.6]
  assign _T_873 = $signed(_T_871) & -33'sh1000; // @[Parameters.scala 137:52:freechips.rocketchip.system.DefaultRV32Config.fir@208362.6]
  assign _T_874 = $signed(_T_873) == 33'sh0; // @[Parameters.scala 137:67:freechips.rocketchip.system.DefaultRV32Config.fir@208363.6]
  assign _T_875 = io_in_b_bits_address ^ 32'hc000000; // @[Parameters.scala 137:31:freechips.rocketchip.system.DefaultRV32Config.fir@208364.6]
  assign _T_876 = {1'b0,$signed(_T_875)}; // @[Parameters.scala 137:49:freechips.rocketchip.system.DefaultRV32Config.fir@208365.6]
  assign _T_878 = $signed(_T_876) & -33'sh4000000; // @[Parameters.scala 137:52:freechips.rocketchip.system.DefaultRV32Config.fir@208367.6]
  assign _T_879 = $signed(_T_878) == 33'sh0; // @[Parameters.scala 137:67:freechips.rocketchip.system.DefaultRV32Config.fir@208368.6]
  assign _T_880 = io_in_b_bits_address ^ 32'h2000000; // @[Parameters.scala 137:31:freechips.rocketchip.system.DefaultRV32Config.fir@208369.6]
  assign _T_881 = {1'b0,$signed(_T_880)}; // @[Parameters.scala 137:49:freechips.rocketchip.system.DefaultRV32Config.fir@208370.6]
  assign _T_883 = $signed(_T_881) & -33'sh10000; // @[Parameters.scala 137:52:freechips.rocketchip.system.DefaultRV32Config.fir@208372.6]
  assign _T_884 = $signed(_T_883) == 33'sh0; // @[Parameters.scala 137:67:freechips.rocketchip.system.DefaultRV32Config.fir@208373.6]
  assign _T_888 = $signed(_T_844) & -33'sh1000; // @[Parameters.scala 137:52:freechips.rocketchip.system.DefaultRV32Config.fir@208377.6]
  assign _T_889 = $signed(_T_888) == 33'sh0; // @[Parameters.scala 137:67:freechips.rocketchip.system.DefaultRV32Config.fir@208378.6]
  assign _T_890 = io_in_b_bits_address ^ 32'h10000; // @[Parameters.scala 137:31:freechips.rocketchip.system.DefaultRV32Config.fir@208379.6]
  assign _T_891 = {1'b0,$signed(_T_890)}; // @[Parameters.scala 137:49:freechips.rocketchip.system.DefaultRV32Config.fir@208380.6]
  assign _T_893 = $signed(_T_891) & -33'sh10000; // @[Parameters.scala 137:52:freechips.rocketchip.system.DefaultRV32Config.fir@208382.6]
  assign _T_894 = $signed(_T_893) == 33'sh0; // @[Parameters.scala 137:67:freechips.rocketchip.system.DefaultRV32Config.fir@208383.6]
  assign _T_895 = io_in_b_bits_address ^ 32'h80000000; // @[Parameters.scala 137:31:freechips.rocketchip.system.DefaultRV32Config.fir@208384.6]
  assign _T_896 = {1'b0,$signed(_T_895)}; // @[Parameters.scala 137:49:freechips.rocketchip.system.DefaultRV32Config.fir@208385.6]
  assign _T_898 = $signed(_T_896) & -33'sh10000000; // @[Parameters.scala 137:52:freechips.rocketchip.system.DefaultRV32Config.fir@208387.6]
  assign _T_899 = $signed(_T_898) == 33'sh0; // @[Parameters.scala 137:67:freechips.rocketchip.system.DefaultRV32Config.fir@208388.6]
  assign _T_900 = io_in_b_bits_address ^ 32'h60000000; // @[Parameters.scala 137:31:freechips.rocketchip.system.DefaultRV32Config.fir@208389.6]
  assign _T_901 = {1'b0,$signed(_T_900)}; // @[Parameters.scala 137:49:freechips.rocketchip.system.DefaultRV32Config.fir@208390.6]
  assign _T_903 = $signed(_T_901) & -33'sh20000000; // @[Parameters.scala 137:52:freechips.rocketchip.system.DefaultRV32Config.fir@208392.6]
  assign _T_904 = $signed(_T_903) == 33'sh0; // @[Parameters.scala 137:67:freechips.rocketchip.system.DefaultRV32Config.fir@208393.6]
  assign _T_906 = _T_874 | _T_879; // @[Parameters.scala 535:64:freechips.rocketchip.system.DefaultRV32Config.fir@208403.6]
  assign _T_907 = _T_906 | _T_884; // @[Parameters.scala 535:64:freechips.rocketchip.system.DefaultRV32Config.fir@208404.6]
  assign _T_908 = _T_907 | _T_889; // @[Parameters.scala 535:64:freechips.rocketchip.system.DefaultRV32Config.fir@208405.6]
  assign _T_909 = _T_908 | _T_894; // @[Parameters.scala 535:64:freechips.rocketchip.system.DefaultRV32Config.fir@208406.6]
  assign _T_910 = _T_909 | _T_899; // @[Parameters.scala 535:64:freechips.rocketchip.system.DefaultRV32Config.fir@208407.6]
  assign _T_911 = _T_910 | _T_904; // @[Parameters.scala 535:64:freechips.rocketchip.system.DefaultRV32Config.fir@208408.6]
  assign _T_913 = 27'hfff << io_in_b_bits_size; // @[package.scala 207:77:freechips.rocketchip.system.DefaultRV32Config.fir@208410.6]
  assign _T_915 = ~_T_913[11:0]; // @[package.scala 207:46:freechips.rocketchip.system.DefaultRV32Config.fir@208412.6]
  assign _GEN_72 = {{20'd0}, _T_915}; // @[Edges.scala 22:16:freechips.rocketchip.system.DefaultRV32Config.fir@208413.6]
  assign _T_916 = io_in_b_bits_address & _GEN_72; // @[Edges.scala 22:16:freechips.rocketchip.system.DefaultRV32Config.fir@208413.6]
  assign _T_917 = _T_916 == 32'h0; // @[Edges.scala 22:24:freechips.rocketchip.system.DefaultRV32Config.fir@208414.6]
  assign _T_920 = 2'h1 << io_in_b_bits_size[0]; // @[OneHot.scala 65:12:freechips.rocketchip.system.DefaultRV32Config.fir@208417.6]
  assign _T_922 = _T_920 | 2'h1; // @[Misc.scala 201:81:freechips.rocketchip.system.DefaultRV32Config.fir@208419.6]
  assign _T_923 = io_in_b_bits_size >= 4'h2; // @[Misc.scala 205:21:freechips.rocketchip.system.DefaultRV32Config.fir@208420.6]
  assign _T_926 = ~io_in_b_bits_address[1]; // @[Misc.scala 210:20:freechips.rocketchip.system.DefaultRV32Config.fir@208423.6]
  assign _T_928 = _T_922[1] & _T_926; // @[Misc.scala 214:38:freechips.rocketchip.system.DefaultRV32Config.fir@208425.6]
  assign _T_929 = _T_923 | _T_928; // @[Misc.scala 214:29:freechips.rocketchip.system.DefaultRV32Config.fir@208426.6]
  assign _T_931 = _T_922[1] & io_in_b_bits_address[1]; // @[Misc.scala 214:38:freechips.rocketchip.system.DefaultRV32Config.fir@208428.6]
  assign _T_932 = _T_923 | _T_931; // @[Misc.scala 214:29:freechips.rocketchip.system.DefaultRV32Config.fir@208429.6]
  assign _T_935 = ~io_in_b_bits_address[0]; // @[Misc.scala 210:20:freechips.rocketchip.system.DefaultRV32Config.fir@208432.6]
  assign _T_936 = _T_926 & _T_935; // @[Misc.scala 213:27:freechips.rocketchip.system.DefaultRV32Config.fir@208433.6]
  assign _T_937 = _T_922[0] & _T_936; // @[Misc.scala 214:38:freechips.rocketchip.system.DefaultRV32Config.fir@208434.6]
  assign _T_938 = _T_929 | _T_937; // @[Misc.scala 214:29:freechips.rocketchip.system.DefaultRV32Config.fir@208435.6]
  assign _T_939 = _T_926 & io_in_b_bits_address[0]; // @[Misc.scala 213:27:freechips.rocketchip.system.DefaultRV32Config.fir@208436.6]
  assign _T_940 = _T_922[0] & _T_939; // @[Misc.scala 214:38:freechips.rocketchip.system.DefaultRV32Config.fir@208437.6]
  assign _T_941 = _T_929 | _T_940; // @[Misc.scala 214:29:freechips.rocketchip.system.DefaultRV32Config.fir@208438.6]
  assign _T_942 = io_in_b_bits_address[1] & _T_935; // @[Misc.scala 213:27:freechips.rocketchip.system.DefaultRV32Config.fir@208439.6]
  assign _T_943 = _T_922[0] & _T_942; // @[Misc.scala 214:38:freechips.rocketchip.system.DefaultRV32Config.fir@208440.6]
  assign _T_944 = _T_932 | _T_943; // @[Misc.scala 214:29:freechips.rocketchip.system.DefaultRV32Config.fir@208441.6]
  assign _T_945 = io_in_b_bits_address[1] & io_in_b_bits_address[0]; // @[Misc.scala 213:27:freechips.rocketchip.system.DefaultRV32Config.fir@208442.6]
  assign _T_946 = _T_922[0] & _T_945; // @[Misc.scala 214:38:freechips.rocketchip.system.DefaultRV32Config.fir@208443.6]
  assign _T_947 = _T_932 | _T_946; // @[Misc.scala 214:29:freechips.rocketchip.system.DefaultRV32Config.fir@208444.6]
  assign _T_950 = {_T_947,_T_944,_T_941,_T_938}; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@208447.6]
  assign _T_957 = _T_857 ? 2'h2 : 2'h0; // @[Mux.scala 27:72:freechips.rocketchip.system.DefaultRV32Config.fir@208458.6]
  assign _GEN_73 = {{1'd0}, _T_849}; // @[Mux.scala 27:72:freechips.rocketchip.system.DefaultRV32Config.fir@208460.6]
  assign _T_959 = _GEN_73 | _T_957; // @[Mux.scala 27:72:freechips.rocketchip.system.DefaultRV32Config.fir@208460.6]
  assign _T_961 = _T_959 == io_in_b_bits_source; // @[Monitor.scala 162:113:freechips.rocketchip.system.DefaultRV32Config.fir@208463.6]
  assign _T_962 = io_in_b_bits_opcode == 3'h6; // @[Monitor.scala 164:25:freechips.rocketchip.system.DefaultRV32Config.fir@208464.6]
  assign _T_967 = 4'h6 == io_in_b_bits_size; // @[Parameters.scala 92:48:freechips.rocketchip.system.DefaultRV32Config.fir@208474.8]
  assign _T_968 = _T_841 & _T_967; // @[Mux.scala 27:72:freechips.rocketchip.system.DefaultRV32Config.fir@208475.8]
  assign _T_975 = _T_968 | reset; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@208483.8]
  assign _T_976 = ~_T_975; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@208484.8]
  assign _T_978 = _T_911 | reset; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@208490.8]
  assign _T_979 = ~_T_978; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@208491.8]
  assign _T_981 = _T_961 | reset; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@208497.8]
  assign _T_982 = ~_T_981; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@208498.8]
  assign _T_984 = _T_917 | reset; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@208504.8]
  assign _T_985 = ~_T_984; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@208505.8]
  assign _T_986 = io_in_b_bits_param <= 2'h2; // @[Bundles.scala 104:26:freechips.rocketchip.system.DefaultRV32Config.fir@208510.8]
  assign _T_988 = _T_986 | reset; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@208512.8]
  assign _T_989 = ~_T_988; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@208513.8]
  assign _T_990 = io_in_b_bits_mask == _T_950; // @[Monitor.scala 170:30:freechips.rocketchip.system.DefaultRV32Config.fir@208518.8]
  assign _T_992 = _T_990 | reset; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@208520.8]
  assign _T_993 = ~_T_992; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@208521.8]
  assign _T_994 = ~io_in_b_bits_corrupt; // @[Monitor.scala 171:18:freechips.rocketchip.system.DefaultRV32Config.fir@208526.8]
  assign _T_996 = _T_994 | reset; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@208528.8]
  assign _T_997 = ~_T_996; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@208529.8]
  assign _T_998 = io_in_b_bits_opcode == 3'h4; // @[Monitor.scala 174:25:freechips.rocketchip.system.DefaultRV32Config.fir@208535.6]
  assign _T_1001 = ~reset; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@208539.8]
  assign _T_1011 = io_in_b_bits_param == 2'h0; // @[Monitor.scala 179:31:freechips.rocketchip.system.DefaultRV32Config.fir@208565.8]
  assign _T_1013 = _T_1011 | reset; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@208567.8]
  assign _T_1014 = ~_T_1013; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@208568.8]
  assign _T_1023 = io_in_b_bits_opcode == 3'h0; // @[Monitor.scala 184:25:freechips.rocketchip.system.DefaultRV32Config.fir@208590.6]
  assign _T_1044 = io_in_b_bits_opcode == 3'h1; // @[Monitor.scala 193:25:freechips.rocketchip.system.DefaultRV32Config.fir@208637.6]
  assign _T_1061 = ~_T_950; // @[Monitor.scala 199:33:freechips.rocketchip.system.DefaultRV32Config.fir@208675.8]
  assign _T_1062 = io_in_b_bits_mask & _T_1061; // @[Monitor.scala 199:31:freechips.rocketchip.system.DefaultRV32Config.fir@208676.8]
  assign _T_1063 = _T_1062 == 4'h0; // @[Monitor.scala 199:40:freechips.rocketchip.system.DefaultRV32Config.fir@208677.8]
  assign _T_1065 = _T_1063 | reset; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@208679.8]
  assign _T_1066 = ~_T_1065; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@208680.8]
  assign _T_1067 = io_in_b_bits_opcode == 3'h2; // @[Monitor.scala 202:25:freechips.rocketchip.system.DefaultRV32Config.fir@208686.6]
  assign _T_1088 = io_in_b_bits_opcode == 3'h3; // @[Monitor.scala 211:25:freechips.rocketchip.system.DefaultRV32Config.fir@208733.6]
  assign _T_1109 = io_in_b_bits_opcode == 3'h5; // @[Monitor.scala 220:25:freechips.rocketchip.system.DefaultRV32Config.fir@208780.6]
  assign _T_1134 = io_in_c_bits_source == 2'h0; // @[Parameters.scala 47:9:freechips.rocketchip.system.DefaultRV32Config.fir@208837.6]
  assign _T_1135 = io_in_c_bits_source == 2'h1; // @[Parameters.scala 47:9:freechips.rocketchip.system.DefaultRV32Config.fir@208838.6]
  assign _T_1136 = io_in_c_bits_source == 2'h2; // @[Parameters.scala 47:9:freechips.rocketchip.system.DefaultRV32Config.fir@208839.6]
  assign _T_1138 = _T_1134 | _T_1135; // @[Parameters.scala 924:46:freechips.rocketchip.system.DefaultRV32Config.fir@208845.6]
  assign _T_1139 = _T_1138 | _T_1136; // @[Parameters.scala 924:46:freechips.rocketchip.system.DefaultRV32Config.fir@208846.6]
  assign _T_1141 = 27'hfff << io_in_c_bits_size; // @[package.scala 207:77:freechips.rocketchip.system.DefaultRV32Config.fir@208848.6]
  assign _T_1143 = ~_T_1141[11:0]; // @[package.scala 207:46:freechips.rocketchip.system.DefaultRV32Config.fir@208850.6]
  assign _GEN_74 = {{20'd0}, _T_1143}; // @[Edges.scala 22:16:freechips.rocketchip.system.DefaultRV32Config.fir@208851.6]
  assign _T_1144 = io_in_c_bits_address & _GEN_74; // @[Edges.scala 22:16:freechips.rocketchip.system.DefaultRV32Config.fir@208851.6]
  assign _T_1145 = _T_1144 == 32'h0; // @[Edges.scala 22:24:freechips.rocketchip.system.DefaultRV32Config.fir@208852.6]
  assign _T_1146 = io_in_c_bits_address ^ 32'h3000; // @[Parameters.scala 137:31:freechips.rocketchip.system.DefaultRV32Config.fir@208853.6]
  assign _T_1147 = {1'b0,$signed(_T_1146)}; // @[Parameters.scala 137:49:freechips.rocketchip.system.DefaultRV32Config.fir@208854.6]
  assign _T_1149 = $signed(_T_1147) & -33'sh1000; // @[Parameters.scala 137:52:freechips.rocketchip.system.DefaultRV32Config.fir@208856.6]
  assign _T_1150 = $signed(_T_1149) == 33'sh0; // @[Parameters.scala 137:67:freechips.rocketchip.system.DefaultRV32Config.fir@208857.6]
  assign _T_1151 = io_in_c_bits_address ^ 32'hc000000; // @[Parameters.scala 137:31:freechips.rocketchip.system.DefaultRV32Config.fir@208858.6]
  assign _T_1152 = {1'b0,$signed(_T_1151)}; // @[Parameters.scala 137:49:freechips.rocketchip.system.DefaultRV32Config.fir@208859.6]
  assign _T_1154 = $signed(_T_1152) & -33'sh4000000; // @[Parameters.scala 137:52:freechips.rocketchip.system.DefaultRV32Config.fir@208861.6]
  assign _T_1155 = $signed(_T_1154) == 33'sh0; // @[Parameters.scala 137:67:freechips.rocketchip.system.DefaultRV32Config.fir@208862.6]
  assign _T_1156 = io_in_c_bits_address ^ 32'h2000000; // @[Parameters.scala 137:31:freechips.rocketchip.system.DefaultRV32Config.fir@208863.6]
  assign _T_1157 = {1'b0,$signed(_T_1156)}; // @[Parameters.scala 137:49:freechips.rocketchip.system.DefaultRV32Config.fir@208864.6]
  assign _T_1159 = $signed(_T_1157) & -33'sh10000; // @[Parameters.scala 137:52:freechips.rocketchip.system.DefaultRV32Config.fir@208866.6]
  assign _T_1160 = $signed(_T_1159) == 33'sh0; // @[Parameters.scala 137:67:freechips.rocketchip.system.DefaultRV32Config.fir@208867.6]
  assign _T_1162 = {1'b0,$signed(io_in_c_bits_address)}; // @[Parameters.scala 137:49:freechips.rocketchip.system.DefaultRV32Config.fir@208869.6]
  assign _T_1164 = $signed(_T_1162) & -33'sh1000; // @[Parameters.scala 137:52:freechips.rocketchip.system.DefaultRV32Config.fir@208871.6]
  assign _T_1165 = $signed(_T_1164) == 33'sh0; // @[Parameters.scala 137:67:freechips.rocketchip.system.DefaultRV32Config.fir@208872.6]
  assign _T_1166 = io_in_c_bits_address ^ 32'h10000; // @[Parameters.scala 137:31:freechips.rocketchip.system.DefaultRV32Config.fir@208873.6]
  assign _T_1167 = {1'b0,$signed(_T_1166)}; // @[Parameters.scala 137:49:freechips.rocketchip.system.DefaultRV32Config.fir@208874.6]
  assign _T_1169 = $signed(_T_1167) & -33'sh10000; // @[Parameters.scala 137:52:freechips.rocketchip.system.DefaultRV32Config.fir@208876.6]
  assign _T_1170 = $signed(_T_1169) == 33'sh0; // @[Parameters.scala 137:67:freechips.rocketchip.system.DefaultRV32Config.fir@208877.6]
  assign _T_1171 = io_in_c_bits_address ^ 32'h80000000; // @[Parameters.scala 137:31:freechips.rocketchip.system.DefaultRV32Config.fir@208878.6]
  assign _T_1172 = {1'b0,$signed(_T_1171)}; // @[Parameters.scala 137:49:freechips.rocketchip.system.DefaultRV32Config.fir@208879.6]
  assign _T_1174 = $signed(_T_1172) & -33'sh10000000; // @[Parameters.scala 137:52:freechips.rocketchip.system.DefaultRV32Config.fir@208881.6]
  assign _T_1175 = $signed(_T_1174) == 33'sh0; // @[Parameters.scala 137:67:freechips.rocketchip.system.DefaultRV32Config.fir@208882.6]
  assign _T_1176 = io_in_c_bits_address ^ 32'h60000000; // @[Parameters.scala 137:31:freechips.rocketchip.system.DefaultRV32Config.fir@208883.6]
  assign _T_1177 = {1'b0,$signed(_T_1176)}; // @[Parameters.scala 137:49:freechips.rocketchip.system.DefaultRV32Config.fir@208884.6]
  assign _T_1179 = $signed(_T_1177) & -33'sh20000000; // @[Parameters.scala 137:52:freechips.rocketchip.system.DefaultRV32Config.fir@208886.6]
  assign _T_1180 = $signed(_T_1179) == 33'sh0; // @[Parameters.scala 137:67:freechips.rocketchip.system.DefaultRV32Config.fir@208887.6]
  assign _T_1182 = _T_1150 | _T_1155; // @[Parameters.scala 535:64:freechips.rocketchip.system.DefaultRV32Config.fir@208897.6]
  assign _T_1183 = _T_1182 | _T_1160; // @[Parameters.scala 535:64:freechips.rocketchip.system.DefaultRV32Config.fir@208898.6]
  assign _T_1184 = _T_1183 | _T_1165; // @[Parameters.scala 535:64:freechips.rocketchip.system.DefaultRV32Config.fir@208899.6]
  assign _T_1185 = _T_1184 | _T_1170; // @[Parameters.scala 535:64:freechips.rocketchip.system.DefaultRV32Config.fir@208900.6]
  assign _T_1186 = _T_1185 | _T_1175; // @[Parameters.scala 535:64:freechips.rocketchip.system.DefaultRV32Config.fir@208901.6]
  assign _T_1187 = _T_1186 | _T_1180; // @[Parameters.scala 535:64:freechips.rocketchip.system.DefaultRV32Config.fir@208902.6]
  assign _T_1217 = io_in_c_bits_opcode == 3'h4; // @[Monitor.scala 239:25:freechips.rocketchip.system.DefaultRV32Config.fir@208936.6]
  assign _T_1219 = _T_1187 | reset; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@208939.8]
  assign _T_1220 = ~_T_1219; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@208940.8]
  assign _T_1222 = _T_1139 | reset; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@208946.8]
  assign _T_1223 = ~_T_1222; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@208947.8]
  assign _T_1224 = io_in_c_bits_size >= 4'h2; // @[Monitor.scala 242:30:freechips.rocketchip.system.DefaultRV32Config.fir@208952.8]
  assign _T_1226 = _T_1224 | reset; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@208954.8]
  assign _T_1227 = ~_T_1226; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@208955.8]
  assign _T_1229 = _T_1145 | reset; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@208961.8]
  assign _T_1230 = ~_T_1229; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@208962.8]
  assign _T_1231 = io_in_c_bits_param <= 3'h5; // @[Bundles.scala 122:29:freechips.rocketchip.system.DefaultRV32Config.fir@208967.8]
  assign _T_1233 = _T_1231 | reset; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@208969.8]
  assign _T_1234 = ~_T_1233; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@208970.8]
  assign _T_1239 = io_in_c_bits_opcode == 3'h5; // @[Monitor.scala 248:25:freechips.rocketchip.system.DefaultRV32Config.fir@208984.6]
  assign _T_1257 = io_in_c_bits_opcode == 3'h6; // @[Monitor.scala 256:25:freechips.rocketchip.system.DefaultRV32Config.fir@209024.6]
  assign _T_1296 = io_in_c_bits_size <= 4'h6; // @[Parameters.scala 93:42:freechips.rocketchip.system.DefaultRV32Config.fir@209064.8]
  assign _T_1304 = _T_1296 & _T_1175; // @[Parameters.scala 551:56:freechips.rocketchip.system.DefaultRV32Config.fir@209072.8]
  assign _T_1308 = _T_1304 | reset; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@209076.8]
  assign _T_1309 = ~_T_1308; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@209077.8]
  assign _T_1314 = 4'h6 == io_in_c_bits_size; // @[Parameters.scala 92:48:freechips.rocketchip.system.DefaultRV32Config.fir@209090.8]
  assign _T_1315 = _T_1134 & _T_1314; // @[Mux.scala 27:72:freechips.rocketchip.system.DefaultRV32Config.fir@209091.8]
  assign _T_1322 = _T_1315 | reset; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@209099.8]
  assign _T_1323 = ~_T_1322; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@209100.8]
  assign _T_1334 = io_in_c_bits_param <= 3'h2; // @[Bundles.scala 116:29:freechips.rocketchip.system.DefaultRV32Config.fir@209127.8]
  assign _T_1336 = _T_1334 | reset; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@209129.8]
  assign _T_1337 = ~_T_1336; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@209130.8]
  assign _T_1342 = io_in_c_bits_opcode == 3'h7; // @[Monitor.scala 266:25:freechips.rocketchip.system.DefaultRV32Config.fir@209144.6]
  assign _T_1423 = io_in_c_bits_opcode == 3'h0; // @[Monitor.scala 275:25:freechips.rocketchip.system.DefaultRV32Config.fir@209256.6]
  assign _T_1433 = io_in_c_bits_param == 3'h0; // @[Monitor.scala 279:31:freechips.rocketchip.system.DefaultRV32Config.fir@209279.8]
  assign _T_1435 = _T_1433 | reset; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@209281.8]
  assign _T_1436 = ~_T_1435; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@209282.8]
  assign _T_1441 = io_in_c_bits_opcode == 3'h1; // @[Monitor.scala 283:25:freechips.rocketchip.system.DefaultRV32Config.fir@209296.6]
  assign _T_1455 = io_in_c_bits_opcode == 3'h2; // @[Monitor.scala 290:25:freechips.rocketchip.system.DefaultRV32Config.fir@209328.6]
  assign _T_1477 = io_in_a_ready & io_in_a_valid; // @[Decoupled.scala 40:37:freechips.rocketchip.system.DefaultRV32Config.fir@209379.4]
  assign _T_1484 = ~io_in_a_bits_opcode[2]; // @[Edges.scala 93:28:freechips.rocketchip.system.DefaultRV32Config.fir@209386.4]
  assign _T_1488 = _T_1486 - 10'h1; // @[Edges.scala 231:28:freechips.rocketchip.system.DefaultRV32Config.fir@209390.4]
  assign _T_1489 = _T_1486 == 10'h0; // @[Edges.scala 232:25:freechips.rocketchip.system.DefaultRV32Config.fir@209391.4]
  assign _T_1502 = ~_T_1489; // @[Monitor.scala 386:22:freechips.rocketchip.system.DefaultRV32Config.fir@209407.4]
  assign _T_1503 = io_in_a_valid & _T_1502; // @[Monitor.scala 386:19:freechips.rocketchip.system.DefaultRV32Config.fir@209408.4]
  assign _T_1504 = io_in_a_bits_opcode == _T_1497; // @[Monitor.scala 387:32:freechips.rocketchip.system.DefaultRV32Config.fir@209410.6]
  assign _T_1506 = _T_1504 | reset; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@209412.6]
  assign _T_1507 = ~_T_1506; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@209413.6]
  assign _T_1508 = io_in_a_bits_param == _T_1498; // @[Monitor.scala 388:32:freechips.rocketchip.system.DefaultRV32Config.fir@209418.6]
  assign _T_1510 = _T_1508 | reset; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@209420.6]
  assign _T_1511 = ~_T_1510; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@209421.6]
  assign _T_1512 = io_in_a_bits_size == _T_1499; // @[Monitor.scala 389:32:freechips.rocketchip.system.DefaultRV32Config.fir@209426.6]
  assign _T_1514 = _T_1512 | reset; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@209428.6]
  assign _T_1515 = ~_T_1514; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@209429.6]
  assign _T_1516 = io_in_a_bits_source == _T_1500; // @[Monitor.scala 390:32:freechips.rocketchip.system.DefaultRV32Config.fir@209434.6]
  assign _T_1518 = _T_1516 | reset; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@209436.6]
  assign _T_1519 = ~_T_1518; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@209437.6]
  assign _T_1520 = io_in_a_bits_address == _T_1501; // @[Monitor.scala 391:32:freechips.rocketchip.system.DefaultRV32Config.fir@209442.6]
  assign _T_1522 = _T_1520 | reset; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@209444.6]
  assign _T_1523 = ~_T_1522; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@209445.6]
  assign _T_1525 = _T_1477 & _T_1489; // @[Monitor.scala 393:20:freechips.rocketchip.system.DefaultRV32Config.fir@209452.4]
  assign _T_1526 = io_in_d_ready & io_in_d_valid; // @[Decoupled.scala 40:37:freechips.rocketchip.system.DefaultRV32Config.fir@209460.4]
  assign _T_1528 = 27'hfff << io_in_d_bits_size; // @[package.scala 207:77:freechips.rocketchip.system.DefaultRV32Config.fir@209462.4]
  assign _T_1530 = ~_T_1528[11:0]; // @[package.scala 207:46:freechips.rocketchip.system.DefaultRV32Config.fir@209464.4]
  assign _T_1536 = _T_1534 - 10'h1; // @[Edges.scala 231:28:freechips.rocketchip.system.DefaultRV32Config.fir@209470.4]
  assign _T_1537 = _T_1534 == 10'h0; // @[Edges.scala 232:25:freechips.rocketchip.system.DefaultRV32Config.fir@209471.4]
  assign _T_1551 = ~_T_1537; // @[Monitor.scala 538:22:freechips.rocketchip.system.DefaultRV32Config.fir@209488.4]
  assign _T_1552 = io_in_d_valid & _T_1551; // @[Monitor.scala 538:19:freechips.rocketchip.system.DefaultRV32Config.fir@209489.4]
  assign _T_1553 = io_in_d_bits_opcode == _T_1545; // @[Monitor.scala 539:29:freechips.rocketchip.system.DefaultRV32Config.fir@209491.6]
  assign _T_1555 = _T_1553 | reset; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@209493.6]
  assign _T_1556 = ~_T_1555; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@209494.6]
  assign _T_1557 = io_in_d_bits_param == _T_1546; // @[Monitor.scala 540:29:freechips.rocketchip.system.DefaultRV32Config.fir@209499.6]
  assign _T_1559 = _T_1557 | reset; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@209501.6]
  assign _T_1560 = ~_T_1559; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@209502.6]
  assign _T_1561 = io_in_d_bits_size == _T_1547; // @[Monitor.scala 541:29:freechips.rocketchip.system.DefaultRV32Config.fir@209507.6]
  assign _T_1563 = _T_1561 | reset; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@209509.6]
  assign _T_1564 = ~_T_1563; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@209510.6]
  assign _T_1565 = io_in_d_bits_source == _T_1548; // @[Monitor.scala 542:29:freechips.rocketchip.system.DefaultRV32Config.fir@209515.6]
  assign _T_1567 = _T_1565 | reset; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@209517.6]
  assign _T_1568 = ~_T_1567; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@209518.6]
  assign _T_1569 = io_in_d_bits_sink == _T_1549; // @[Monitor.scala 543:29:freechips.rocketchip.system.DefaultRV32Config.fir@209523.6]
  assign _T_1571 = _T_1569 | reset; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@209525.6]
  assign _T_1572 = ~_T_1571; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@209526.6]
  assign _T_1573 = io_in_d_bits_denied == _T_1550; // @[Monitor.scala 544:29:freechips.rocketchip.system.DefaultRV32Config.fir@209531.6]
  assign _T_1575 = _T_1573 | reset; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@209533.6]
  assign _T_1576 = ~_T_1575; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@209534.6]
  assign _T_1578 = _T_1526 & _T_1537; // @[Monitor.scala 546:20:freechips.rocketchip.system.DefaultRV32Config.fir@209541.4]
  assign _T_1579 = io_in_b_ready & io_in_b_valid; // @[Decoupled.scala 40:37:freechips.rocketchip.system.DefaultRV32Config.fir@209550.4]
  assign _T_1590 = _T_1588 - 10'h1; // @[Edges.scala 231:28:freechips.rocketchip.system.DefaultRV32Config.fir@209561.4]
  assign _T_1591 = _T_1588 == 10'h0; // @[Edges.scala 232:25:freechips.rocketchip.system.DefaultRV32Config.fir@209562.4]
  assign _T_1604 = ~_T_1591; // @[Monitor.scala 409:22:freechips.rocketchip.system.DefaultRV32Config.fir@209578.4]
  assign _T_1605 = io_in_b_valid & _T_1604; // @[Monitor.scala 409:19:freechips.rocketchip.system.DefaultRV32Config.fir@209579.4]
  assign _T_1606 = io_in_b_bits_opcode == _T_1599; // @[Monitor.scala 410:32:freechips.rocketchip.system.DefaultRV32Config.fir@209581.6]
  assign _T_1608 = _T_1606 | reset; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@209583.6]
  assign _T_1609 = ~_T_1608; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@209584.6]
  assign _T_1610 = io_in_b_bits_param == _T_1600; // @[Monitor.scala 411:32:freechips.rocketchip.system.DefaultRV32Config.fir@209589.6]
  assign _T_1612 = _T_1610 | reset; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@209591.6]
  assign _T_1613 = ~_T_1612; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@209592.6]
  assign _T_1614 = io_in_b_bits_size == _T_1601; // @[Monitor.scala 412:32:freechips.rocketchip.system.DefaultRV32Config.fir@209597.6]
  assign _T_1616 = _T_1614 | reset; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@209599.6]
  assign _T_1617 = ~_T_1616; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@209600.6]
  assign _T_1618 = io_in_b_bits_source == _T_1602; // @[Monitor.scala 413:32:freechips.rocketchip.system.DefaultRV32Config.fir@209605.6]
  assign _T_1620 = _T_1618 | reset; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@209607.6]
  assign _T_1621 = ~_T_1620; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@209608.6]
  assign _T_1622 = io_in_b_bits_address == _T_1603; // @[Monitor.scala 414:32:freechips.rocketchip.system.DefaultRV32Config.fir@209613.6]
  assign _T_1624 = _T_1622 | reset; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@209615.6]
  assign _T_1625 = ~_T_1624; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@209616.6]
  assign _T_1627 = _T_1579 & _T_1591; // @[Monitor.scala 416:20:freechips.rocketchip.system.DefaultRV32Config.fir@209623.4]
  assign _T_1628 = io_in_c_ready & io_in_c_valid; // @[Decoupled.scala 40:37:freechips.rocketchip.system.DefaultRV32Config.fir@209631.4]
  assign _T_1638 = _T_1636 - 10'h1; // @[Edges.scala 231:28:freechips.rocketchip.system.DefaultRV32Config.fir@209641.4]
  assign _T_1639 = _T_1636 == 10'h0; // @[Edges.scala 232:25:freechips.rocketchip.system.DefaultRV32Config.fir@209642.4]
  assign _T_1652 = ~_T_1639; // @[Monitor.scala 514:22:freechips.rocketchip.system.DefaultRV32Config.fir@209658.4]
  assign _T_1653 = io_in_c_valid & _T_1652; // @[Monitor.scala 514:19:freechips.rocketchip.system.DefaultRV32Config.fir@209659.4]
  assign _T_1654 = io_in_c_bits_opcode == _T_1647; // @[Monitor.scala 515:32:freechips.rocketchip.system.DefaultRV32Config.fir@209661.6]
  assign _T_1656 = _T_1654 | reset; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@209663.6]
  assign _T_1657 = ~_T_1656; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@209664.6]
  assign _T_1658 = io_in_c_bits_param == _T_1648; // @[Monitor.scala 516:32:freechips.rocketchip.system.DefaultRV32Config.fir@209669.6]
  assign _T_1660 = _T_1658 | reset; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@209671.6]
  assign _T_1661 = ~_T_1660; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@209672.6]
  assign _T_1662 = io_in_c_bits_size == _T_1649; // @[Monitor.scala 517:32:freechips.rocketchip.system.DefaultRV32Config.fir@209677.6]
  assign _T_1664 = _T_1662 | reset; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@209679.6]
  assign _T_1665 = ~_T_1664; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@209680.6]
  assign _T_1666 = io_in_c_bits_source == _T_1650; // @[Monitor.scala 518:32:freechips.rocketchip.system.DefaultRV32Config.fir@209685.6]
  assign _T_1668 = _T_1666 | reset; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@209687.6]
  assign _T_1669 = ~_T_1668; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@209688.6]
  assign _T_1670 = io_in_c_bits_address == _T_1651; // @[Monitor.scala 519:32:freechips.rocketchip.system.DefaultRV32Config.fir@209693.6]
  assign _T_1672 = _T_1670 | reset; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@209695.6]
  assign _T_1673 = ~_T_1672; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@209696.6]
  assign _T_1675 = _T_1628 & _T_1639; // @[Monitor.scala 521:20:freechips.rocketchip.system.DefaultRV32Config.fir@209703.4]
  assign _T_1687 = _T_1685 - 10'h1; // @[Edges.scala 231:28:freechips.rocketchip.system.DefaultRV32Config.fir@209725.4]
  assign a_first = _T_1685 == 10'h0; // @[Edges.scala 232:25:freechips.rocketchip.system.DefaultRV32Config.fir@209726.4]
  assign _T_1705 = _T_1703 - 10'h1; // @[Edges.scala 231:28:freechips.rocketchip.system.DefaultRV32Config.fir@209747.4]
  assign d_first = _T_1703 == 10'h0; // @[Edges.scala 232:25:freechips.rocketchip.system.DefaultRV32Config.fir@209748.4]
  assign _GEN_75 = {io_in_d_bits_source, 2'h0}; // @[Monitor.scala 629:69:freechips.rocketchip.system.DefaultRV32Config.fir@209767.4]
  assign _T_1713 = {{1'd0}, _GEN_75}; // @[Monitor.scala 629:69:freechips.rocketchip.system.DefaultRV32Config.fir@209767.4]
  assign _T_1714 = inflight_opcodes >> _T_1713; // @[Monitor.scala 629:44:freechips.rocketchip.system.DefaultRV32Config.fir@209768.4]
  assign _T_1718 = 16'h10 - 16'h1; // @[Monitor.scala 606:57:freechips.rocketchip.system.DefaultRV32Config.fir@209772.4]
  assign _GEN_76 = {{4'd0}, _T_1714}; // @[Monitor.scala 629:97:freechips.rocketchip.system.DefaultRV32Config.fir@209773.4]
  assign _T_1719 = _GEN_76 & _T_1718; // @[Monitor.scala 629:97:freechips.rocketchip.system.DefaultRV32Config.fir@209773.4]
  assign _T_1720 = {{1'd0}, _T_1719[15:1]}; // @[Monitor.scala 629:152:freechips.rocketchip.system.DefaultRV32Config.fir@209774.4]
  assign _T_1721 = {io_in_d_bits_source, 3'h0}; // @[Monitor.scala 633:65:freechips.rocketchip.system.DefaultRV32Config.fir@209778.4]
  assign _T_1722 = inflight_sizes >> _T_1721; // @[Monitor.scala 633:40:freechips.rocketchip.system.DefaultRV32Config.fir@209779.4]
  assign _T_1726 = 16'h100 - 16'h1; // @[Monitor.scala 606:57:freechips.rocketchip.system.DefaultRV32Config.fir@209783.4]
  assign _GEN_78 = {{8'd0}, _T_1726}; // @[Monitor.scala 633:91:freechips.rocketchip.system.DefaultRV32Config.fir@209784.4]
  assign _T_1727 = _T_1722 & _GEN_78; // @[Monitor.scala 633:91:freechips.rocketchip.system.DefaultRV32Config.fir@209784.4]
  assign _T_1728 = {{1'd0}, _T_1727[23:1]}; // @[Monitor.scala 633:144:freechips.rocketchip.system.DefaultRV32Config.fir@209785.4]
  assign _T_1732 = _T_1477 & a_first; // @[Monitor.scala 643:27:freechips.rocketchip.system.DefaultRV32Config.fir@209810.4]
  assign _T_1734 = 4'h1 << io_in_a_bits_source; // @[OneHot.scala 58:35:freechips.rocketchip.system.DefaultRV32Config.fir@209813.6]
  assign _T_1735 = {io_in_a_bits_opcode, 1'h0}; // @[Monitor.scala 645:53:freechips.rocketchip.system.DefaultRV32Config.fir@209815.6]
  assign _T_1736 = _T_1735 | 4'h1; // @[Monitor.scala 645:61:freechips.rocketchip.system.DefaultRV32Config.fir@209816.6]
  assign _T_1737 = {io_in_a_bits_size, 1'h0}; // @[Monitor.scala 646:49:freechips.rocketchip.system.DefaultRV32Config.fir@209818.6]
  assign _T_1738 = _T_1737 | 5'h1; // @[Monitor.scala 646:57:freechips.rocketchip.system.DefaultRV32Config.fir@209819.6]
  assign _GEN_80 = {io_in_a_bits_source, 2'h0}; // @[Monitor.scala 647:72:freechips.rocketchip.system.DefaultRV32Config.fir@209821.6]
  assign _T_1739 = {{1'd0}, _GEN_80}; // @[Monitor.scala 647:72:freechips.rocketchip.system.DefaultRV32Config.fir@209821.6]
  assign a_opcodes_set_interm = _T_1732 ? _T_1736 : 4'h0; // @[Monitor.scala 643:72:freechips.rocketchip.system.DefaultRV32Config.fir@209812.4]
  assign _GEN_81 = {{31'd0}, a_opcodes_set_interm}; // @[Monitor.scala 647:47:freechips.rocketchip.system.DefaultRV32Config.fir@209822.6]
  assign _T_1740 = _GEN_81 << _T_1739; // @[Monitor.scala 647:47:freechips.rocketchip.system.DefaultRV32Config.fir@209822.6]
  assign _T_1741 = {io_in_a_bits_source, 3'h0}; // @[Monitor.scala 648:68:freechips.rocketchip.system.DefaultRV32Config.fir@209824.6]
  assign a_sizes_set_interm = _T_1732 ? _T_1738 : 5'h0; // @[Monitor.scala 643:72:freechips.rocketchip.system.DefaultRV32Config.fir@209812.4]
  assign _GEN_82 = {{31'd0}, a_sizes_set_interm}; // @[Monitor.scala 648:43:freechips.rocketchip.system.DefaultRV32Config.fir@209825.6]
  assign _T_1742 = _GEN_82 << _T_1741; // @[Monitor.scala 648:43:freechips.rocketchip.system.DefaultRV32Config.fir@209825.6]
  assign _T_1743 = inflight >> io_in_a_bits_source; // @[Monitor.scala 649:26:freechips.rocketchip.system.DefaultRV32Config.fir@209827.6]
  assign _T_1745 = ~_T_1743[0]; // @[Monitor.scala 649:17:freechips.rocketchip.system.DefaultRV32Config.fir@209829.6]
  assign _T_1747 = _T_1745 | reset; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@209831.6]
  assign _T_1748 = ~_T_1747; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@209832.6]
  assign _GEN_27 = _T_1732 ? _T_1734 : 4'h0; // @[Monitor.scala 643:72:freechips.rocketchip.system.DefaultRV32Config.fir@209812.4]
  assign _GEN_30 = _T_1732 ? _T_1740 : 35'h0; // @[Monitor.scala 643:72:freechips.rocketchip.system.DefaultRV32Config.fir@209812.4]
  assign _GEN_31 = _T_1732 ? _T_1742 : 36'h0; // @[Monitor.scala 643:72:freechips.rocketchip.system.DefaultRV32Config.fir@209812.4]
  assign _T_1751 = _T_1526 & d_first; // @[Monitor.scala 660:27:freechips.rocketchip.system.DefaultRV32Config.fir@209846.4]
  assign _T_1753 = ~_T_708; // @[Monitor.scala 660:75:freechips.rocketchip.system.DefaultRV32Config.fir@209848.4]
  assign _T_1754 = _T_1751 & _T_1753; // @[Monitor.scala 660:72:freechips.rocketchip.system.DefaultRV32Config.fir@209849.4]
  assign _T_1755 = 4'h1 << io_in_d_bits_source; // @[OneHot.scala 58:35:freechips.rocketchip.system.DefaultRV32Config.fir@209851.6]
  assign _GEN_84 = {{31'd0}, _T_1718}; // @[Monitor.scala 662:76:freechips.rocketchip.system.DefaultRV32Config.fir@209858.6]
  assign _T_1761 = _GEN_84 << _T_1713; // @[Monitor.scala 662:76:freechips.rocketchip.system.DefaultRV32Config.fir@209858.6]
  assign _GEN_85 = {{31'd0}, _T_1726}; // @[Monitor.scala 663:72:freechips.rocketchip.system.DefaultRV32Config.fir@209865.6]
  assign _T_1767 = _GEN_85 << _T_1721; // @[Monitor.scala 663:72:freechips.rocketchip.system.DefaultRV32Config.fir@209865.6]
  assign _GEN_32 = _T_1754 ? _T_1755 : 4'h0; // @[Monitor.scala 660:91:freechips.rocketchip.system.DefaultRV32Config.fir@209850.4]
  assign _GEN_33 = _T_1754 ? _T_1761 : 47'h0; // @[Monitor.scala 660:91:freechips.rocketchip.system.DefaultRV32Config.fir@209850.4]
  assign _GEN_34 = _T_1754 ? _T_1767 : 47'h0; // @[Monitor.scala 660:91:freechips.rocketchip.system.DefaultRV32Config.fir@209850.4]
  assign _T_1768 = io_in_d_valid & d_first; // @[Monitor.scala 665:26:freechips.rocketchip.system.DefaultRV32Config.fir@209868.4]
  assign _T_1771 = _T_1768 & _T_1753; // @[Monitor.scala 665:71:freechips.rocketchip.system.DefaultRV32Config.fir@209871.4]
  assign _T_1772 = inflight >> io_in_d_bits_source; // @[Monitor.scala 666:25:freechips.rocketchip.system.DefaultRV32Config.fir@209873.6]
  assign _T_1774 = io_in_a_bits_source == io_in_d_bits_source; // @[Monitor.scala 666:93:freechips.rocketchip.system.DefaultRV32Config.fir@209875.6]
  assign _T_1775 = io_in_a_valid & _T_1774; // @[Monitor.scala 666:68:freechips.rocketchip.system.DefaultRV32Config.fir@209876.6]
  assign _T_1776 = io_in_a_bits_size == io_in_d_bits_size; // @[Monitor.scala 666:142:freechips.rocketchip.system.DefaultRV32Config.fir@209877.6]
  assign _T_1777 = _T_1775 & _T_1776; // @[Monitor.scala 666:119:freechips.rocketchip.system.DefaultRV32Config.fir@209878.6]
  assign _T_1778 = _T_1777 & a_first; // @[Monitor.scala 666:166:freechips.rocketchip.system.DefaultRV32Config.fir@209879.6]
  assign _T_1779 = _T_1772[0] | _T_1778; // @[Monitor.scala 666:49:freechips.rocketchip.system.DefaultRV32Config.fir@209880.6]
  assign _T_1781 = _T_1779 | reset; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@209882.6]
  assign _T_1782 = ~_T_1781; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@209883.6]
  assign a_opcode_lookup = _T_1720[3:0]; // @[:freechips.rocketchip.system.DefaultRV32Config.fir@209765.4 :freechips.rocketchip.system.DefaultRV32Config.fir@209766.4 Monitor.scala 629:21:freechips.rocketchip.system.DefaultRV32Config.fir@209775.4]
  assign _GEN_37 = 3'h2 == a_opcode_lookup[2:0] ? 3'h1 : 3'h0; // @[Monitor.scala 667:37:freechips.rocketchip.system.DefaultRV32Config.fir@209889.6]
  assign _GEN_38 = 3'h3 == a_opcode_lookup[2:0] ? 3'h1 : _GEN_37; // @[Monitor.scala 667:37:freechips.rocketchip.system.DefaultRV32Config.fir@209889.6]
  assign _GEN_39 = 3'h4 == a_opcode_lookup[2:0] ? 3'h1 : _GEN_38; // @[Monitor.scala 667:37:freechips.rocketchip.system.DefaultRV32Config.fir@209889.6]
  assign _GEN_40 = 3'h5 == a_opcode_lookup[2:0] ? 3'h2 : _GEN_39; // @[Monitor.scala 667:37:freechips.rocketchip.system.DefaultRV32Config.fir@209889.6]
  assign _GEN_41 = 3'h6 == a_opcode_lookup[2:0] ? 3'h4 : _GEN_40; // @[Monitor.scala 667:37:freechips.rocketchip.system.DefaultRV32Config.fir@209889.6]
  assign _GEN_42 = 3'h7 == a_opcode_lookup[2:0] ? 3'h4 : _GEN_41; // @[Monitor.scala 667:37:freechips.rocketchip.system.DefaultRV32Config.fir@209889.6]
  assign _T_1784 = io_in_d_bits_opcode == _GEN_42; // @[Monitor.scala 667:37:freechips.rocketchip.system.DefaultRV32Config.fir@209889.6]
  assign _GEN_49 = 3'h6 == a_opcode_lookup[2:0] ? 3'h5 : _GEN_40; // @[Monitor.scala 667:96:freechips.rocketchip.system.DefaultRV32Config.fir@209891.6]
  assign _GEN_50 = 3'h7 == a_opcode_lookup[2:0] ? 3'h4 : _GEN_49; // @[Monitor.scala 667:96:freechips.rocketchip.system.DefaultRV32Config.fir@209891.6]
  assign _T_1786 = io_in_d_bits_opcode == _GEN_50; // @[Monitor.scala 667:96:freechips.rocketchip.system.DefaultRV32Config.fir@209891.6]
  assign _T_1787 = _T_1784 | _T_1786; // @[Monitor.scala 667:71:freechips.rocketchip.system.DefaultRV32Config.fir@209892.6]
  assign _GEN_53 = 3'h2 == io_in_a_bits_opcode ? 3'h1 : 3'h0; // @[Monitor.scala 668:60:freechips.rocketchip.system.DefaultRV32Config.fir@209893.6]
  assign _GEN_54 = 3'h3 == io_in_a_bits_opcode ? 3'h1 : _GEN_53; // @[Monitor.scala 668:60:freechips.rocketchip.system.DefaultRV32Config.fir@209893.6]
  assign _GEN_55 = 3'h4 == io_in_a_bits_opcode ? 3'h1 : _GEN_54; // @[Monitor.scala 668:60:freechips.rocketchip.system.DefaultRV32Config.fir@209893.6]
  assign _GEN_56 = 3'h5 == io_in_a_bits_opcode ? 3'h2 : _GEN_55; // @[Monitor.scala 668:60:freechips.rocketchip.system.DefaultRV32Config.fir@209893.6]
  assign _GEN_57 = 3'h6 == io_in_a_bits_opcode ? 3'h4 : _GEN_56; // @[Monitor.scala 668:60:freechips.rocketchip.system.DefaultRV32Config.fir@209893.6]
  assign _GEN_58 = 3'h7 == io_in_a_bits_opcode ? 3'h4 : _GEN_57; // @[Monitor.scala 668:60:freechips.rocketchip.system.DefaultRV32Config.fir@209893.6]
  assign _T_1788 = io_in_d_bits_opcode == _GEN_58; // @[Monitor.scala 668:60:freechips.rocketchip.system.DefaultRV32Config.fir@209893.6]
  assign _GEN_65 = 3'h6 == io_in_a_bits_opcode ? 3'h5 : _GEN_56; // @[Monitor.scala 668:124:freechips.rocketchip.system.DefaultRV32Config.fir@209894.6]
  assign _GEN_66 = 3'h7 == io_in_a_bits_opcode ? 3'h4 : _GEN_65; // @[Monitor.scala 668:124:freechips.rocketchip.system.DefaultRV32Config.fir@209894.6]
  assign _T_1789 = io_in_d_bits_opcode == _GEN_66; // @[Monitor.scala 668:124:freechips.rocketchip.system.DefaultRV32Config.fir@209894.6]
  assign _T_1790 = _T_1788 | _T_1789; // @[Monitor.scala 668:99:freechips.rocketchip.system.DefaultRV32Config.fir@209895.6]
  assign _T_1791 = io_in_a_valid & _T_1790; // @[Monitor.scala 668:34:freechips.rocketchip.system.DefaultRV32Config.fir@209896.6]
  assign _T_1792 = _T_1787 | _T_1791; // @[Monitor.scala 668:15:freechips.rocketchip.system.DefaultRV32Config.fir@209897.6]
  assign _T_1794 = _T_1792 | reset; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@209899.6]
  assign _T_1795 = ~_T_1794; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@209900.6]
  assign a_size_lookup = _T_1728[7:0]; // @[:freechips.rocketchip.system.DefaultRV32Config.fir@209776.4 :freechips.rocketchip.system.DefaultRV32Config.fir@209777.4 Monitor.scala 633:19:freechips.rocketchip.system.DefaultRV32Config.fir@209786.4]
  assign _GEN_86 = {{4'd0}, io_in_d_bits_size}; // @[Monitor.scala 670:34:freechips.rocketchip.system.DefaultRV32Config.fir@209905.6]
  assign _T_1796 = _GEN_86 == a_size_lookup; // @[Monitor.scala 670:34:freechips.rocketchip.system.DefaultRV32Config.fir@209905.6]
  assign _T_1798 = io_in_a_valid & _T_1776; // @[Monitor.scala 670:72:freechips.rocketchip.system.DefaultRV32Config.fir@209907.6]
  assign _T_1799 = _T_1796 | _T_1798; // @[Monitor.scala 670:53:freechips.rocketchip.system.DefaultRV32Config.fir@209908.6]
  assign _T_1801 = _T_1799 | reset; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@209910.6]
  assign _T_1802 = ~_T_1801; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@209911.6]
  assign _T_1804 = _T_1768 & a_first; // @[Monitor.scala 672:36:freechips.rocketchip.system.DefaultRV32Config.fir@209918.4]
  assign _T_1805 = _T_1804 & io_in_a_valid; // @[Monitor.scala 672:47:freechips.rocketchip.system.DefaultRV32Config.fir@209919.4]
  assign _T_1807 = _T_1805 & _T_1774; // @[Monitor.scala 672:65:freechips.rocketchip.system.DefaultRV32Config.fir@209921.4]
  assign _T_1809 = _T_1807 & _T_1753; // @[Monitor.scala 672:116:freechips.rocketchip.system.DefaultRV32Config.fir@209923.4]
  assign _T_1810 = ~io_in_d_ready; // @[Monitor.scala 673:15:freechips.rocketchip.system.DefaultRV32Config.fir@209925.6]
  assign _T_1811 = _T_1810 | io_in_a_ready; // @[Monitor.scala 673:32:freechips.rocketchip.system.DefaultRV32Config.fir@209926.6]
  assign _T_1813 = _T_1811 | reset; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@209928.6]
  assign _T_1814 = ~_T_1813; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@209929.6]
  assign a_set = _GEN_27[2:0]; // @[:freechips.rocketchip.system.DefaultRV32Config.fir@209759.4 :freechips.rocketchip.system.DefaultRV32Config.fir@209760.4 Monitor.scala 644:13:freechips.rocketchip.system.DefaultRV32Config.fir@209814.6]
  assign d_clr = _GEN_32[2:0]; // @[:freechips.rocketchip.system.DefaultRV32Config.fir@209838.4 :freechips.rocketchip.system.DefaultRV32Config.fir@209839.4 Monitor.scala 661:13:freechips.rocketchip.system.DefaultRV32Config.fir@209852.6]
  assign _T_1815 = a_set != d_clr; // @[Monitor.scala 677:20:freechips.rocketchip.system.DefaultRV32Config.fir@209935.4]
  assign _T_1816 = |a_set; // @[Monitor.scala 677:40:freechips.rocketchip.system.DefaultRV32Config.fir@209936.4]
  assign _T_1817 = ~_T_1816; // @[Monitor.scala 677:33:freechips.rocketchip.system.DefaultRV32Config.fir@209937.4]
  assign _T_1818 = _T_1815 | _T_1817; // @[Monitor.scala 677:30:freechips.rocketchip.system.DefaultRV32Config.fir@209938.4]
  assign _T_1820 = _T_1818 | reset; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@209940.4]
  assign _T_1821 = ~_T_1820; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@209941.4]
  assign _T_1822 = inflight | a_set; // @[Monitor.scala 680:27:freechips.rocketchip.system.DefaultRV32Config.fir@209946.4]
  assign _T_1823 = ~d_clr; // @[Monitor.scala 680:38:freechips.rocketchip.system.DefaultRV32Config.fir@209947.4]
  assign _T_1824 = _T_1822 & _T_1823; // @[Monitor.scala 680:36:freechips.rocketchip.system.DefaultRV32Config.fir@209948.4]
  assign a_opcodes_set = _GEN_30[11:0]; // @[:freechips.rocketchip.system.DefaultRV32Config.fir@209761.4 :freechips.rocketchip.system.DefaultRV32Config.fir@209762.4 Monitor.scala 647:21:freechips.rocketchip.system.DefaultRV32Config.fir@209823.6]
  assign _T_1825 = inflight_opcodes | a_opcodes_set; // @[Monitor.scala 681:43:freechips.rocketchip.system.DefaultRV32Config.fir@209950.4]
  assign d_opcodes_clr = _GEN_33[11:0]; // @[:freechips.rocketchip.system.DefaultRV32Config.fir@209840.4 :freechips.rocketchip.system.DefaultRV32Config.fir@209841.4 Monitor.scala 662:21:freechips.rocketchip.system.DefaultRV32Config.fir@209859.6]
  assign _T_1826 = ~d_opcodes_clr; // @[Monitor.scala 681:62:freechips.rocketchip.system.DefaultRV32Config.fir@209951.4]
  assign _T_1827 = _T_1825 & _T_1826; // @[Monitor.scala 681:60:freechips.rocketchip.system.DefaultRV32Config.fir@209952.4]
  assign a_sizes_set = _GEN_31[23:0]; // @[:freechips.rocketchip.system.DefaultRV32Config.fir@209763.4 :freechips.rocketchip.system.DefaultRV32Config.fir@209764.4 Monitor.scala 648:19:freechips.rocketchip.system.DefaultRV32Config.fir@209826.6]
  assign _T_1828 = inflight_sizes | a_sizes_set; // @[Monitor.scala 682:39:freechips.rocketchip.system.DefaultRV32Config.fir@209954.4]
  assign d_sizes_clr = _GEN_34[23:0]; // @[:freechips.rocketchip.system.DefaultRV32Config.fir@209842.4 :freechips.rocketchip.system.DefaultRV32Config.fir@209843.4 Monitor.scala 663:19:freechips.rocketchip.system.DefaultRV32Config.fir@209866.6]
  assign _T_1829 = ~d_sizes_clr; // @[Monitor.scala 682:56:freechips.rocketchip.system.DefaultRV32Config.fir@209955.4]
  assign _T_1830 = _T_1828 & _T_1829; // @[Monitor.scala 682:54:freechips.rocketchip.system.DefaultRV32Config.fir@209956.4]
  assign _T_1832 = |inflight; // @[Monitor.scala 687:26:freechips.rocketchip.system.DefaultRV32Config.fir@209961.4]
  assign _T_1833 = ~_T_1832; // @[Monitor.scala 687:16:freechips.rocketchip.system.DefaultRV32Config.fir@209962.4]
  assign _T_1834 = plusarg_reader_out == 32'h0; // @[Monitor.scala 687:39:freechips.rocketchip.system.DefaultRV32Config.fir@209963.4]
  assign _T_1835 = _T_1833 | _T_1834; // @[Monitor.scala 687:30:freechips.rocketchip.system.DefaultRV32Config.fir@209964.4]
  assign _T_1836 = _T_1831 < plusarg_reader_out; // @[Monitor.scala 687:59:freechips.rocketchip.system.DefaultRV32Config.fir@209965.4]
  assign _T_1837 = _T_1835 | _T_1836; // @[Monitor.scala 687:47:freechips.rocketchip.system.DefaultRV32Config.fir@209966.4]
  assign _T_1839 = _T_1837 | reset; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@209968.4]
  assign _T_1840 = ~_T_1839; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@209969.4]
  assign _T_1842 = _T_1831 + 32'h1; // @[Monitor.scala 689:26:freechips.rocketchip.system.DefaultRV32Config.fir@209975.4]
  assign _T_1845 = _T_1477 | _T_1526; // @[Monitor.scala 690:27:freechips.rocketchip.system.DefaultRV32Config.fir@209979.4]
  assign _T_1857 = _T_1855 - 10'h1; // @[Edges.scala 231:28:freechips.rocketchip.system.DefaultRV32Config.fir@209994.4]
  assign _T_1858 = _T_1855 == 10'h0; // @[Edges.scala 232:25:freechips.rocketchip.system.DefaultRV32Config.fir@209995.4]
  assign _T_1868 = _T_1526 & _T_1858; // @[Monitor.scala 700:27:freechips.rocketchip.system.DefaultRV32Config.fir@210009.4]
  assign _T_1871 = ~io_in_d_bits_opcode[1]; // @[Edges.scala 72:43:freechips.rocketchip.system.DefaultRV32Config.fir@210012.4]
  assign _T_1872 = io_in_d_bits_opcode[2] & _T_1871; // @[Edges.scala 72:40:freechips.rocketchip.system.DefaultRV32Config.fir@210013.4]
  assign _T_1873 = _T_1868 & _T_1872; // @[Monitor.scala 700:38:freechips.rocketchip.system.DefaultRV32Config.fir@210014.4]
  assign _T_1874 = 4'h1 << io_in_d_bits_sink; // @[OneHot.scala 58:35:freechips.rocketchip.system.DefaultRV32Config.fir@210016.6]
  assign _T_1875 = _T_1846 >> io_in_d_bits_sink; // @[Monitor.scala 702:23:freechips.rocketchip.system.DefaultRV32Config.fir@210018.6]
  assign _T_1877 = ~_T_1875[0]; // @[Monitor.scala 702:14:freechips.rocketchip.system.DefaultRV32Config.fir@210020.6]
  assign _T_1879 = _T_1877 | reset; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@210022.6]
  assign _T_1880 = ~_T_1879; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@210023.6]
  assign _GEN_69 = _T_1873 ? _T_1874 : 4'h0; // @[Monitor.scala 700:72:freechips.rocketchip.system.DefaultRV32Config.fir@210015.4]
  assign _T_1882 = io_in_e_ready & io_in_e_valid; // @[Decoupled.scala 40:37:freechips.rocketchip.system.DefaultRV32Config.fir@210031.4]
  assign _T_1885 = 4'h1 << io_in_e_bits_sink; // @[OneHot.scala 58:35:freechips.rocketchip.system.DefaultRV32Config.fir@210035.6]
  assign _T_1886 = _GEN_69 | _T_1846; // @[Monitor.scala 708:24:freechips.rocketchip.system.DefaultRV32Config.fir@210037.6]
  assign _T_1887 = _T_1886 >> io_in_e_bits_sink; // @[Monitor.scala 708:35:freechips.rocketchip.system.DefaultRV32Config.fir@210038.6]
  assign _T_1890 = _T_1887[0] | reset; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@210041.6]
  assign _T_1891 = ~_T_1890; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@210042.6]
  assign _GEN_70 = _T_1882 ? _T_1885 : 4'h0; // @[Monitor.scala 706:73:freechips.rocketchip.system.DefaultRV32Config.fir@210034.4]
  assign _T_1892 = _T_1846 | _GEN_69; // @[Monitor.scala 713:27:freechips.rocketchip.system.DefaultRV32Config.fir@210048.4]
  assign _T_1893 = ~_GEN_70; // @[Monitor.scala 713:38:freechips.rocketchip.system.DefaultRV32Config.fir@210049.4]
  assign _T_1894 = _T_1892 & _T_1893; // @[Monitor.scala 713:36:freechips.rocketchip.system.DefaultRV32Config.fir@210050.4]
  assign _GEN_87 = io_in_a_valid & _T_78; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@207244.10]
  assign _GEN_103 = io_in_a_valid & _T_168; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@207373.10]
  assign _GEN_121 = io_in_a_valid & _T_262; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@207513.10]
  assign _GEN_133 = io_in_a_valid & _T_336; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@207620.10]
  assign _GEN_143 = io_in_a_valid & _T_413; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@207719.10]
  assign _GEN_153 = io_in_a_valid & _T_492; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@207810.10]
  assign _GEN_163 = io_in_a_valid & _T_559; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@207899.10]
  assign _GEN_173 = io_in_a_valid & _T_626; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@207988.10]
  assign _GEN_185 = io_in_d_valid & _T_708; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@208057.10]
  assign _GEN_195 = io_in_d_valid & _T_728; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@208099.10]
  assign _GEN_205 = io_in_d_valid & _T_756; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@208157.10]
  assign _GEN_215 = io_in_d_valid & _T_785; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@208216.10]
  assign _GEN_221 = io_in_d_valid & _T_802; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@208251.10]
  assign _GEN_227 = io_in_d_valid & _T_820; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@208287.10]
  assign _GEN_233 = io_in_b_valid & _T_962; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@208486.10]
  assign _GEN_247 = io_in_b_valid & _T_998; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@208541.10]
  assign _GEN_261 = io_in_b_valid & _T_1023; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@208596.10]
  assign _GEN_273 = io_in_b_valid & _T_1044; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@208643.10]
  assign _GEN_285 = io_in_b_valid & _T_1067; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@208692.10]
  assign _GEN_295 = io_in_b_valid & _T_1088; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@208739.10]
  assign _GEN_305 = io_in_b_valid & _T_1109; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@208786.10]
  assign _GEN_317 = io_in_c_valid & _T_1217; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@208942.10]
  assign _GEN_327 = io_in_c_valid & _T_1239; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@208990.10]
  assign _GEN_337 = io_in_c_valid & _T_1257; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@209079.10]
  assign _GEN_349 = io_in_c_valid & _T_1342; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@209199.10]
  assign _GEN_361 = io_in_c_valid & _T_1423; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@209262.10]
  assign _GEN_369 = io_in_c_valid & _T_1441; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@209302.10]
  assign _GEN_377 = io_in_c_valid & _T_1455; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@209334.10]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_1486 = _RAND_0[9:0];
  _RAND_1 = {1{`RANDOM}};
  _T_1497 = _RAND_1[2:0];
  _RAND_2 = {1{`RANDOM}};
  _T_1498 = _RAND_2[2:0];
  _RAND_3 = {1{`RANDOM}};
  _T_1499 = _RAND_3[3:0];
  _RAND_4 = {1{`RANDOM}};
  _T_1500 = _RAND_4[1:0];
  _RAND_5 = {1{`RANDOM}};
  _T_1501 = _RAND_5[31:0];
  _RAND_6 = {1{`RANDOM}};
  _T_1534 = _RAND_6[9:0];
  _RAND_7 = {1{`RANDOM}};
  _T_1545 = _RAND_7[2:0];
  _RAND_8 = {1{`RANDOM}};
  _T_1546 = _RAND_8[1:0];
  _RAND_9 = {1{`RANDOM}};
  _T_1547 = _RAND_9[3:0];
  _RAND_10 = {1{`RANDOM}};
  _T_1548 = _RAND_10[1:0];
  _RAND_11 = {1{`RANDOM}};
  _T_1549 = _RAND_11[1:0];
  _RAND_12 = {1{`RANDOM}};
  _T_1550 = _RAND_12[0:0];
  _RAND_13 = {1{`RANDOM}};
  _T_1588 = _RAND_13[9:0];
  _RAND_14 = {1{`RANDOM}};
  _T_1599 = _RAND_14[2:0];
  _RAND_15 = {1{`RANDOM}};
  _T_1600 = _RAND_15[1:0];
  _RAND_16 = {1{`RANDOM}};
  _T_1601 = _RAND_16[3:0];
  _RAND_17 = {1{`RANDOM}};
  _T_1602 = _RAND_17[1:0];
  _RAND_18 = {1{`RANDOM}};
  _T_1603 = _RAND_18[31:0];
  _RAND_19 = {1{`RANDOM}};
  _T_1636 = _RAND_19[9:0];
  _RAND_20 = {1{`RANDOM}};
  _T_1647 = _RAND_20[2:0];
  _RAND_21 = {1{`RANDOM}};
  _T_1648 = _RAND_21[2:0];
  _RAND_22 = {1{`RANDOM}};
  _T_1649 = _RAND_22[3:0];
  _RAND_23 = {1{`RANDOM}};
  _T_1650 = _RAND_23[1:0];
  _RAND_24 = {1{`RANDOM}};
  _T_1651 = _RAND_24[31:0];
  _RAND_25 = {1{`RANDOM}};
  inflight = _RAND_25[2:0];
  _RAND_26 = {1{`RANDOM}};
  inflight_opcodes = _RAND_26[11:0];
  _RAND_27 = {1{`RANDOM}};
  inflight_sizes = _RAND_27[23:0];
  _RAND_28 = {1{`RANDOM}};
  _T_1685 = _RAND_28[9:0];
  _RAND_29 = {1{`RANDOM}};
  _T_1703 = _RAND_29[9:0];
  _RAND_30 = {1{`RANDOM}};
  _T_1831 = _RAND_30[31:0];
  _RAND_31 = {1{`RANDOM}};
  _T_1846 = _RAND_31[3:0];
  _RAND_32 = {1{`RANDOM}};
  _T_1855 = _RAND_32[9:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      _T_1486 <= 10'h0;
    end else if (_T_1477) begin
      if (_T_1489) begin
        if (_T_1484) begin
          _T_1486 <= _T_13[11:2];
        end else begin
          _T_1486 <= 10'h0;
        end
      end else begin
        _T_1486 <= _T_1488;
      end
    end
    if (_T_1525) begin
      _T_1497 <= io_in_a_bits_opcode;
    end
    if (_T_1525) begin
      _T_1498 <= io_in_a_bits_param;
    end
    if (_T_1525) begin
      _T_1499 <= io_in_a_bits_size;
    end
    if (_T_1525) begin
      _T_1500 <= io_in_a_bits_source;
    end
    if (_T_1525) begin
      _T_1501 <= io_in_a_bits_address;
    end
    if (reset) begin
      _T_1534 <= 10'h0;
    end else if (_T_1526) begin
      if (_T_1537) begin
        if (io_in_d_bits_opcode[0]) begin
          _T_1534 <= _T_1530[11:2];
        end else begin
          _T_1534 <= 10'h0;
        end
      end else begin
        _T_1534 <= _T_1536;
      end
    end
    if (_T_1578) begin
      _T_1545 <= io_in_d_bits_opcode;
    end
    if (_T_1578) begin
      _T_1546 <= io_in_d_bits_param;
    end
    if (_T_1578) begin
      _T_1547 <= io_in_d_bits_size;
    end
    if (_T_1578) begin
      _T_1548 <= io_in_d_bits_source;
    end
    if (_T_1578) begin
      _T_1549 <= io_in_d_bits_sink;
    end
    if (_T_1578) begin
      _T_1550 <= io_in_d_bits_denied;
    end
    if (reset) begin
      _T_1588 <= 10'h0;
    end else if (_T_1579) begin
      if (_T_1591) begin
        _T_1588 <= 10'h0;
      end else begin
        _T_1588 <= _T_1590;
      end
    end
    if (_T_1627) begin
      _T_1599 <= io_in_b_bits_opcode;
    end
    if (_T_1627) begin
      _T_1600 <= io_in_b_bits_param;
    end
    if (_T_1627) begin
      _T_1601 <= io_in_b_bits_size;
    end
    if (_T_1627) begin
      _T_1602 <= io_in_b_bits_source;
    end
    if (_T_1627) begin
      _T_1603 <= io_in_b_bits_address;
    end
    if (reset) begin
      _T_1636 <= 10'h0;
    end else if (_T_1628) begin
      if (_T_1639) begin
        if (io_in_c_bits_opcode[0]) begin
          _T_1636 <= _T_1143[11:2];
        end else begin
          _T_1636 <= 10'h0;
        end
      end else begin
        _T_1636 <= _T_1638;
      end
    end
    if (_T_1675) begin
      _T_1647 <= io_in_c_bits_opcode;
    end
    if (_T_1675) begin
      _T_1648 <= io_in_c_bits_param;
    end
    if (_T_1675) begin
      _T_1649 <= io_in_c_bits_size;
    end
    if (_T_1675) begin
      _T_1650 <= io_in_c_bits_source;
    end
    if (_T_1675) begin
      _T_1651 <= io_in_c_bits_address;
    end
    if (reset) begin
      inflight <= 3'h0;
    end else begin
      inflight <= _T_1824;
    end
    if (reset) begin
      inflight_opcodes <= 12'h0;
    end else begin
      inflight_opcodes <= _T_1827;
    end
    if (reset) begin
      inflight_sizes <= 24'h0;
    end else begin
      inflight_sizes <= _T_1830;
    end
    if (reset) begin
      _T_1685 <= 10'h0;
    end else if (_T_1477) begin
      if (a_first) begin
        if (_T_1484) begin
          _T_1685 <= _T_13[11:2];
        end else begin
          _T_1685 <= 10'h0;
        end
      end else begin
        _T_1685 <= _T_1687;
      end
    end
    if (reset) begin
      _T_1703 <= 10'h0;
    end else if (_T_1526) begin
      if (d_first) begin
        if (io_in_d_bits_opcode[0]) begin
          _T_1703 <= _T_1530[11:2];
        end else begin
          _T_1703 <= 10'h0;
        end
      end else begin
        _T_1703 <= _T_1705;
      end
    end
    if (reset) begin
      _T_1831 <= 32'h0;
    end else if (_T_1845) begin
      _T_1831 <= 32'h0;
    end else begin
      _T_1831 <= _T_1842;
    end
    if (reset) begin
      _T_1846 <= 4'h0;
    end else begin
      _T_1846 <= _T_1894;
    end
    if (reset) begin
      _T_1855 <= 10'h0;
    end else if (_T_1526) begin
      if (_T_1858) begin
        if (io_in_d_bits_opcode[0]) begin
          _T_1855 <= _T_1530[11:2];
        end else begin
          _T_1855 <= 10'h0;
        end
      end else begin
        _T_1855 <= _T_1857;
      end
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_87 & _T_130) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel carries AcquireBlock type unsupported by manager (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@207244.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_87 & _T_130) begin
          $fatal; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@207245.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_87 & _T_144) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel carries AcquireBlock from a client which does not support Probe (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@207267.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_87 & _T_144) begin
          $fatal; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@207268.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_87 & _T_147) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel AcquireBlock carries invalid source ID (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@207274.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_87 & _T_147) begin
          $fatal; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@207275.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_87 & _T_151) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel AcquireBlock smaller than a beat (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@207282.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_87 & _T_151) begin
          $fatal; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@207283.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_87 & _T_154) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel AcquireBlock address not aligned to size (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@207289.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_87 & _T_154) begin
          $fatal; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@207290.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_87 & _T_158) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel AcquireBlock carries invalid grow param (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@207297.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_87 & _T_158) begin
          $fatal; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@207298.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_87 & _T_163) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel AcquireBlock contains invalid mask (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@207306.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_87 & _T_163) begin
          $fatal; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@207307.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_87 & _T_167) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel AcquireBlock is corrupt (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@207314.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_87 & _T_167) begin
          $fatal; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@207315.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_103 & _T_130) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel carries AcquirePerm type unsupported by manager (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@207373.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_103 & _T_130) begin
          $fatal; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@207374.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_103 & _T_144) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel carries AcquirePerm from a client which does not support Probe (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@207396.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_103 & _T_144) begin
          $fatal; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@207397.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_103 & _T_147) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel AcquirePerm carries invalid source ID (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@207403.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_103 & _T_147) begin
          $fatal; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@207404.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_103 & _T_151) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel AcquirePerm smaller than a beat (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@207411.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_103 & _T_151) begin
          $fatal; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@207412.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_103 & _T_154) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel AcquirePerm address not aligned to size (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@207418.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_103 & _T_154) begin
          $fatal; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@207419.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_103 & _T_158) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel AcquirePerm carries invalid grow param (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@207426.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_103 & _T_158) begin
          $fatal; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@207427.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_103 & _T_252) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel AcquirePerm requests NtoB (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@207434.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_103 & _T_252) begin
          $fatal; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@207435.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_103 & _T_163) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel AcquirePerm contains invalid mask (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@207443.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_103 & _T_163) begin
          $fatal; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@207444.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_103 & _T_167) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel AcquirePerm is corrupt (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@207451.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_103 & _T_167) begin
          $fatal; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@207452.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_121 & _T_317) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel carries Get type unsupported by manager (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@207513.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_121 & _T_317) begin
          $fatal; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@207514.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_121 & _T_147) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel Get carries invalid source ID (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@207520.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_121 & _T_147) begin
          $fatal; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@207521.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_121 & _T_154) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel Get address not aligned to size (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@207527.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_121 & _T_154) begin
          $fatal; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@207528.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_121 & _T_327) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel Get carries invalid param (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@207535.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_121 & _T_327) begin
          $fatal; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@207536.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_121 & _T_331) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel Get contains invalid mask (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@207543.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_121 & _T_331) begin
          $fatal; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@207544.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_121 & _T_167) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel Get is corrupt (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@207551.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_121 & _T_167) begin
          $fatal; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@207552.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_133 & _T_398) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel carries PutFull type unsupported by manager (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@207620.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_133 & _T_398) begin
          $fatal; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@207621.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_133 & _T_147) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel PutFull carries invalid source ID (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@207627.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_133 & _T_147) begin
          $fatal; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@207628.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_133 & _T_154) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel PutFull address not aligned to size (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@207634.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_133 & _T_154) begin
          $fatal; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@207635.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_133 & _T_327) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel PutFull carries invalid param (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@207642.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_133 & _T_327) begin
          $fatal; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@207643.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_133 & _T_331) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel PutFull contains invalid mask (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@207650.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_133 & _T_331) begin
          $fatal; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@207651.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_143 & _T_398) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel carries PutPartial type unsupported by manager (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@207719.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_143 & _T_398) begin
          $fatal; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@207720.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_143 & _T_147) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel PutPartial carries invalid source ID (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@207726.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_143 & _T_147) begin
          $fatal; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@207727.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_143 & _T_154) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel PutPartial address not aligned to size (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@207733.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_143 & _T_154) begin
          $fatal; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@207734.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_143 & _T_327) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel PutPartial carries invalid param (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@207741.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_143 & _T_327) begin
          $fatal; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@207742.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_143 & _T_491) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel PutPartial contains invalid mask (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@207751.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_143 & _T_491) begin
          $fatal; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@207752.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_153 & _T_544) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel carries Arithmetic type unsupported by manager (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@207810.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_153 & _T_544) begin
          $fatal; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@207811.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_153 & _T_147) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel Arithmetic carries invalid source ID (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@207817.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_153 & _T_147) begin
          $fatal; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@207818.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_153 & _T_154) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel Arithmetic address not aligned to size (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@207824.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_153 & _T_154) begin
          $fatal; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@207825.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_153 & _T_554) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel Arithmetic carries invalid opcode param (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@207832.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_153 & _T_554) begin
          $fatal; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@207833.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_153 & _T_331) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel Arithmetic contains invalid mask (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@207840.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_153 & _T_331) begin
          $fatal; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@207841.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_163 & _T_544) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel carries Logical type unsupported by manager (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@207899.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_163 & _T_544) begin
          $fatal; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@207900.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_163 & _T_147) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel Logical carries invalid source ID (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@207906.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_163 & _T_147) begin
          $fatal; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@207907.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_163 & _T_154) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel Logical address not aligned to size (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@207913.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_163 & _T_154) begin
          $fatal; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@207914.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_163 & _T_621) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel Logical carries invalid opcode param (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@207921.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_163 & _T_621) begin
          $fatal; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@207922.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_163 & _T_331) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel Logical contains invalid mask (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@207929.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_163 & _T_331) begin
          $fatal; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@207930.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_173 & _T_678) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel carries Hint type unsupported by manager (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@207988.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_173 & _T_678) begin
          $fatal; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@207989.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_173 & _T_147) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel Hint carries invalid source ID (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@207995.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_173 & _T_147) begin
          $fatal; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@207996.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_173 & _T_154) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel Hint address not aligned to size (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@208002.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_173 & _T_154) begin
          $fatal; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@208003.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_173 & _T_688) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel Hint carries invalid opcode param (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@208010.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_173 & _T_688) begin
          $fatal; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@208011.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_173 & _T_331) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel Hint contains invalid mask (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@208018.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_173 & _T_331) begin
          $fatal; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@208019.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_173 & _T_167) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel Hint is corrupt (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@208026.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_173 & _T_167) begin
          $fatal; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@208027.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_d_valid & _T_700) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel has invalid opcode (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:51 assert(cond, message)\n"); // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@208037.8]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_d_valid & _T_700) begin
          $fatal; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@208038.8]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_185 & _T_711) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel ReleaseAck carries invalid source ID (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:51 assert(cond, message)\n"); // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@208057.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_185 & _T_711) begin
          $fatal; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@208058.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_185 & _T_715) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel ReleaseAck smaller than a beat (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:51 assert(cond, message)\n"); // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@208065.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_185 & _T_715) begin
          $fatal; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@208066.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_185 & _T_719) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel ReleaseeAck carries invalid param (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:51 assert(cond, message)\n"); // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@208073.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_185 & _T_719) begin
          $fatal; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@208074.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_185 & _T_723) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel ReleaseAck is corrupt (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:51 assert(cond, message)\n"); // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@208081.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_185 & _T_723) begin
          $fatal; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@208082.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_185 & _T_727) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel ReleaseAck is denied (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:51 assert(cond, message)\n"); // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@208089.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_185 & _T_727) begin
          $fatal; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@208090.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_195 & _T_711) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel Grant carries invalid source ID (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:51 assert(cond, message)\n"); // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@208099.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_195 & _T_711) begin
          $fatal; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@208100.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_195 & _T_715) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel Grant smaller than a beat (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:51 assert(cond, message)\n"); // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@208114.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_195 & _T_715) begin
          $fatal; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@208115.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_195 & _T_742) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel Grant carries invalid cap param (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:51 assert(cond, message)\n"); // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@208122.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_195 & _T_742) begin
          $fatal; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@208123.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_195 & _T_746) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel Grant carries toN param (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:51 assert(cond, message)\n"); // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@208130.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_195 & _T_746) begin
          $fatal; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@208131.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_195 & _T_723) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel Grant is corrupt (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:51 assert(cond, message)\n"); // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@208138.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_195 & _T_723) begin
          $fatal; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@208139.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_205 & _T_711) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel GrantData carries invalid source ID (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:51 assert(cond, message)\n"); // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@208157.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_205 & _T_711) begin
          $fatal; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@208158.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_205 & _T_715) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel GrantData smaller than a beat (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:51 assert(cond, message)\n"); // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@208172.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_205 & _T_715) begin
          $fatal; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@208173.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_205 & _T_742) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel GrantData carries invalid cap param (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:51 assert(cond, message)\n"); // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@208180.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_205 & _T_742) begin
          $fatal; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@208181.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_205 & _T_746) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel GrantData carries toN param (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:51 assert(cond, message)\n"); // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@208188.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_205 & _T_746) begin
          $fatal; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@208189.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_205 & _T_779) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel GrantData is denied but not corrupt (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:51 assert(cond, message)\n"); // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@208197.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_205 & _T_779) begin
          $fatal; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@208198.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_215 & _T_711) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel AccessAck carries invalid source ID (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:51 assert(cond, message)\n"); // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@208216.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_215 & _T_711) begin
          $fatal; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@208217.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_215 & _T_719) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel AccessAck carries invalid param (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:51 assert(cond, message)\n"); // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@208224.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_215 & _T_719) begin
          $fatal; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@208225.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_215 & _T_723) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel AccessAck is corrupt (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:51 assert(cond, message)\n"); // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@208232.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_215 & _T_723) begin
          $fatal; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@208233.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_221 & _T_711) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel AccessAckData carries invalid source ID (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:51 assert(cond, message)\n"); // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@208251.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_221 & _T_711) begin
          $fatal; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@208252.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_221 & _T_719) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel AccessAckData carries invalid param (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:51 assert(cond, message)\n"); // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@208259.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_221 & _T_719) begin
          $fatal; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@208260.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_221 & _T_779) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel AccessAckData is denied but not corrupt (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:51 assert(cond, message)\n"); // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@208268.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_221 & _T_779) begin
          $fatal; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@208269.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_227 & _T_711) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel HintAck carries invalid source ID (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:51 assert(cond, message)\n"); // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@208287.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_227 & _T_711) begin
          $fatal; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@208288.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_227 & _T_719) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel HintAck carries invalid param (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:51 assert(cond, message)\n"); // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@208295.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_227 & _T_719) begin
          $fatal; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@208296.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_227 & _T_723) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel HintAck is corrupt (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:51 assert(cond, message)\n"); // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@208303.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_227 & _T_723) begin
          $fatal; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@208304.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_b_valid & _T_840) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel has invalid opcode (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@208323.8]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_b_valid & _T_840) begin
          $fatal; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@208324.8]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_233 & _T_976) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel carries Probe type unsupported by client (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@208486.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_233 & _T_976) begin
          $fatal; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@208487.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_233 & _T_979) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel Probe carries unmanaged address (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@208493.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_233 & _T_979) begin
          $fatal; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@208494.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_233 & _T_982) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel Probe carries source that is not first source (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@208500.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_233 & _T_982) begin
          $fatal; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@208501.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_233 & _T_985) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel Probe address not aligned to size (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@208507.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_233 & _T_985) begin
          $fatal; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@208508.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_233 & _T_989) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel Probe carries invalid cap param (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@208515.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_233 & _T_989) begin
          $fatal; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@208516.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_233 & _T_993) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel Probe contains invalid mask (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@208523.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_233 & _T_993) begin
          $fatal; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@208524.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_233 & _T_997) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel Probe is corrupt (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@208531.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_233 & _T_997) begin
          $fatal; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@208532.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_247 & _T_1001) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel carries Get type unsupported by client (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@208541.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_247 & _T_1001) begin
          $fatal; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@208542.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_247 & _T_979) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel Get carries unmanaged address (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@208548.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_247 & _T_979) begin
          $fatal; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@208549.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_247 & _T_982) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel Get carries source that is not first source (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@208555.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_247 & _T_982) begin
          $fatal; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@208556.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_247 & _T_985) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel Get address not aligned to size (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@208562.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_247 & _T_985) begin
          $fatal; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@208563.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_247 & _T_1014) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel Get carries invalid param (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@208570.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_247 & _T_1014) begin
          $fatal; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@208571.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_247 & _T_993) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel Get contains invalid mask (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@208578.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_247 & _T_993) begin
          $fatal; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@208579.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_247 & _T_997) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel Get is corrupt (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@208586.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_247 & _T_997) begin
          $fatal; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@208587.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_261 & _T_1001) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel carries PutFull type unsupported by client (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@208596.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_261 & _T_1001) begin
          $fatal; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@208597.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_261 & _T_979) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel PutFull carries unmanaged address (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@208603.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_261 & _T_979) begin
          $fatal; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@208604.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_261 & _T_982) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel PutFull carries source that is not first source (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@208610.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_261 & _T_982) begin
          $fatal; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@208611.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_261 & _T_985) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel PutFull address not aligned to size (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@208617.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_261 & _T_985) begin
          $fatal; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@208618.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_261 & _T_1014) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel PutFull carries invalid param (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@208625.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_261 & _T_1014) begin
          $fatal; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@208626.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_261 & _T_993) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel PutFull contains invalid mask (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@208633.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_261 & _T_993) begin
          $fatal; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@208634.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_273 & _T_1001) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel carries PutPartial type unsupported by client (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@208643.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_273 & _T_1001) begin
          $fatal; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@208644.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_273 & _T_979) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel PutPartial carries unmanaged address (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@208650.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_273 & _T_979) begin
          $fatal; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@208651.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_273 & _T_982) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel PutPartial carries source that is not first source (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@208657.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_273 & _T_982) begin
          $fatal; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@208658.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_273 & _T_985) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel PutPartial address not aligned to size (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@208664.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_273 & _T_985) begin
          $fatal; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@208665.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_273 & _T_1014) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel PutPartial carries invalid param (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@208672.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_273 & _T_1014) begin
          $fatal; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@208673.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_273 & _T_1066) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel PutPartial contains invalid mask (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@208682.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_273 & _T_1066) begin
          $fatal; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@208683.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_285 & _T_1001) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel carries Arithmetic type unsupported by client (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@208692.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_285 & _T_1001) begin
          $fatal; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@208693.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_285 & _T_979) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel Arithmetic carries unmanaged address (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@208699.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_285 & _T_979) begin
          $fatal; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@208700.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_285 & _T_982) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel Arithmetic carries source that is not first source (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@208706.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_285 & _T_982) begin
          $fatal; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@208707.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_285 & _T_985) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel Arithmetic address not aligned to size (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@208713.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_285 & _T_985) begin
          $fatal; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@208714.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_285 & _T_993) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel Arithmetic contains invalid mask (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@208729.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_285 & _T_993) begin
          $fatal; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@208730.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_295 & _T_1001) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel carries Logical type unsupported by client (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@208739.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_295 & _T_1001) begin
          $fatal; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@208740.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_295 & _T_979) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel Logical carries unmanaged address (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@208746.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_295 & _T_979) begin
          $fatal; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@208747.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_295 & _T_982) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel Logical carries source that is not first source (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@208753.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_295 & _T_982) begin
          $fatal; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@208754.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_295 & _T_985) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel Logical address not aligned to size (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@208760.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_295 & _T_985) begin
          $fatal; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@208761.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_295 & _T_993) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel Logical contains invalid mask (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@208776.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_295 & _T_993) begin
          $fatal; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@208777.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_305 & _T_1001) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel carries Hint type unsupported by client (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@208786.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_305 & _T_1001) begin
          $fatal; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@208787.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_305 & _T_979) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel Hint carries unmanaged address (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@208793.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_305 & _T_979) begin
          $fatal; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@208794.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_305 & _T_982) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel Hint carries source that is not first source (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@208800.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_305 & _T_982) begin
          $fatal; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@208801.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_305 & _T_985) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel Hint address not aligned to size (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@208807.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_305 & _T_985) begin
          $fatal; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@208808.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_305 & _T_993) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel Hint contains invalid mask (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@208815.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_305 & _T_993) begin
          $fatal; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@208816.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_305 & _T_997) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel Hint is corrupt (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@208823.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_305 & _T_997) begin
          $fatal; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@208824.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_317 & _T_1220) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel ProbeAck carries unmanaged address (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@208942.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_317 & _T_1220) begin
          $fatal; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@208943.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_317 & _T_1223) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel ProbeAck carries invalid source ID (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@208949.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_317 & _T_1223) begin
          $fatal; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@208950.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_317 & _T_1227) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel ProbeAck smaller than a beat (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@208957.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_317 & _T_1227) begin
          $fatal; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@208958.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_317 & _T_1230) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel ProbeAck address not aligned to size (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@208964.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_317 & _T_1230) begin
          $fatal; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@208965.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_317 & _T_1234) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel ProbeAck carries invalid report param (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@208972.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_317 & _T_1234) begin
          $fatal; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@208973.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_327 & _T_1220) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel ProbeAckData carries unmanaged address (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@208990.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_327 & _T_1220) begin
          $fatal; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@208991.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_327 & _T_1223) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel ProbeAckData carries invalid source ID (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@208997.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_327 & _T_1223) begin
          $fatal; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@208998.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_327 & _T_1227) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel ProbeAckData smaller than a beat (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@209005.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_327 & _T_1227) begin
          $fatal; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@209006.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_327 & _T_1230) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel ProbeAckData address not aligned to size (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@209012.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_327 & _T_1230) begin
          $fatal; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@209013.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_327 & _T_1234) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel ProbeAckData carries invalid report param (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@209020.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_327 & _T_1234) begin
          $fatal; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@209021.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_337 & _T_1309) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel carries Release type unsupported by manager (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@209079.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_337 & _T_1309) begin
          $fatal; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@209080.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_337 & _T_1323) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel carries Release from a client which does not support Probe (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@209102.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_337 & _T_1323) begin
          $fatal; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@209103.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_337 & _T_1223) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel Release carries invalid source ID (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@209109.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_337 & _T_1223) begin
          $fatal; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@209110.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_337 & _T_1227) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel Release smaller than a beat (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@209117.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_337 & _T_1227) begin
          $fatal; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@209118.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_337 & _T_1230) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel Release address not aligned to size (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@209124.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_337 & _T_1230) begin
          $fatal; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@209125.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_337 & _T_1337) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel Release carries invalid shrink param (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@209132.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_337 & _T_1337) begin
          $fatal; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@209133.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_349 & _T_1309) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel carries ReleaseData type unsupported by manager (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@209199.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_349 & _T_1309) begin
          $fatal; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@209200.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_349 & _T_1323) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel carries Release from a client which does not support Probe (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@209222.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_349 & _T_1323) begin
          $fatal; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@209223.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_349 & _T_1223) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel ReleaseData carries invalid source ID (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@209229.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_349 & _T_1223) begin
          $fatal; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@209230.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_349 & _T_1227) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel ReleaseData smaller than a beat (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@209237.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_349 & _T_1227) begin
          $fatal; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@209238.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_349 & _T_1230) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel ReleaseData address not aligned to size (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@209244.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_349 & _T_1230) begin
          $fatal; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@209245.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_349 & _T_1337) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel ReleaseData carries invalid shrink param (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@209252.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_349 & _T_1337) begin
          $fatal; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@209253.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_361 & _T_1220) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel AccessAck carries unmanaged address (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@209262.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_361 & _T_1220) begin
          $fatal; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@209263.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_361 & _T_1223) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel AccessAck carries invalid source ID (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@209269.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_361 & _T_1223) begin
          $fatal; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@209270.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_361 & _T_1230) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel AccessAck address not aligned to size (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@209276.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_361 & _T_1230) begin
          $fatal; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@209277.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_361 & _T_1436) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel AccessAck carries invalid param (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@209284.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_361 & _T_1436) begin
          $fatal; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@209285.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_369 & _T_1220) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel AccessAckData carries unmanaged address (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@209302.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_369 & _T_1220) begin
          $fatal; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@209303.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_369 & _T_1223) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel AccessAckData carries invalid source ID (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@209309.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_369 & _T_1223) begin
          $fatal; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@209310.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_369 & _T_1230) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel AccessAckData address not aligned to size (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@209316.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_369 & _T_1230) begin
          $fatal; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@209317.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_369 & _T_1436) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel AccessAckData carries invalid param (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@209324.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_369 & _T_1436) begin
          $fatal; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@209325.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_377 & _T_1220) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel HintAck carries unmanaged address (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@209334.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_377 & _T_1220) begin
          $fatal; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@209335.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_377 & _T_1223) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel HintAck carries invalid source ID (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@209341.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_377 & _T_1223) begin
          $fatal; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@209342.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_377 & _T_1230) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel HintAck address not aligned to size (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@209348.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_377 & _T_1230) begin
          $fatal; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@209349.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_377 & _T_1436) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel HintAck carries invalid param (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@209356.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_377 & _T_1436) begin
          $fatal; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@209357.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1503 & _T_1507) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel opcode changed within multibeat operation (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@209415.8]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_1503 & _T_1507) begin
          $fatal; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@209416.8]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1503 & _T_1511) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel param changed within multibeat operation (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@209423.8]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_1503 & _T_1511) begin
          $fatal; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@209424.8]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1503 & _T_1515) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel size changed within multibeat operation (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@209431.8]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_1503 & _T_1515) begin
          $fatal; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@209432.8]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1503 & _T_1519) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel source changed within multibeat operation (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@209439.8]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_1503 & _T_1519) begin
          $fatal; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@209440.8]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1503 & _T_1523) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel address changed with multibeat operation (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@209447.8]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_1503 & _T_1523) begin
          $fatal; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@209448.8]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1552 & _T_1556) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel opcode changed within multibeat operation (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:51 assert(cond, message)\n"); // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@209496.8]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_1552 & _T_1556) begin
          $fatal; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@209497.8]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1552 & _T_1560) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel param changed within multibeat operation (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:51 assert(cond, message)\n"); // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@209504.8]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_1552 & _T_1560) begin
          $fatal; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@209505.8]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1552 & _T_1564) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel size changed within multibeat operation (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:51 assert(cond, message)\n"); // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@209512.8]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_1552 & _T_1564) begin
          $fatal; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@209513.8]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1552 & _T_1568) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel source changed within multibeat operation (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:51 assert(cond, message)\n"); // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@209520.8]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_1552 & _T_1568) begin
          $fatal; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@209521.8]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1552 & _T_1572) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel sink changed with multibeat operation (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:51 assert(cond, message)\n"); // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@209528.8]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_1552 & _T_1572) begin
          $fatal; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@209529.8]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1552 & _T_1576) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel denied changed with multibeat operation (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:51 assert(cond, message)\n"); // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@209536.8]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_1552 & _T_1576) begin
          $fatal; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@209537.8]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1605 & _T_1609) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel opcode changed within multibeat operation (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@209586.8]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_1605 & _T_1609) begin
          $fatal; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@209587.8]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1605 & _T_1613) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel param changed within multibeat operation (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@209594.8]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_1605 & _T_1613) begin
          $fatal; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@209595.8]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1605 & _T_1617) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel size changed within multibeat operation (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@209602.8]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_1605 & _T_1617) begin
          $fatal; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@209603.8]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1605 & _T_1621) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel source changed within multibeat operation (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@209610.8]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_1605 & _T_1621) begin
          $fatal; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@209611.8]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1605 & _T_1625) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel addresss changed with multibeat operation (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@209618.8]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_1605 & _T_1625) begin
          $fatal; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@209619.8]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1653 & _T_1657) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel opcode changed within multibeat operation (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@209666.8]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_1653 & _T_1657) begin
          $fatal; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@209667.8]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1653 & _T_1661) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel param changed within multibeat operation (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@209674.8]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_1653 & _T_1661) begin
          $fatal; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@209675.8]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1653 & _T_1665) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel size changed within multibeat operation (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@209682.8]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_1653 & _T_1665) begin
          $fatal; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@209683.8]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1653 & _T_1669) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel source changed within multibeat operation (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@209690.8]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_1653 & _T_1669) begin
          $fatal; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@209691.8]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1653 & _T_1673) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel address changed with multibeat operation (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@209698.8]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_1653 & _T_1673) begin
          $fatal; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@209699.8]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1732 & _T_1748) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel re-used a source ID (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@209834.8]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_1732 & _T_1748) begin
          $fatal; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@209835.8]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1771 & _T_1782) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel acknowledged for nothing inflight (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:51 assert(cond, message)\n"); // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@209885.8]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_1771 & _T_1782) begin
          $fatal; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@209886.8]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1771 & _T_1795) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel contains improper opcode response (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:51 assert(cond, message)\n"); // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@209902.8]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_1771 & _T_1795) begin
          $fatal; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@209903.8]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1771 & _T_1802) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel contains improper response size (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:51 assert(cond, message)\n"); // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@209913.8]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_1771 & _T_1802) begin
          $fatal; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@209914.8]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1809 & _T_1814) begin
          $fwrite(32'h80000002,"Assertion failed: ready check\n    at Monitor.scala:51 assert(cond, message)\n"); // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@209931.8]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_1809 & _T_1814) begin
          $fatal; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@209932.8]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1821) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' and 'D' concurrent, despite minlatency 3 (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:51 assert(cond, message)\n"); // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@209943.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_1821) begin
          $fatal; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@209944.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1840) begin
          $fwrite(32'h80000002,"Assertion failed: TileLink timeout expired (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@209971.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_1840) begin
          $fatal; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@209972.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1873 & _T_1880) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel re-used a sink ID (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:51 assert(cond, message)\n"); // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@210025.8]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_1873 & _T_1880) begin
          $fatal; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@210026.8]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1882 & _T_1891) begin
          $fwrite(32'h80000002,"Assertion failed: 'E' channel acknowledged for nothing inflight (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@210044.8]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_1882 & _T_1891) begin
          $fatal; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@210045.8]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
  end
endmodule
