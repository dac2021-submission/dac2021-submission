module SimpleClockGroupSource( // @[:freechips.rocketchip.system.DefaultRV32Config.fir@20.2]
  input   clock, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@21.4]
  input   reset, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@22.4]
  output  auto_out_member_5_clock, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@23.4]
  output  auto_out_member_5_reset, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@23.4]
  output  auto_out_member_4_clock, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@23.4]
  output  auto_out_member_4_reset, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@23.4]
  output  auto_out_member_3_clock, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@23.4]
  output  auto_out_member_3_reset, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@23.4]
  output  auto_out_member_2_clock, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@23.4]
  output  auto_out_member_2_reset, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@23.4]
  output  auto_out_member_1_clock, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@23.4]
  output  auto_out_member_1_reset, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@23.4]
  output  auto_out_member_0_clock, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@23.4]
  output  auto_out_member_0_reset // @[:freechips.rocketchip.system.DefaultRV32Config.fir@23.4]
);
  assign auto_out_member_5_clock = clock; // @[LazyModule.scala 305:12:freechips.rocketchip.system.DefaultRV32Config.fir@30.4]
  assign auto_out_member_5_reset = reset; // @[LazyModule.scala 305:12:freechips.rocketchip.system.DefaultRV32Config.fir@30.4]
  assign auto_out_member_4_clock = clock; // @[LazyModule.scala 305:12:freechips.rocketchip.system.DefaultRV32Config.fir@30.4]
  assign auto_out_member_4_reset = reset; // @[LazyModule.scala 305:12:freechips.rocketchip.system.DefaultRV32Config.fir@30.4]
  assign auto_out_member_3_clock = clock; // @[LazyModule.scala 305:12:freechips.rocketchip.system.DefaultRV32Config.fir@30.4]
  assign auto_out_member_3_reset = reset; // @[LazyModule.scala 305:12:freechips.rocketchip.system.DefaultRV32Config.fir@30.4]
  assign auto_out_member_2_clock = clock; // @[LazyModule.scala 305:12:freechips.rocketchip.system.DefaultRV32Config.fir@30.4]
  assign auto_out_member_2_reset = reset; // @[LazyModule.scala 305:12:freechips.rocketchip.system.DefaultRV32Config.fir@30.4]
  assign auto_out_member_1_clock = clock; // @[LazyModule.scala 305:12:freechips.rocketchip.system.DefaultRV32Config.fir@30.4]
  assign auto_out_member_1_reset = reset; // @[LazyModule.scala 305:12:freechips.rocketchip.system.DefaultRV32Config.fir@30.4]
  assign auto_out_member_0_clock = clock; // @[LazyModule.scala 305:12:freechips.rocketchip.system.DefaultRV32Config.fir@30.4]
  assign auto_out_member_0_reset = reset; // @[LazyModule.scala 305:12:freechips.rocketchip.system.DefaultRV32Config.fir@30.4]
endmodule
