module TLMonitor_3( // @[:freechips.rocketchip.system.DefaultRV32Config.fir@9350.2]
  input         clock, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@9351.4]
  input         reset, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@9352.4]
  input         io_in_a_ready, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@9353.4]
  input         io_in_a_valid, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@9353.4]
  input  [2:0]  io_in_a_bits_opcode, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@9353.4]
  input  [2:0]  io_in_a_bits_param, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@9353.4]
  input  [3:0]  io_in_a_bits_size, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@9353.4]
  input  [1:0]  io_in_a_bits_source, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@9353.4]
  input  [31:0] io_in_a_bits_address, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@9353.4]
  input  [3:0]  io_in_a_bits_mask, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@9353.4]
  input         io_in_a_bits_corrupt, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@9353.4]
  input         io_in_b_ready, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@9353.4]
  input         io_in_b_valid, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@9353.4]
  input  [1:0]  io_in_b_bits_param, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@9353.4]
  input  [31:0] io_in_b_bits_address, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@9353.4]
  input         io_in_c_ready, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@9353.4]
  input         io_in_c_valid, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@9353.4]
  input  [2:0]  io_in_c_bits_opcode, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@9353.4]
  input  [2:0]  io_in_c_bits_param, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@9353.4]
  input  [3:0]  io_in_c_bits_size, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@9353.4]
  input  [1:0]  io_in_c_bits_source, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@9353.4]
  input  [31:0] io_in_c_bits_address, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@9353.4]
  input         io_in_c_bits_corrupt, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@9353.4]
  input         io_in_d_ready, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@9353.4]
  input         io_in_d_valid, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@9353.4]
  input  [2:0]  io_in_d_bits_opcode, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@9353.4]
  input  [1:0]  io_in_d_bits_param, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@9353.4]
  input  [3:0]  io_in_d_bits_size, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@9353.4]
  input  [1:0]  io_in_d_bits_source, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@9353.4]
  input  [1:0]  io_in_d_bits_sink, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@9353.4]
  input         io_in_d_bits_denied, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@9353.4]
  input         io_in_d_bits_corrupt, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@9353.4]
  input         io_in_e_valid, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@9353.4]
  input  [1:0]  io_in_e_bits_sink // @[:freechips.rocketchip.system.DefaultRV32Config.fir@9353.4]
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
`endif // RANDOMIZE_REG_INIT
  wire [31:0] plusarg_reader_out; // @[PlusArg.scala 80:11:freechips.rocketchip.system.DefaultRV32Config.fir@12216.4]
  wire  _T_4; // @[Parameters.scala 47:9:freechips.rocketchip.system.DefaultRV32Config.fir@9364.6]
  wire  _T_5; // @[Parameters.scala 47:9:freechips.rocketchip.system.DefaultRV32Config.fir@9365.6]
  wire  _T_6; // @[Parameters.scala 47:9:freechips.rocketchip.system.DefaultRV32Config.fir@9366.6]
  wire  _T_8; // @[Parameters.scala 924:46:freechips.rocketchip.system.DefaultRV32Config.fir@9372.6]
  wire  _T_9; // @[Parameters.scala 924:46:freechips.rocketchip.system.DefaultRV32Config.fir@9373.6]
  wire [26:0] _T_11; // @[package.scala 207:77:freechips.rocketchip.system.DefaultRV32Config.fir@9375.6]
  wire [11:0] _T_13; // @[package.scala 207:46:freechips.rocketchip.system.DefaultRV32Config.fir@9377.6]
  wire [31:0] _GEN_71; // @[Edges.scala 22:16:freechips.rocketchip.system.DefaultRV32Config.fir@9378.6]
  wire [31:0] _T_14; // @[Edges.scala 22:16:freechips.rocketchip.system.DefaultRV32Config.fir@9378.6]
  wire  _T_15; // @[Edges.scala 22:24:freechips.rocketchip.system.DefaultRV32Config.fir@9379.6]
  wire [1:0] _T_18; // @[OneHot.scala 65:12:freechips.rocketchip.system.DefaultRV32Config.fir@9382.6]
  wire [1:0] _T_20; // @[Misc.scala 201:81:freechips.rocketchip.system.DefaultRV32Config.fir@9384.6]
  wire  _T_21; // @[Misc.scala 205:21:freechips.rocketchip.system.DefaultRV32Config.fir@9385.6]
  wire  _T_24; // @[Misc.scala 210:20:freechips.rocketchip.system.DefaultRV32Config.fir@9388.6]
  wire  _T_26; // @[Misc.scala 214:38:freechips.rocketchip.system.DefaultRV32Config.fir@9390.6]
  wire  _T_27; // @[Misc.scala 214:29:freechips.rocketchip.system.DefaultRV32Config.fir@9391.6]
  wire  _T_29; // @[Misc.scala 214:38:freechips.rocketchip.system.DefaultRV32Config.fir@9393.6]
  wire  _T_30; // @[Misc.scala 214:29:freechips.rocketchip.system.DefaultRV32Config.fir@9394.6]
  wire  _T_33; // @[Misc.scala 210:20:freechips.rocketchip.system.DefaultRV32Config.fir@9397.6]
  wire  _T_34; // @[Misc.scala 213:27:freechips.rocketchip.system.DefaultRV32Config.fir@9398.6]
  wire  _T_35; // @[Misc.scala 214:38:freechips.rocketchip.system.DefaultRV32Config.fir@9399.6]
  wire  _T_36; // @[Misc.scala 214:29:freechips.rocketchip.system.DefaultRV32Config.fir@9400.6]
  wire  _T_37; // @[Misc.scala 213:27:freechips.rocketchip.system.DefaultRV32Config.fir@9401.6]
  wire  _T_38; // @[Misc.scala 214:38:freechips.rocketchip.system.DefaultRV32Config.fir@9402.6]
  wire  _T_39; // @[Misc.scala 214:29:freechips.rocketchip.system.DefaultRV32Config.fir@9403.6]
  wire  _T_40; // @[Misc.scala 213:27:freechips.rocketchip.system.DefaultRV32Config.fir@9404.6]
  wire  _T_41; // @[Misc.scala 214:38:freechips.rocketchip.system.DefaultRV32Config.fir@9405.6]
  wire  _T_42; // @[Misc.scala 214:29:freechips.rocketchip.system.DefaultRV32Config.fir@9406.6]
  wire  _T_43; // @[Misc.scala 213:27:freechips.rocketchip.system.DefaultRV32Config.fir@9407.6]
  wire  _T_44; // @[Misc.scala 214:38:freechips.rocketchip.system.DefaultRV32Config.fir@9408.6]
  wire  _T_45; // @[Misc.scala 214:29:freechips.rocketchip.system.DefaultRV32Config.fir@9409.6]
  wire [3:0] _T_48; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@9412.6]
  wire [32:0] _T_52; // @[Parameters.scala 137:49:freechips.rocketchip.system.DefaultRV32Config.fir@9416.6]
  wire  _T_78; // @[Monitor.scala 79:25:freechips.rocketchip.system.DefaultRV32Config.fir@9446.6]
  wire [32:0] _T_83; // @[Parameters.scala 137:52:freechips.rocketchip.system.DefaultRV32Config.fir@9452.8]
  wire  _T_84; // @[Parameters.scala 137:67:freechips.rocketchip.system.DefaultRV32Config.fir@9453.8]
  wire [31:0] _T_85; // @[Parameters.scala 137:31:freechips.rocketchip.system.DefaultRV32Config.fir@9454.8]
  wire [32:0] _T_86; // @[Parameters.scala 137:49:freechips.rocketchip.system.DefaultRV32Config.fir@9455.8]
  wire [32:0] _T_88; // @[Parameters.scala 137:52:freechips.rocketchip.system.DefaultRV32Config.fir@9457.8]
  wire  _T_89; // @[Parameters.scala 137:67:freechips.rocketchip.system.DefaultRV32Config.fir@9458.8]
  wire [31:0] _T_90; // @[Parameters.scala 137:31:freechips.rocketchip.system.DefaultRV32Config.fir@9459.8]
  wire [32:0] _T_91; // @[Parameters.scala 137:49:freechips.rocketchip.system.DefaultRV32Config.fir@9460.8]
  wire [32:0] _T_93; // @[Parameters.scala 137:52:freechips.rocketchip.system.DefaultRV32Config.fir@9462.8]
  wire  _T_94; // @[Parameters.scala 137:67:freechips.rocketchip.system.DefaultRV32Config.fir@9463.8]
  wire [31:0] _T_95; // @[Parameters.scala 137:31:freechips.rocketchip.system.DefaultRV32Config.fir@9464.8]
  wire [32:0] _T_96; // @[Parameters.scala 137:49:freechips.rocketchip.system.DefaultRV32Config.fir@9465.8]
  wire [32:0] _T_98; // @[Parameters.scala 137:52:freechips.rocketchip.system.DefaultRV32Config.fir@9467.8]
  wire  _T_99; // @[Parameters.scala 137:67:freechips.rocketchip.system.DefaultRV32Config.fir@9468.8]
  wire [31:0] _T_100; // @[Parameters.scala 137:31:freechips.rocketchip.system.DefaultRV32Config.fir@9469.8]
  wire [32:0] _T_101; // @[Parameters.scala 137:49:freechips.rocketchip.system.DefaultRV32Config.fir@9470.8]
  wire [32:0] _T_103; // @[Parameters.scala 137:52:freechips.rocketchip.system.DefaultRV32Config.fir@9472.8]
  wire  _T_104; // @[Parameters.scala 137:67:freechips.rocketchip.system.DefaultRV32Config.fir@9473.8]
  wire [31:0] _T_105; // @[Parameters.scala 137:31:freechips.rocketchip.system.DefaultRV32Config.fir@9474.8]
  wire [32:0] _T_106; // @[Parameters.scala 137:49:freechips.rocketchip.system.DefaultRV32Config.fir@9475.8]
  wire [32:0] _T_108; // @[Parameters.scala 137:52:freechips.rocketchip.system.DefaultRV32Config.fir@9477.8]
  wire  _T_109; // @[Parameters.scala 137:67:freechips.rocketchip.system.DefaultRV32Config.fir@9478.8]
  wire  _T_110; // @[Parameters.scala 552:42:freechips.rocketchip.system.DefaultRV32Config.fir@9479.8]
  wire  _T_117; // @[Parameters.scala 93:42:freechips.rocketchip.system.DefaultRV32Config.fir@9486.8]
  wire [31:0] _T_120; // @[Parameters.scala 137:31:freechips.rocketchip.system.DefaultRV32Config.fir@9489.8]
  wire [32:0] _T_121; // @[Parameters.scala 137:49:freechips.rocketchip.system.DefaultRV32Config.fir@9490.8]
  wire [32:0] _T_123; // @[Parameters.scala 137:52:freechips.rocketchip.system.DefaultRV32Config.fir@9492.8]
  wire  _T_124; // @[Parameters.scala 137:67:freechips.rocketchip.system.DefaultRV32Config.fir@9493.8]
  wire  _T_125; // @[Parameters.scala 551:56:freechips.rocketchip.system.DefaultRV32Config.fir@9494.8]
  wire  _T_129; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@9498.8]
  wire  _T_130; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@9499.8]
  wire  _T_135; // @[Parameters.scala 92:48:freechips.rocketchip.system.DefaultRV32Config.fir@9512.8]
  wire  _T_136; // @[Mux.scala 27:72:freechips.rocketchip.system.DefaultRV32Config.fir@9513.8]
  wire  _T_143; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@9521.8]
  wire  _T_144; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@9522.8]
  wire  _T_146; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@9528.8]
  wire  _T_147; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@9529.8]
  wire  _T_150; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@9536.8]
  wire  _T_151; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@9537.8]
  wire  _T_153; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@9543.8]
  wire  _T_154; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@9544.8]
  wire  _T_155; // @[Bundles.scala 110:27:freechips.rocketchip.system.DefaultRV32Config.fir@9549.8]
  wire  _T_157; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@9551.8]
  wire  _T_158; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@9552.8]
  wire [3:0] _T_159; // @[Monitor.scala 86:18:freechips.rocketchip.system.DefaultRV32Config.fir@9557.8]
  wire  _T_160; // @[Monitor.scala 86:31:freechips.rocketchip.system.DefaultRV32Config.fir@9558.8]
  wire  _T_162; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@9560.8]
  wire  _T_163; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@9561.8]
  wire  _T_164; // @[Monitor.scala 87:18:freechips.rocketchip.system.DefaultRV32Config.fir@9566.8]
  wire  _T_166; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@9568.8]
  wire  _T_167; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@9569.8]
  wire  _T_168; // @[Monitor.scala 90:25:freechips.rocketchip.system.DefaultRV32Config.fir@9575.6]
  wire  _T_249; // @[Monitor.scala 97:31:freechips.rocketchip.system.DefaultRV32Config.fir@9686.8]
  wire  _T_251; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@9688.8]
  wire  _T_252; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@9689.8]
  wire  _T_262; // @[Monitor.scala 102:25:freechips.rocketchip.system.DefaultRV32Config.fir@9712.6]
  wire  _T_264; // @[Parameters.scala 93:42:freechips.rocketchip.system.DefaultRV32Config.fir@9715.8]
  wire  _T_272; // @[Parameters.scala 551:56:freechips.rocketchip.system.DefaultRV32Config.fir@9723.8]
  wire  _T_307; // @[Parameters.scala 552:42:freechips.rocketchip.system.DefaultRV32Config.fir@9758.8]
  wire  _T_308; // @[Parameters.scala 552:42:freechips.rocketchip.system.DefaultRV32Config.fir@9759.8]
  wire  _T_309; // @[Parameters.scala 552:42:freechips.rocketchip.system.DefaultRV32Config.fir@9760.8]
  wire  _T_310; // @[Parameters.scala 552:42:freechips.rocketchip.system.DefaultRV32Config.fir@9761.8]
  wire  _T_311; // @[Parameters.scala 552:42:freechips.rocketchip.system.DefaultRV32Config.fir@9762.8]
  wire  _T_312; // @[Parameters.scala 551:56:freechips.rocketchip.system.DefaultRV32Config.fir@9763.8]
  wire  _T_314; // @[Parameters.scala 553:30:freechips.rocketchip.system.DefaultRV32Config.fir@9765.8]
  wire  _T_316; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@9767.8]
  wire  _T_317; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@9768.8]
  wire  _T_324; // @[Monitor.scala 106:31:freechips.rocketchip.system.DefaultRV32Config.fir@9787.8]
  wire  _T_326; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@9789.8]
  wire  _T_327; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@9790.8]
  wire  _T_328; // @[Monitor.scala 107:30:freechips.rocketchip.system.DefaultRV32Config.fir@9795.8]
  wire  _T_330; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@9797.8]
  wire  _T_331; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@9798.8]
  wire  _T_336; // @[Monitor.scala 111:25:freechips.rocketchip.system.DefaultRV32Config.fir@9812.6]
  wire  _T_371; // @[Parameters.scala 552:42:freechips.rocketchip.system.DefaultRV32Config.fir@9848.8]
  wire  _T_372; // @[Parameters.scala 552:42:freechips.rocketchip.system.DefaultRV32Config.fir@9849.8]
  wire  _T_373; // @[Parameters.scala 552:42:freechips.rocketchip.system.DefaultRV32Config.fir@9850.8]
  wire  _T_374; // @[Parameters.scala 551:56:freechips.rocketchip.system.DefaultRV32Config.fir@9851.8]
  wire  _T_383; // @[Parameters.scala 93:42:freechips.rocketchip.system.DefaultRV32Config.fir@9860.8]
  wire  _T_391; // @[Parameters.scala 551:56:freechips.rocketchip.system.DefaultRV32Config.fir@9868.8]
  wire  _T_393; // @[Parameters.scala 553:30:freechips.rocketchip.system.DefaultRV32Config.fir@9870.8]
  wire  _T_395; // @[Parameters.scala 553:30:freechips.rocketchip.system.DefaultRV32Config.fir@9872.8]
  wire  _T_397; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@9874.8]
  wire  _T_398; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@9875.8]
  wire  _T_413; // @[Monitor.scala 119:25:freechips.rocketchip.system.DefaultRV32Config.fir@9911.6]
  wire [3:0] _T_486; // @[Monitor.scala 124:33:freechips.rocketchip.system.DefaultRV32Config.fir@10001.8]
  wire [3:0] _T_487; // @[Monitor.scala 124:31:freechips.rocketchip.system.DefaultRV32Config.fir@10002.8]
  wire  _T_488; // @[Monitor.scala 124:40:freechips.rocketchip.system.DefaultRV32Config.fir@10003.8]
  wire  _T_490; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@10005.8]
  wire  _T_491; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@10006.8]
  wire  _T_492; // @[Monitor.scala 127:25:freechips.rocketchip.system.DefaultRV32Config.fir@10012.6]
  wire  _T_494; // @[Parameters.scala 93:42:freechips.rocketchip.system.DefaultRV32Config.fir@10015.8]
  wire  _T_518; // @[Parameters.scala 552:42:freechips.rocketchip.system.DefaultRV32Config.fir@10039.8]
  wire  _T_519; // @[Parameters.scala 552:42:freechips.rocketchip.system.DefaultRV32Config.fir@10040.8]
  wire  _T_520; // @[Parameters.scala 551:56:freechips.rocketchip.system.DefaultRV32Config.fir@10041.8]
  wire  _T_543; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@10064.8]
  wire  _T_544; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@10065.8]
  wire  _T_551; // @[Bundles.scala 140:33:freechips.rocketchip.system.DefaultRV32Config.fir@10084.8]
  wire  _T_553; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@10086.8]
  wire  _T_554; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@10087.8]
  wire  _T_559; // @[Monitor.scala 135:25:freechips.rocketchip.system.DefaultRV32Config.fir@10101.6]
  wire  _T_618; // @[Bundles.scala 147:30:freechips.rocketchip.system.DefaultRV32Config.fir@10173.8]
  wire  _T_620; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@10175.8]
  wire  _T_621; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@10176.8]
  wire  _T_626; // @[Monitor.scala 143:25:freechips.rocketchip.system.DefaultRV32Config.fir@10190.6]
  wire  _T_677; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@10242.8]
  wire  _T_678; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@10243.8]
  wire  _T_685; // @[Bundles.scala 160:28:freechips.rocketchip.system.DefaultRV32Config.fir@10262.8]
  wire  _T_687; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@10264.8]
  wire  _T_688; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@10265.8]
  wire  _T_697; // @[Bundles.scala 44:24:freechips.rocketchip.system.DefaultRV32Config.fir@10289.6]
  wire  _T_699; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@10291.6]
  wire  _T_700; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@10292.6]
  wire  _T_701; // @[Parameters.scala 47:9:freechips.rocketchip.system.DefaultRV32Config.fir@10297.6]
  wire  _T_702; // @[Parameters.scala 47:9:freechips.rocketchip.system.DefaultRV32Config.fir@10298.6]
  wire  _T_703; // @[Parameters.scala 47:9:freechips.rocketchip.system.DefaultRV32Config.fir@10299.6]
  wire  _T_705; // @[Parameters.scala 924:46:freechips.rocketchip.system.DefaultRV32Config.fir@10305.6]
  wire  _T_706; // @[Parameters.scala 924:46:freechips.rocketchip.system.DefaultRV32Config.fir@10306.6]
  wire  _T_708; // @[Monitor.scala 307:25:freechips.rocketchip.system.DefaultRV32Config.fir@10308.6]
  wire  _T_710; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@10311.8]
  wire  _T_711; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@10312.8]
  wire  _T_712; // @[Monitor.scala 309:27:freechips.rocketchip.system.DefaultRV32Config.fir@10317.8]
  wire  _T_714; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@10319.8]
  wire  _T_715; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@10320.8]
  wire  _T_716; // @[Monitor.scala 310:28:freechips.rocketchip.system.DefaultRV32Config.fir@10325.8]
  wire  _T_718; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@10327.8]
  wire  _T_719; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@10328.8]
  wire  _T_720; // @[Monitor.scala 311:15:freechips.rocketchip.system.DefaultRV32Config.fir@10333.8]
  wire  _T_722; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@10335.8]
  wire  _T_723; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@10336.8]
  wire  _T_724; // @[Monitor.scala 312:15:freechips.rocketchip.system.DefaultRV32Config.fir@10341.8]
  wire  _T_726; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@10343.8]
  wire  _T_727; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@10344.8]
  wire  _T_728; // @[Monitor.scala 315:25:freechips.rocketchip.system.DefaultRV32Config.fir@10350.6]
  wire  _T_739; // @[Bundles.scala 104:26:freechips.rocketchip.system.DefaultRV32Config.fir@10374.8]
  wire  _T_741; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@10376.8]
  wire  _T_742; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@10377.8]
  wire  _T_743; // @[Monitor.scala 320:28:freechips.rocketchip.system.DefaultRV32Config.fir@10382.8]
  wire  _T_745; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@10384.8]
  wire  _T_746; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@10385.8]
  wire  _T_756; // @[Monitor.scala 325:25:freechips.rocketchip.system.DefaultRV32Config.fir@10408.6]
  wire  _T_776; // @[Monitor.scala 331:30:freechips.rocketchip.system.DefaultRV32Config.fir@10449.8]
  wire  _T_778; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@10451.8]
  wire  _T_779; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@10452.8]
  wire  _T_785; // @[Monitor.scala 335:25:freechips.rocketchip.system.DefaultRV32Config.fir@10467.6]
  wire  _T_802; // @[Monitor.scala 343:25:freechips.rocketchip.system.DefaultRV32Config.fir@10502.6]
  wire  _T_820; // @[Monitor.scala 351:25:freechips.rocketchip.system.DefaultRV32Config.fir@10538.6]
  wire [32:0] _T_844; // @[Parameters.scala 137:49:freechips.rocketchip.system.DefaultRV32Config.fir@10586.6]
  wire [31:0] _T_870; // @[Parameters.scala 137:31:freechips.rocketchip.system.DefaultRV32Config.fir@10616.6]
  wire [32:0] _T_871; // @[Parameters.scala 137:49:freechips.rocketchip.system.DefaultRV32Config.fir@10617.6]
  wire [32:0] _T_873; // @[Parameters.scala 137:52:freechips.rocketchip.system.DefaultRV32Config.fir@10619.6]
  wire  _T_874; // @[Parameters.scala 137:67:freechips.rocketchip.system.DefaultRV32Config.fir@10620.6]
  wire [31:0] _T_875; // @[Parameters.scala 137:31:freechips.rocketchip.system.DefaultRV32Config.fir@10621.6]
  wire [32:0] _T_876; // @[Parameters.scala 137:49:freechips.rocketchip.system.DefaultRV32Config.fir@10622.6]
  wire [32:0] _T_878; // @[Parameters.scala 137:52:freechips.rocketchip.system.DefaultRV32Config.fir@10624.6]
  wire  _T_879; // @[Parameters.scala 137:67:freechips.rocketchip.system.DefaultRV32Config.fir@10625.6]
  wire [31:0] _T_880; // @[Parameters.scala 137:31:freechips.rocketchip.system.DefaultRV32Config.fir@10626.6]
  wire [32:0] _T_881; // @[Parameters.scala 137:49:freechips.rocketchip.system.DefaultRV32Config.fir@10627.6]
  wire [32:0] _T_883; // @[Parameters.scala 137:52:freechips.rocketchip.system.DefaultRV32Config.fir@10629.6]
  wire  _T_884; // @[Parameters.scala 137:67:freechips.rocketchip.system.DefaultRV32Config.fir@10630.6]
  wire [32:0] _T_888; // @[Parameters.scala 137:52:freechips.rocketchip.system.DefaultRV32Config.fir@10634.6]
  wire  _T_889; // @[Parameters.scala 137:67:freechips.rocketchip.system.DefaultRV32Config.fir@10635.6]
  wire [31:0] _T_890; // @[Parameters.scala 137:31:freechips.rocketchip.system.DefaultRV32Config.fir@10636.6]
  wire [32:0] _T_891; // @[Parameters.scala 137:49:freechips.rocketchip.system.DefaultRV32Config.fir@10637.6]
  wire [32:0] _T_893; // @[Parameters.scala 137:52:freechips.rocketchip.system.DefaultRV32Config.fir@10639.6]
  wire  _T_894; // @[Parameters.scala 137:67:freechips.rocketchip.system.DefaultRV32Config.fir@10640.6]
  wire [31:0] _T_895; // @[Parameters.scala 137:31:freechips.rocketchip.system.DefaultRV32Config.fir@10641.6]
  wire [32:0] _T_896; // @[Parameters.scala 137:49:freechips.rocketchip.system.DefaultRV32Config.fir@10642.6]
  wire [32:0] _T_898; // @[Parameters.scala 137:52:freechips.rocketchip.system.DefaultRV32Config.fir@10644.6]
  wire  _T_899; // @[Parameters.scala 137:67:freechips.rocketchip.system.DefaultRV32Config.fir@10645.6]
  wire [31:0] _T_900; // @[Parameters.scala 137:31:freechips.rocketchip.system.DefaultRV32Config.fir@10646.6]
  wire [32:0] _T_901; // @[Parameters.scala 137:49:freechips.rocketchip.system.DefaultRV32Config.fir@10647.6]
  wire [32:0] _T_903; // @[Parameters.scala 137:52:freechips.rocketchip.system.DefaultRV32Config.fir@10649.6]
  wire  _T_904; // @[Parameters.scala 137:67:freechips.rocketchip.system.DefaultRV32Config.fir@10650.6]
  wire  _T_906; // @[Parameters.scala 535:64:freechips.rocketchip.system.DefaultRV32Config.fir@10660.6]
  wire  _T_907; // @[Parameters.scala 535:64:freechips.rocketchip.system.DefaultRV32Config.fir@10661.6]
  wire  _T_908; // @[Parameters.scala 535:64:freechips.rocketchip.system.DefaultRV32Config.fir@10662.6]
  wire  _T_909; // @[Parameters.scala 535:64:freechips.rocketchip.system.DefaultRV32Config.fir@10663.6]
  wire  _T_910; // @[Parameters.scala 535:64:freechips.rocketchip.system.DefaultRV32Config.fir@10664.6]
  wire  _T_911; // @[Parameters.scala 535:64:freechips.rocketchip.system.DefaultRV32Config.fir@10665.6]
  wire [31:0] _T_916; // @[Edges.scala 22:16:freechips.rocketchip.system.DefaultRV32Config.fir@10670.6]
  wire  _T_917; // @[Edges.scala 22:24:freechips.rocketchip.system.DefaultRV32Config.fir@10671.6]
  wire  _T_978; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@10747.8]
  wire  _T_979; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@10748.8]
  wire  _T_984; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@10761.8]
  wire  _T_985; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@10762.8]
  wire  _T_986; // @[Bundles.scala 104:26:freechips.rocketchip.system.DefaultRV32Config.fir@10767.8]
  wire  _T_988; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@10769.8]
  wire  _T_989; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@10770.8]
  wire  _T_1134; // @[Parameters.scala 47:9:freechips.rocketchip.system.DefaultRV32Config.fir@11094.6]
  wire  _T_1135; // @[Parameters.scala 47:9:freechips.rocketchip.system.DefaultRV32Config.fir@11095.6]
  wire  _T_1136; // @[Parameters.scala 47:9:freechips.rocketchip.system.DefaultRV32Config.fir@11096.6]
  wire  _T_1138; // @[Parameters.scala 924:46:freechips.rocketchip.system.DefaultRV32Config.fir@11102.6]
  wire  _T_1139; // @[Parameters.scala 924:46:freechips.rocketchip.system.DefaultRV32Config.fir@11103.6]
  wire [26:0] _T_1141; // @[package.scala 207:77:freechips.rocketchip.system.DefaultRV32Config.fir@11105.6]
  wire [11:0] _T_1143; // @[package.scala 207:46:freechips.rocketchip.system.DefaultRV32Config.fir@11107.6]
  wire [31:0] _GEN_72; // @[Edges.scala 22:16:freechips.rocketchip.system.DefaultRV32Config.fir@11108.6]
  wire [31:0] _T_1144; // @[Edges.scala 22:16:freechips.rocketchip.system.DefaultRV32Config.fir@11108.6]
  wire  _T_1145; // @[Edges.scala 22:24:freechips.rocketchip.system.DefaultRV32Config.fir@11109.6]
  wire [31:0] _T_1146; // @[Parameters.scala 137:31:freechips.rocketchip.system.DefaultRV32Config.fir@11110.6]
  wire [32:0] _T_1147; // @[Parameters.scala 137:49:freechips.rocketchip.system.DefaultRV32Config.fir@11111.6]
  wire [32:0] _T_1149; // @[Parameters.scala 137:52:freechips.rocketchip.system.DefaultRV32Config.fir@11113.6]
  wire  _T_1150; // @[Parameters.scala 137:67:freechips.rocketchip.system.DefaultRV32Config.fir@11114.6]
  wire [31:0] _T_1151; // @[Parameters.scala 137:31:freechips.rocketchip.system.DefaultRV32Config.fir@11115.6]
  wire [32:0] _T_1152; // @[Parameters.scala 137:49:freechips.rocketchip.system.DefaultRV32Config.fir@11116.6]
  wire [32:0] _T_1154; // @[Parameters.scala 137:52:freechips.rocketchip.system.DefaultRV32Config.fir@11118.6]
  wire  _T_1155; // @[Parameters.scala 137:67:freechips.rocketchip.system.DefaultRV32Config.fir@11119.6]
  wire [31:0] _T_1156; // @[Parameters.scala 137:31:freechips.rocketchip.system.DefaultRV32Config.fir@11120.6]
  wire [32:0] _T_1157; // @[Parameters.scala 137:49:freechips.rocketchip.system.DefaultRV32Config.fir@11121.6]
  wire [32:0] _T_1159; // @[Parameters.scala 137:52:freechips.rocketchip.system.DefaultRV32Config.fir@11123.6]
  wire  _T_1160; // @[Parameters.scala 137:67:freechips.rocketchip.system.DefaultRV32Config.fir@11124.6]
  wire [32:0] _T_1162; // @[Parameters.scala 137:49:freechips.rocketchip.system.DefaultRV32Config.fir@11126.6]
  wire [32:0] _T_1164; // @[Parameters.scala 137:52:freechips.rocketchip.system.DefaultRV32Config.fir@11128.6]
  wire  _T_1165; // @[Parameters.scala 137:67:freechips.rocketchip.system.DefaultRV32Config.fir@11129.6]
  wire [31:0] _T_1166; // @[Parameters.scala 137:31:freechips.rocketchip.system.DefaultRV32Config.fir@11130.6]
  wire [32:0] _T_1167; // @[Parameters.scala 137:49:freechips.rocketchip.system.DefaultRV32Config.fir@11131.6]
  wire [32:0] _T_1169; // @[Parameters.scala 137:52:freechips.rocketchip.system.DefaultRV32Config.fir@11133.6]
  wire  _T_1170; // @[Parameters.scala 137:67:freechips.rocketchip.system.DefaultRV32Config.fir@11134.6]
  wire [31:0] _T_1171; // @[Parameters.scala 137:31:freechips.rocketchip.system.DefaultRV32Config.fir@11135.6]
  wire [32:0] _T_1172; // @[Parameters.scala 137:49:freechips.rocketchip.system.DefaultRV32Config.fir@11136.6]
  wire [32:0] _T_1174; // @[Parameters.scala 137:52:freechips.rocketchip.system.DefaultRV32Config.fir@11138.6]
  wire  _T_1175; // @[Parameters.scala 137:67:freechips.rocketchip.system.DefaultRV32Config.fir@11139.6]
  wire [31:0] _T_1176; // @[Parameters.scala 137:31:freechips.rocketchip.system.DefaultRV32Config.fir@11140.6]
  wire [32:0] _T_1177; // @[Parameters.scala 137:49:freechips.rocketchip.system.DefaultRV32Config.fir@11141.6]
  wire [32:0] _T_1179; // @[Parameters.scala 137:52:freechips.rocketchip.system.DefaultRV32Config.fir@11143.6]
  wire  _T_1180; // @[Parameters.scala 137:67:freechips.rocketchip.system.DefaultRV32Config.fir@11144.6]
  wire  _T_1182; // @[Parameters.scala 535:64:freechips.rocketchip.system.DefaultRV32Config.fir@11154.6]
  wire  _T_1183; // @[Parameters.scala 535:64:freechips.rocketchip.system.DefaultRV32Config.fir@11155.6]
  wire  _T_1184; // @[Parameters.scala 535:64:freechips.rocketchip.system.DefaultRV32Config.fir@11156.6]
  wire  _T_1185; // @[Parameters.scala 535:64:freechips.rocketchip.system.DefaultRV32Config.fir@11157.6]
  wire  _T_1186; // @[Parameters.scala 535:64:freechips.rocketchip.system.DefaultRV32Config.fir@11158.6]
  wire  _T_1187; // @[Parameters.scala 535:64:freechips.rocketchip.system.DefaultRV32Config.fir@11159.6]
  wire  _T_1217; // @[Monitor.scala 239:25:freechips.rocketchip.system.DefaultRV32Config.fir@11193.6]
  wire  _T_1219; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@11196.8]
  wire  _T_1220; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@11197.8]
  wire  _T_1222; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@11203.8]
  wire  _T_1223; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@11204.8]
  wire  _T_1224; // @[Monitor.scala 242:30:freechips.rocketchip.system.DefaultRV32Config.fir@11209.8]
  wire  _T_1226; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@11211.8]
  wire  _T_1227; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@11212.8]
  wire  _T_1229; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@11218.8]
  wire  _T_1230; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@11219.8]
  wire  _T_1231; // @[Bundles.scala 122:29:freechips.rocketchip.system.DefaultRV32Config.fir@11224.8]
  wire  _T_1233; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@11226.8]
  wire  _T_1234; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@11227.8]
  wire  _T_1235; // @[Monitor.scala 245:18:freechips.rocketchip.system.DefaultRV32Config.fir@11232.8]
  wire  _T_1237; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@11234.8]
  wire  _T_1238; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@11235.8]
  wire  _T_1239; // @[Monitor.scala 248:25:freechips.rocketchip.system.DefaultRV32Config.fir@11241.6]
  wire  _T_1257; // @[Monitor.scala 256:25:freechips.rocketchip.system.DefaultRV32Config.fir@11281.6]
  wire  _T_1296; // @[Parameters.scala 93:42:freechips.rocketchip.system.DefaultRV32Config.fir@11321.8]
  wire  _T_1304; // @[Parameters.scala 551:56:freechips.rocketchip.system.DefaultRV32Config.fir@11329.8]
  wire  _T_1308; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@11333.8]
  wire  _T_1309; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@11334.8]
  wire  _T_1314; // @[Parameters.scala 92:48:freechips.rocketchip.system.DefaultRV32Config.fir@11347.8]
  wire  _T_1315; // @[Mux.scala 27:72:freechips.rocketchip.system.DefaultRV32Config.fir@11348.8]
  wire  _T_1322; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@11356.8]
  wire  _T_1323; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@11357.8]
  wire  _T_1334; // @[Bundles.scala 116:29:freechips.rocketchip.system.DefaultRV32Config.fir@11384.8]
  wire  _T_1336; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@11386.8]
  wire  _T_1337; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@11387.8]
  wire  _T_1342; // @[Monitor.scala 266:25:freechips.rocketchip.system.DefaultRV32Config.fir@11401.6]
  wire  _T_1423; // @[Monitor.scala 275:25:freechips.rocketchip.system.DefaultRV32Config.fir@11513.6]
  wire  _T_1433; // @[Monitor.scala 279:31:freechips.rocketchip.system.DefaultRV32Config.fir@11536.8]
  wire  _T_1435; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@11538.8]
  wire  _T_1436; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@11539.8]
  wire  _T_1441; // @[Monitor.scala 283:25:freechips.rocketchip.system.DefaultRV32Config.fir@11553.6]
  wire  _T_1455; // @[Monitor.scala 290:25:freechips.rocketchip.system.DefaultRV32Config.fir@11585.6]
  wire  _T_1477; // @[Decoupled.scala 40:37:freechips.rocketchip.system.DefaultRV32Config.fir@11636.4]
  wire  _T_1484; // @[Edges.scala 93:28:freechips.rocketchip.system.DefaultRV32Config.fir@11643.4]
  reg [9:0] _T_1486; // @[Edges.scala 230:27:freechips.rocketchip.system.DefaultRV32Config.fir@11645.4]
  wire [9:0] _T_1488; // @[Edges.scala 231:28:freechips.rocketchip.system.DefaultRV32Config.fir@11647.4]
  wire  _T_1489; // @[Edges.scala 232:25:freechips.rocketchip.system.DefaultRV32Config.fir@11648.4]
  reg [2:0] _T_1497; // @[Monitor.scala 381:22:freechips.rocketchip.system.DefaultRV32Config.fir@11659.4]
  reg [2:0] _T_1498; // @[Monitor.scala 382:22:freechips.rocketchip.system.DefaultRV32Config.fir@11660.4]
  reg [3:0] _T_1499; // @[Monitor.scala 383:22:freechips.rocketchip.system.DefaultRV32Config.fir@11661.4]
  reg [1:0] _T_1500; // @[Monitor.scala 384:22:freechips.rocketchip.system.DefaultRV32Config.fir@11662.4]
  reg [31:0] _T_1501; // @[Monitor.scala 385:22:freechips.rocketchip.system.DefaultRV32Config.fir@11663.4]
  wire  _T_1502; // @[Monitor.scala 386:22:freechips.rocketchip.system.DefaultRV32Config.fir@11664.4]
  wire  _T_1503; // @[Monitor.scala 386:19:freechips.rocketchip.system.DefaultRV32Config.fir@11665.4]
  wire  _T_1504; // @[Monitor.scala 387:32:freechips.rocketchip.system.DefaultRV32Config.fir@11667.6]
  wire  _T_1506; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@11669.6]
  wire  _T_1507; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@11670.6]
  wire  _T_1508; // @[Monitor.scala 388:32:freechips.rocketchip.system.DefaultRV32Config.fir@11675.6]
  wire  _T_1510; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@11677.6]
  wire  _T_1511; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@11678.6]
  wire  _T_1512; // @[Monitor.scala 389:32:freechips.rocketchip.system.DefaultRV32Config.fir@11683.6]
  wire  _T_1514; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@11685.6]
  wire  _T_1515; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@11686.6]
  wire  _T_1516; // @[Monitor.scala 390:32:freechips.rocketchip.system.DefaultRV32Config.fir@11691.6]
  wire  _T_1518; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@11693.6]
  wire  _T_1519; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@11694.6]
  wire  _T_1520; // @[Monitor.scala 391:32:freechips.rocketchip.system.DefaultRV32Config.fir@11699.6]
  wire  _T_1522; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@11701.6]
  wire  _T_1523; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@11702.6]
  wire  _T_1525; // @[Monitor.scala 393:20:freechips.rocketchip.system.DefaultRV32Config.fir@11709.4]
  wire  _T_1526; // @[Decoupled.scala 40:37:freechips.rocketchip.system.DefaultRV32Config.fir@11717.4]
  wire [26:0] _T_1528; // @[package.scala 207:77:freechips.rocketchip.system.DefaultRV32Config.fir@11719.4]
  wire [11:0] _T_1530; // @[package.scala 207:46:freechips.rocketchip.system.DefaultRV32Config.fir@11721.4]
  reg [9:0] _T_1534; // @[Edges.scala 230:27:freechips.rocketchip.system.DefaultRV32Config.fir@11725.4]
  wire [9:0] _T_1536; // @[Edges.scala 231:28:freechips.rocketchip.system.DefaultRV32Config.fir@11727.4]
  wire  _T_1537; // @[Edges.scala 232:25:freechips.rocketchip.system.DefaultRV32Config.fir@11728.4]
  reg [2:0] _T_1545; // @[Monitor.scala 532:22:freechips.rocketchip.system.DefaultRV32Config.fir@11739.4]
  reg [1:0] _T_1546; // @[Monitor.scala 533:22:freechips.rocketchip.system.DefaultRV32Config.fir@11740.4]
  reg [3:0] _T_1547; // @[Monitor.scala 534:22:freechips.rocketchip.system.DefaultRV32Config.fir@11741.4]
  reg [1:0] _T_1548; // @[Monitor.scala 535:22:freechips.rocketchip.system.DefaultRV32Config.fir@11742.4]
  reg [1:0] _T_1549; // @[Monitor.scala 536:22:freechips.rocketchip.system.DefaultRV32Config.fir@11743.4]
  reg  _T_1550; // @[Monitor.scala 537:22:freechips.rocketchip.system.DefaultRV32Config.fir@11744.4]
  wire  _T_1551; // @[Monitor.scala 538:22:freechips.rocketchip.system.DefaultRV32Config.fir@11745.4]
  wire  _T_1552; // @[Monitor.scala 538:19:freechips.rocketchip.system.DefaultRV32Config.fir@11746.4]
  wire  _T_1553; // @[Monitor.scala 539:29:freechips.rocketchip.system.DefaultRV32Config.fir@11748.6]
  wire  _T_1555; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@11750.6]
  wire  _T_1556; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@11751.6]
  wire  _T_1557; // @[Monitor.scala 540:29:freechips.rocketchip.system.DefaultRV32Config.fir@11756.6]
  wire  _T_1559; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@11758.6]
  wire  _T_1560; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@11759.6]
  wire  _T_1561; // @[Monitor.scala 541:29:freechips.rocketchip.system.DefaultRV32Config.fir@11764.6]
  wire  _T_1563; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@11766.6]
  wire  _T_1564; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@11767.6]
  wire  _T_1565; // @[Monitor.scala 542:29:freechips.rocketchip.system.DefaultRV32Config.fir@11772.6]
  wire  _T_1567; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@11774.6]
  wire  _T_1568; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@11775.6]
  wire  _T_1569; // @[Monitor.scala 543:29:freechips.rocketchip.system.DefaultRV32Config.fir@11780.6]
  wire  _T_1571; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@11782.6]
  wire  _T_1572; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@11783.6]
  wire  _T_1573; // @[Monitor.scala 544:29:freechips.rocketchip.system.DefaultRV32Config.fir@11788.6]
  wire  _T_1575; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@11790.6]
  wire  _T_1576; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@11791.6]
  wire  _T_1578; // @[Monitor.scala 546:20:freechips.rocketchip.system.DefaultRV32Config.fir@11798.4]
  wire  _T_1579; // @[Decoupled.scala 40:37:freechips.rocketchip.system.DefaultRV32Config.fir@11807.4]
  reg [9:0] _T_1588; // @[Edges.scala 230:27:freechips.rocketchip.system.DefaultRV32Config.fir@11816.4]
  wire [9:0] _T_1590; // @[Edges.scala 231:28:freechips.rocketchip.system.DefaultRV32Config.fir@11818.4]
  wire  _T_1591; // @[Edges.scala 232:25:freechips.rocketchip.system.DefaultRV32Config.fir@11819.4]
  reg [1:0] _T_1600; // @[Monitor.scala 405:22:freechips.rocketchip.system.DefaultRV32Config.fir@11831.4]
  reg [31:0] _T_1603; // @[Monitor.scala 408:22:freechips.rocketchip.system.DefaultRV32Config.fir@11834.4]
  wire  _T_1604; // @[Monitor.scala 409:22:freechips.rocketchip.system.DefaultRV32Config.fir@11835.4]
  wire  _T_1605; // @[Monitor.scala 409:19:freechips.rocketchip.system.DefaultRV32Config.fir@11836.4]
  wire  _T_1610; // @[Monitor.scala 411:32:freechips.rocketchip.system.DefaultRV32Config.fir@11846.6]
  wire  _T_1612; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@11848.6]
  wire  _T_1613; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@11849.6]
  wire  _T_1622; // @[Monitor.scala 414:32:freechips.rocketchip.system.DefaultRV32Config.fir@11870.6]
  wire  _T_1624; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@11872.6]
  wire  _T_1625; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@11873.6]
  wire  _T_1627; // @[Monitor.scala 416:20:freechips.rocketchip.system.DefaultRV32Config.fir@11880.4]
  wire  _T_1628; // @[Decoupled.scala 40:37:freechips.rocketchip.system.DefaultRV32Config.fir@11888.4]
  reg [9:0] _T_1636; // @[Edges.scala 230:27:freechips.rocketchip.system.DefaultRV32Config.fir@11896.4]
  wire [9:0] _T_1638; // @[Edges.scala 231:28:freechips.rocketchip.system.DefaultRV32Config.fir@11898.4]
  wire  _T_1639; // @[Edges.scala 232:25:freechips.rocketchip.system.DefaultRV32Config.fir@11899.4]
  reg [2:0] _T_1647; // @[Monitor.scala 509:22:freechips.rocketchip.system.DefaultRV32Config.fir@11910.4]
  reg [2:0] _T_1648; // @[Monitor.scala 510:22:freechips.rocketchip.system.DefaultRV32Config.fir@11911.4]
  reg [3:0] _T_1649; // @[Monitor.scala 511:22:freechips.rocketchip.system.DefaultRV32Config.fir@11912.4]
  reg [1:0] _T_1650; // @[Monitor.scala 512:22:freechips.rocketchip.system.DefaultRV32Config.fir@11913.4]
  reg [31:0] _T_1651; // @[Monitor.scala 513:22:freechips.rocketchip.system.DefaultRV32Config.fir@11914.4]
  wire  _T_1652; // @[Monitor.scala 514:22:freechips.rocketchip.system.DefaultRV32Config.fir@11915.4]
  wire  _T_1653; // @[Monitor.scala 514:19:freechips.rocketchip.system.DefaultRV32Config.fir@11916.4]
  wire  _T_1654; // @[Monitor.scala 515:32:freechips.rocketchip.system.DefaultRV32Config.fir@11918.6]
  wire  _T_1656; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@11920.6]
  wire  _T_1657; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@11921.6]
  wire  _T_1658; // @[Monitor.scala 516:32:freechips.rocketchip.system.DefaultRV32Config.fir@11926.6]
  wire  _T_1660; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@11928.6]
  wire  _T_1661; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@11929.6]
  wire  _T_1662; // @[Monitor.scala 517:32:freechips.rocketchip.system.DefaultRV32Config.fir@11934.6]
  wire  _T_1664; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@11936.6]
  wire  _T_1665; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@11937.6]
  wire  _T_1666; // @[Monitor.scala 518:32:freechips.rocketchip.system.DefaultRV32Config.fir@11942.6]
  wire  _T_1668; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@11944.6]
  wire  _T_1669; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@11945.6]
  wire  _T_1670; // @[Monitor.scala 519:32:freechips.rocketchip.system.DefaultRV32Config.fir@11950.6]
  wire  _T_1672; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@11952.6]
  wire  _T_1673; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@11953.6]
  wire  _T_1675; // @[Monitor.scala 521:20:freechips.rocketchip.system.DefaultRV32Config.fir@11960.4]
  reg [2:0] inflight; // @[Monitor.scala 608:27:freechips.rocketchip.system.DefaultRV32Config.fir@11968.4]
  reg [11:0] inflight_opcodes; // @[Monitor.scala 610:35:freechips.rocketchip.system.DefaultRV32Config.fir@11969.4]
  reg [23:0] inflight_sizes; // @[Monitor.scala 612:33:freechips.rocketchip.system.DefaultRV32Config.fir@11970.4]
  reg [9:0] _T_1685; // @[Edges.scala 230:27:freechips.rocketchip.system.DefaultRV32Config.fir@11980.4]
  wire [9:0] _T_1687; // @[Edges.scala 231:28:freechips.rocketchip.system.DefaultRV32Config.fir@11982.4]
  wire  a_first; // @[Edges.scala 232:25:freechips.rocketchip.system.DefaultRV32Config.fir@11983.4]
  reg [9:0] _T_1703; // @[Edges.scala 230:27:freechips.rocketchip.system.DefaultRV32Config.fir@12002.4]
  wire [9:0] _T_1705; // @[Edges.scala 231:28:freechips.rocketchip.system.DefaultRV32Config.fir@12004.4]
  wire  d_first; // @[Edges.scala 232:25:freechips.rocketchip.system.DefaultRV32Config.fir@12005.4]
  wire [3:0] _GEN_73; // @[Monitor.scala 629:69:freechips.rocketchip.system.DefaultRV32Config.fir@12024.4]
  wire [4:0] _T_1713; // @[Monitor.scala 629:69:freechips.rocketchip.system.DefaultRV32Config.fir@12024.4]
  wire [11:0] _T_1714; // @[Monitor.scala 629:44:freechips.rocketchip.system.DefaultRV32Config.fir@12025.4]
  wire [15:0] _T_1718; // @[Monitor.scala 606:57:freechips.rocketchip.system.DefaultRV32Config.fir@12029.4]
  wire [15:0] _GEN_74; // @[Monitor.scala 629:97:freechips.rocketchip.system.DefaultRV32Config.fir@12030.4]
  wire [15:0] _T_1719; // @[Monitor.scala 629:97:freechips.rocketchip.system.DefaultRV32Config.fir@12030.4]
  wire [15:0] _T_1720; // @[Monitor.scala 629:152:freechips.rocketchip.system.DefaultRV32Config.fir@12031.4]
  wire [4:0] _T_1721; // @[Monitor.scala 633:65:freechips.rocketchip.system.DefaultRV32Config.fir@12035.4]
  wire [23:0] _T_1722; // @[Monitor.scala 633:40:freechips.rocketchip.system.DefaultRV32Config.fir@12036.4]
  wire [15:0] _T_1726; // @[Monitor.scala 606:57:freechips.rocketchip.system.DefaultRV32Config.fir@12040.4]
  wire [23:0] _GEN_76; // @[Monitor.scala 633:91:freechips.rocketchip.system.DefaultRV32Config.fir@12041.4]
  wire [23:0] _T_1727; // @[Monitor.scala 633:91:freechips.rocketchip.system.DefaultRV32Config.fir@12041.4]
  wire [23:0] _T_1728; // @[Monitor.scala 633:144:freechips.rocketchip.system.DefaultRV32Config.fir@12042.4]
  wire  _T_1732; // @[Monitor.scala 643:27:freechips.rocketchip.system.DefaultRV32Config.fir@12067.4]
  wire [3:0] _T_1734; // @[OneHot.scala 58:35:freechips.rocketchip.system.DefaultRV32Config.fir@12070.6]
  wire [3:0] _T_1735; // @[Monitor.scala 645:53:freechips.rocketchip.system.DefaultRV32Config.fir@12072.6]
  wire [3:0] _T_1736; // @[Monitor.scala 645:61:freechips.rocketchip.system.DefaultRV32Config.fir@12073.6]
  wire [4:0] _T_1737; // @[Monitor.scala 646:49:freechips.rocketchip.system.DefaultRV32Config.fir@12075.6]
  wire [4:0] _T_1738; // @[Monitor.scala 646:57:freechips.rocketchip.system.DefaultRV32Config.fir@12076.6]
  wire [3:0] _GEN_78; // @[Monitor.scala 647:72:freechips.rocketchip.system.DefaultRV32Config.fir@12078.6]
  wire [4:0] _T_1739; // @[Monitor.scala 647:72:freechips.rocketchip.system.DefaultRV32Config.fir@12078.6]
  wire [3:0] a_opcodes_set_interm; // @[Monitor.scala 643:72:freechips.rocketchip.system.DefaultRV32Config.fir@12069.4]
  wire [34:0] _GEN_79; // @[Monitor.scala 647:47:freechips.rocketchip.system.DefaultRV32Config.fir@12079.6]
  wire [34:0] _T_1740; // @[Monitor.scala 647:47:freechips.rocketchip.system.DefaultRV32Config.fir@12079.6]
  wire [4:0] _T_1741; // @[Monitor.scala 648:68:freechips.rocketchip.system.DefaultRV32Config.fir@12081.6]
  wire [4:0] a_sizes_set_interm; // @[Monitor.scala 643:72:freechips.rocketchip.system.DefaultRV32Config.fir@12069.4]
  wire [35:0] _GEN_80; // @[Monitor.scala 648:43:freechips.rocketchip.system.DefaultRV32Config.fir@12082.6]
  wire [35:0] _T_1742; // @[Monitor.scala 648:43:freechips.rocketchip.system.DefaultRV32Config.fir@12082.6]
  wire [2:0] _T_1743; // @[Monitor.scala 649:26:freechips.rocketchip.system.DefaultRV32Config.fir@12084.6]
  wire  _T_1745; // @[Monitor.scala 649:17:freechips.rocketchip.system.DefaultRV32Config.fir@12086.6]
  wire  _T_1747; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@12088.6]
  wire  _T_1748; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@12089.6]
  wire [3:0] _GEN_27; // @[Monitor.scala 643:72:freechips.rocketchip.system.DefaultRV32Config.fir@12069.4]
  wire [34:0] _GEN_30; // @[Monitor.scala 643:72:freechips.rocketchip.system.DefaultRV32Config.fir@12069.4]
  wire [35:0] _GEN_31; // @[Monitor.scala 643:72:freechips.rocketchip.system.DefaultRV32Config.fir@12069.4]
  wire  _T_1751; // @[Monitor.scala 660:27:freechips.rocketchip.system.DefaultRV32Config.fir@12103.4]
  wire  _T_1753; // @[Monitor.scala 660:75:freechips.rocketchip.system.DefaultRV32Config.fir@12105.4]
  wire  _T_1754; // @[Monitor.scala 660:72:freechips.rocketchip.system.DefaultRV32Config.fir@12106.4]
  wire [3:0] _T_1755; // @[OneHot.scala 58:35:freechips.rocketchip.system.DefaultRV32Config.fir@12108.6]
  wire [46:0] _GEN_82; // @[Monitor.scala 662:76:freechips.rocketchip.system.DefaultRV32Config.fir@12115.6]
  wire [46:0] _T_1761; // @[Monitor.scala 662:76:freechips.rocketchip.system.DefaultRV32Config.fir@12115.6]
  wire [46:0] _GEN_83; // @[Monitor.scala 663:72:freechips.rocketchip.system.DefaultRV32Config.fir@12122.6]
  wire [46:0] _T_1767; // @[Monitor.scala 663:72:freechips.rocketchip.system.DefaultRV32Config.fir@12122.6]
  wire [3:0] _GEN_32; // @[Monitor.scala 660:91:freechips.rocketchip.system.DefaultRV32Config.fir@12107.4]
  wire [46:0] _GEN_33; // @[Monitor.scala 660:91:freechips.rocketchip.system.DefaultRV32Config.fir@12107.4]
  wire [46:0] _GEN_34; // @[Monitor.scala 660:91:freechips.rocketchip.system.DefaultRV32Config.fir@12107.4]
  wire  _T_1768; // @[Monitor.scala 665:26:freechips.rocketchip.system.DefaultRV32Config.fir@12125.4]
  wire  _T_1771; // @[Monitor.scala 665:71:freechips.rocketchip.system.DefaultRV32Config.fir@12128.4]
  wire [2:0] _T_1772; // @[Monitor.scala 666:25:freechips.rocketchip.system.DefaultRV32Config.fir@12130.6]
  wire  _T_1774; // @[Monitor.scala 666:93:freechips.rocketchip.system.DefaultRV32Config.fir@12132.6]
  wire  _T_1775; // @[Monitor.scala 666:68:freechips.rocketchip.system.DefaultRV32Config.fir@12133.6]
  wire  _T_1776; // @[Monitor.scala 666:142:freechips.rocketchip.system.DefaultRV32Config.fir@12134.6]
  wire  _T_1777; // @[Monitor.scala 666:119:freechips.rocketchip.system.DefaultRV32Config.fir@12135.6]
  wire  _T_1778; // @[Monitor.scala 666:166:freechips.rocketchip.system.DefaultRV32Config.fir@12136.6]
  wire  _T_1779; // @[Monitor.scala 666:49:freechips.rocketchip.system.DefaultRV32Config.fir@12137.6]
  wire  _T_1781; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@12139.6]
  wire  _T_1782; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@12140.6]
  wire [3:0] a_opcode_lookup; // @[:freechips.rocketchip.system.DefaultRV32Config.fir@12022.4 :freechips.rocketchip.system.DefaultRV32Config.fir@12023.4 Monitor.scala 629:21:freechips.rocketchip.system.DefaultRV32Config.fir@12032.4]
  wire [2:0] _GEN_37; // @[Monitor.scala 667:37:freechips.rocketchip.system.DefaultRV32Config.fir@12146.6]
  wire [2:0] _GEN_38; // @[Monitor.scala 667:37:freechips.rocketchip.system.DefaultRV32Config.fir@12146.6]
  wire [2:0] _GEN_39; // @[Monitor.scala 667:37:freechips.rocketchip.system.DefaultRV32Config.fir@12146.6]
  wire [2:0] _GEN_40; // @[Monitor.scala 667:37:freechips.rocketchip.system.DefaultRV32Config.fir@12146.6]
  wire [2:0] _GEN_41; // @[Monitor.scala 667:37:freechips.rocketchip.system.DefaultRV32Config.fir@12146.6]
  wire [2:0] _GEN_42; // @[Monitor.scala 667:37:freechips.rocketchip.system.DefaultRV32Config.fir@12146.6]
  wire  _T_1784; // @[Monitor.scala 667:37:freechips.rocketchip.system.DefaultRV32Config.fir@12146.6]
  wire [2:0] _GEN_49; // @[Monitor.scala 667:96:freechips.rocketchip.system.DefaultRV32Config.fir@12148.6]
  wire [2:0] _GEN_50; // @[Monitor.scala 667:96:freechips.rocketchip.system.DefaultRV32Config.fir@12148.6]
  wire  _T_1786; // @[Monitor.scala 667:96:freechips.rocketchip.system.DefaultRV32Config.fir@12148.6]
  wire  _T_1787; // @[Monitor.scala 667:71:freechips.rocketchip.system.DefaultRV32Config.fir@12149.6]
  wire [2:0] _GEN_53; // @[Monitor.scala 668:60:freechips.rocketchip.system.DefaultRV32Config.fir@12150.6]
  wire [2:0] _GEN_54; // @[Monitor.scala 668:60:freechips.rocketchip.system.DefaultRV32Config.fir@12150.6]
  wire [2:0] _GEN_55; // @[Monitor.scala 668:60:freechips.rocketchip.system.DefaultRV32Config.fir@12150.6]
  wire [2:0] _GEN_56; // @[Monitor.scala 668:60:freechips.rocketchip.system.DefaultRV32Config.fir@12150.6]
  wire [2:0] _GEN_57; // @[Monitor.scala 668:60:freechips.rocketchip.system.DefaultRV32Config.fir@12150.6]
  wire [2:0] _GEN_58; // @[Monitor.scala 668:60:freechips.rocketchip.system.DefaultRV32Config.fir@12150.6]
  wire  _T_1788; // @[Monitor.scala 668:60:freechips.rocketchip.system.DefaultRV32Config.fir@12150.6]
  wire [2:0] _GEN_65; // @[Monitor.scala 668:124:freechips.rocketchip.system.DefaultRV32Config.fir@12151.6]
  wire [2:0] _GEN_66; // @[Monitor.scala 668:124:freechips.rocketchip.system.DefaultRV32Config.fir@12151.6]
  wire  _T_1789; // @[Monitor.scala 668:124:freechips.rocketchip.system.DefaultRV32Config.fir@12151.6]
  wire  _T_1790; // @[Monitor.scala 668:99:freechips.rocketchip.system.DefaultRV32Config.fir@12152.6]
  wire  _T_1791; // @[Monitor.scala 668:34:freechips.rocketchip.system.DefaultRV32Config.fir@12153.6]
  wire  _T_1792; // @[Monitor.scala 668:15:freechips.rocketchip.system.DefaultRV32Config.fir@12154.6]
  wire  _T_1794; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@12156.6]
  wire  _T_1795; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@12157.6]
  wire [7:0] a_size_lookup; // @[:freechips.rocketchip.system.DefaultRV32Config.fir@12033.4 :freechips.rocketchip.system.DefaultRV32Config.fir@12034.4 Monitor.scala 633:19:freechips.rocketchip.system.DefaultRV32Config.fir@12043.4]
  wire [7:0] _GEN_84; // @[Monitor.scala 670:34:freechips.rocketchip.system.DefaultRV32Config.fir@12162.6]
  wire  _T_1796; // @[Monitor.scala 670:34:freechips.rocketchip.system.DefaultRV32Config.fir@12162.6]
  wire  _T_1798; // @[Monitor.scala 670:72:freechips.rocketchip.system.DefaultRV32Config.fir@12164.6]
  wire  _T_1799; // @[Monitor.scala 670:53:freechips.rocketchip.system.DefaultRV32Config.fir@12165.6]
  wire  _T_1801; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@12167.6]
  wire  _T_1802; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@12168.6]
  wire  _T_1804; // @[Monitor.scala 672:36:freechips.rocketchip.system.DefaultRV32Config.fir@12175.4]
  wire  _T_1805; // @[Monitor.scala 672:47:freechips.rocketchip.system.DefaultRV32Config.fir@12176.4]
  wire  _T_1807; // @[Monitor.scala 672:65:freechips.rocketchip.system.DefaultRV32Config.fir@12178.4]
  wire  _T_1809; // @[Monitor.scala 672:116:freechips.rocketchip.system.DefaultRV32Config.fir@12180.4]
  wire  _T_1810; // @[Monitor.scala 673:15:freechips.rocketchip.system.DefaultRV32Config.fir@12182.6]
  wire  _T_1811; // @[Monitor.scala 673:32:freechips.rocketchip.system.DefaultRV32Config.fir@12183.6]
  wire  _T_1813; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@12185.6]
  wire  _T_1814; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@12186.6]
  wire [2:0] a_set; // @[:freechips.rocketchip.system.DefaultRV32Config.fir@12016.4 :freechips.rocketchip.system.DefaultRV32Config.fir@12017.4 Monitor.scala 644:13:freechips.rocketchip.system.DefaultRV32Config.fir@12071.6]
  wire [2:0] d_clr; // @[:freechips.rocketchip.system.DefaultRV32Config.fir@12095.4 :freechips.rocketchip.system.DefaultRV32Config.fir@12096.4 Monitor.scala 661:13:freechips.rocketchip.system.DefaultRV32Config.fir@12109.6]
  wire  _T_1815; // @[Monitor.scala 677:20:freechips.rocketchip.system.DefaultRV32Config.fir@12192.4]
  wire  _T_1816; // @[Monitor.scala 677:40:freechips.rocketchip.system.DefaultRV32Config.fir@12193.4]
  wire  _T_1817; // @[Monitor.scala 677:33:freechips.rocketchip.system.DefaultRV32Config.fir@12194.4]
  wire  _T_1818; // @[Monitor.scala 677:30:freechips.rocketchip.system.DefaultRV32Config.fir@12195.4]
  wire  _T_1820; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@12197.4]
  wire  _T_1821; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@12198.4]
  wire [2:0] _T_1822; // @[Monitor.scala 680:27:freechips.rocketchip.system.DefaultRV32Config.fir@12203.4]
  wire [2:0] _T_1823; // @[Monitor.scala 680:38:freechips.rocketchip.system.DefaultRV32Config.fir@12204.4]
  wire [2:0] _T_1824; // @[Monitor.scala 680:36:freechips.rocketchip.system.DefaultRV32Config.fir@12205.4]
  wire [11:0] a_opcodes_set; // @[:freechips.rocketchip.system.DefaultRV32Config.fir@12018.4 :freechips.rocketchip.system.DefaultRV32Config.fir@12019.4 Monitor.scala 647:21:freechips.rocketchip.system.DefaultRV32Config.fir@12080.6]
  wire [11:0] _T_1825; // @[Monitor.scala 681:43:freechips.rocketchip.system.DefaultRV32Config.fir@12207.4]
  wire [11:0] d_opcodes_clr; // @[:freechips.rocketchip.system.DefaultRV32Config.fir@12097.4 :freechips.rocketchip.system.DefaultRV32Config.fir@12098.4 Monitor.scala 662:21:freechips.rocketchip.system.DefaultRV32Config.fir@12116.6]
  wire [11:0] _T_1826; // @[Monitor.scala 681:62:freechips.rocketchip.system.DefaultRV32Config.fir@12208.4]
  wire [11:0] _T_1827; // @[Monitor.scala 681:60:freechips.rocketchip.system.DefaultRV32Config.fir@12209.4]
  wire [23:0] a_sizes_set; // @[:freechips.rocketchip.system.DefaultRV32Config.fir@12020.4 :freechips.rocketchip.system.DefaultRV32Config.fir@12021.4 Monitor.scala 648:19:freechips.rocketchip.system.DefaultRV32Config.fir@12083.6]
  wire [23:0] _T_1828; // @[Monitor.scala 682:39:freechips.rocketchip.system.DefaultRV32Config.fir@12211.4]
  wire [23:0] d_sizes_clr; // @[:freechips.rocketchip.system.DefaultRV32Config.fir@12099.4 :freechips.rocketchip.system.DefaultRV32Config.fir@12100.4 Monitor.scala 663:19:freechips.rocketchip.system.DefaultRV32Config.fir@12123.6]
  wire [23:0] _T_1829; // @[Monitor.scala 682:56:freechips.rocketchip.system.DefaultRV32Config.fir@12212.4]
  wire [23:0] _T_1830; // @[Monitor.scala 682:54:freechips.rocketchip.system.DefaultRV32Config.fir@12213.4]
  reg [31:0] _T_1831; // @[Monitor.scala 684:27:freechips.rocketchip.system.DefaultRV32Config.fir@12215.4]
  wire  _T_1832; // @[Monitor.scala 687:26:freechips.rocketchip.system.DefaultRV32Config.fir@12218.4]
  wire  _T_1833; // @[Monitor.scala 687:16:freechips.rocketchip.system.DefaultRV32Config.fir@12219.4]
  wire  _T_1834; // @[Monitor.scala 687:39:freechips.rocketchip.system.DefaultRV32Config.fir@12220.4]
  wire  _T_1835; // @[Monitor.scala 687:30:freechips.rocketchip.system.DefaultRV32Config.fir@12221.4]
  wire  _T_1836; // @[Monitor.scala 687:59:freechips.rocketchip.system.DefaultRV32Config.fir@12222.4]
  wire  _T_1837; // @[Monitor.scala 687:47:freechips.rocketchip.system.DefaultRV32Config.fir@12223.4]
  wire  _T_1839; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@12225.4]
  wire  _T_1840; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@12226.4]
  wire [31:0] _T_1842; // @[Monitor.scala 689:26:freechips.rocketchip.system.DefaultRV32Config.fir@12232.4]
  wire  _T_1845; // @[Monitor.scala 690:27:freechips.rocketchip.system.DefaultRV32Config.fir@12236.4]
  reg [3:0] _T_1846; // @[Monitor.scala 694:27:freechips.rocketchip.system.DefaultRV32Config.fir@12240.4]
  reg [9:0] _T_1855; // @[Edges.scala 230:27:freechips.rocketchip.system.DefaultRV32Config.fir@12249.4]
  wire [9:0] _T_1857; // @[Edges.scala 231:28:freechips.rocketchip.system.DefaultRV32Config.fir@12251.4]
  wire  _T_1858; // @[Edges.scala 232:25:freechips.rocketchip.system.DefaultRV32Config.fir@12252.4]
  wire  _T_1868; // @[Monitor.scala 700:27:freechips.rocketchip.system.DefaultRV32Config.fir@12266.4]
  wire  _T_1871; // @[Edges.scala 72:43:freechips.rocketchip.system.DefaultRV32Config.fir@12269.4]
  wire  _T_1872; // @[Edges.scala 72:40:freechips.rocketchip.system.DefaultRV32Config.fir@12270.4]
  wire  _T_1873; // @[Monitor.scala 700:38:freechips.rocketchip.system.DefaultRV32Config.fir@12271.4]
  wire [3:0] _T_1874; // @[OneHot.scala 58:35:freechips.rocketchip.system.DefaultRV32Config.fir@12273.6]
  wire [3:0] _T_1875; // @[Monitor.scala 702:23:freechips.rocketchip.system.DefaultRV32Config.fir@12275.6]
  wire  _T_1877; // @[Monitor.scala 702:14:freechips.rocketchip.system.DefaultRV32Config.fir@12277.6]
  wire  _T_1879; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@12279.6]
  wire  _T_1880; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@12280.6]
  wire [3:0] _GEN_69; // @[Monitor.scala 700:72:freechips.rocketchip.system.DefaultRV32Config.fir@12272.4]
  wire [3:0] _T_1885; // @[OneHot.scala 58:35:freechips.rocketchip.system.DefaultRV32Config.fir@12292.6]
  wire [3:0] _T_1886; // @[Monitor.scala 708:24:freechips.rocketchip.system.DefaultRV32Config.fir@12294.6]
  wire [3:0] _T_1887; // @[Monitor.scala 708:35:freechips.rocketchip.system.DefaultRV32Config.fir@12295.6]
  wire  _T_1890; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@12298.6]
  wire  _T_1891; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@12299.6]
  wire [3:0] _GEN_70; // @[Monitor.scala 706:73:freechips.rocketchip.system.DefaultRV32Config.fir@12291.4]
  wire [3:0] _T_1892; // @[Monitor.scala 713:27:freechips.rocketchip.system.DefaultRV32Config.fir@12305.4]
  wire [3:0] _T_1893; // @[Monitor.scala 713:38:freechips.rocketchip.system.DefaultRV32Config.fir@12306.4]
  wire [3:0] _T_1894; // @[Monitor.scala 713:36:freechips.rocketchip.system.DefaultRV32Config.fir@12307.4]
  wire  _GEN_85; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@9501.10]
  wire  _GEN_101; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@9630.10]
  wire  _GEN_119; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@9770.10]
  wire  _GEN_131; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@9877.10]
  wire  _GEN_141; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@9976.10]
  wire  _GEN_151; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@10067.10]
  wire  _GEN_161; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@10156.10]
  wire  _GEN_171; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@10245.10]
  wire  _GEN_183; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@10314.10]
  wire  _GEN_193; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@10356.10]
  wire  _GEN_203; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@10414.10]
  wire  _GEN_213; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@10473.10]
  wire  _GEN_219; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@10508.10]
  wire  _GEN_225; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@10544.10]
  wire  _GEN_231; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@11199.10]
  wire  _GEN_243; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@11247.10]
  wire  _GEN_253; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@11336.10]
  wire  _GEN_267; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@11456.10]
  wire  _GEN_279; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@11519.10]
  wire  _GEN_289; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@11559.10]
  wire  _GEN_297; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@11591.10]
  plusarg_reader #(.FORMAT("tilelink_timeout=%d"), .DEFAULT(0), .WIDTH(32)) plusarg_reader ( // @[PlusArg.scala 80:11:freechips.rocketchip.system.DefaultRV32Config.fir@12216.4]
    .out(plusarg_reader_out)
  );
  assign _T_4 = io_in_a_bits_source == 2'h0; // @[Parameters.scala 47:9:freechips.rocketchip.system.DefaultRV32Config.fir@9364.6]
  assign _T_5 = io_in_a_bits_source == 2'h1; // @[Parameters.scala 47:9:freechips.rocketchip.system.DefaultRV32Config.fir@9365.6]
  assign _T_6 = io_in_a_bits_source == 2'h2; // @[Parameters.scala 47:9:freechips.rocketchip.system.DefaultRV32Config.fir@9366.6]
  assign _T_8 = _T_4 | _T_5; // @[Parameters.scala 924:46:freechips.rocketchip.system.DefaultRV32Config.fir@9372.6]
  assign _T_9 = _T_8 | _T_6; // @[Parameters.scala 924:46:freechips.rocketchip.system.DefaultRV32Config.fir@9373.6]
  assign _T_11 = 27'hfff << io_in_a_bits_size; // @[package.scala 207:77:freechips.rocketchip.system.DefaultRV32Config.fir@9375.6]
  assign _T_13 = ~_T_11[11:0]; // @[package.scala 207:46:freechips.rocketchip.system.DefaultRV32Config.fir@9377.6]
  assign _GEN_71 = {{20'd0}, _T_13}; // @[Edges.scala 22:16:freechips.rocketchip.system.DefaultRV32Config.fir@9378.6]
  assign _T_14 = io_in_a_bits_address & _GEN_71; // @[Edges.scala 22:16:freechips.rocketchip.system.DefaultRV32Config.fir@9378.6]
  assign _T_15 = _T_14 == 32'h0; // @[Edges.scala 22:24:freechips.rocketchip.system.DefaultRV32Config.fir@9379.6]
  assign _T_18 = 2'h1 << io_in_a_bits_size[0]; // @[OneHot.scala 65:12:freechips.rocketchip.system.DefaultRV32Config.fir@9382.6]
  assign _T_20 = _T_18 | 2'h1; // @[Misc.scala 201:81:freechips.rocketchip.system.DefaultRV32Config.fir@9384.6]
  assign _T_21 = io_in_a_bits_size >= 4'h2; // @[Misc.scala 205:21:freechips.rocketchip.system.DefaultRV32Config.fir@9385.6]
  assign _T_24 = ~io_in_a_bits_address[1]; // @[Misc.scala 210:20:freechips.rocketchip.system.DefaultRV32Config.fir@9388.6]
  assign _T_26 = _T_20[1] & _T_24; // @[Misc.scala 214:38:freechips.rocketchip.system.DefaultRV32Config.fir@9390.6]
  assign _T_27 = _T_21 | _T_26; // @[Misc.scala 214:29:freechips.rocketchip.system.DefaultRV32Config.fir@9391.6]
  assign _T_29 = _T_20[1] & io_in_a_bits_address[1]; // @[Misc.scala 214:38:freechips.rocketchip.system.DefaultRV32Config.fir@9393.6]
  assign _T_30 = _T_21 | _T_29; // @[Misc.scala 214:29:freechips.rocketchip.system.DefaultRV32Config.fir@9394.6]
  assign _T_33 = ~io_in_a_bits_address[0]; // @[Misc.scala 210:20:freechips.rocketchip.system.DefaultRV32Config.fir@9397.6]
  assign _T_34 = _T_24 & _T_33; // @[Misc.scala 213:27:freechips.rocketchip.system.DefaultRV32Config.fir@9398.6]
  assign _T_35 = _T_20[0] & _T_34; // @[Misc.scala 214:38:freechips.rocketchip.system.DefaultRV32Config.fir@9399.6]
  assign _T_36 = _T_27 | _T_35; // @[Misc.scala 214:29:freechips.rocketchip.system.DefaultRV32Config.fir@9400.6]
  assign _T_37 = _T_24 & io_in_a_bits_address[0]; // @[Misc.scala 213:27:freechips.rocketchip.system.DefaultRV32Config.fir@9401.6]
  assign _T_38 = _T_20[0] & _T_37; // @[Misc.scala 214:38:freechips.rocketchip.system.DefaultRV32Config.fir@9402.6]
  assign _T_39 = _T_27 | _T_38; // @[Misc.scala 214:29:freechips.rocketchip.system.DefaultRV32Config.fir@9403.6]
  assign _T_40 = io_in_a_bits_address[1] & _T_33; // @[Misc.scala 213:27:freechips.rocketchip.system.DefaultRV32Config.fir@9404.6]
  assign _T_41 = _T_20[0] & _T_40; // @[Misc.scala 214:38:freechips.rocketchip.system.DefaultRV32Config.fir@9405.6]
  assign _T_42 = _T_30 | _T_41; // @[Misc.scala 214:29:freechips.rocketchip.system.DefaultRV32Config.fir@9406.6]
  assign _T_43 = io_in_a_bits_address[1] & io_in_a_bits_address[0]; // @[Misc.scala 213:27:freechips.rocketchip.system.DefaultRV32Config.fir@9407.6]
  assign _T_44 = _T_20[0] & _T_43; // @[Misc.scala 214:38:freechips.rocketchip.system.DefaultRV32Config.fir@9408.6]
  assign _T_45 = _T_30 | _T_44; // @[Misc.scala 214:29:freechips.rocketchip.system.DefaultRV32Config.fir@9409.6]
  assign _T_48 = {_T_45,_T_42,_T_39,_T_36}; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@9412.6]
  assign _T_52 = {1'b0,$signed(io_in_a_bits_address)}; // @[Parameters.scala 137:49:freechips.rocketchip.system.DefaultRV32Config.fir@9416.6]
  assign _T_78 = io_in_a_bits_opcode == 3'h6; // @[Monitor.scala 79:25:freechips.rocketchip.system.DefaultRV32Config.fir@9446.6]
  assign _T_83 = $signed(_T_52) & -33'sh1000; // @[Parameters.scala 137:52:freechips.rocketchip.system.DefaultRV32Config.fir@9452.8]
  assign _T_84 = $signed(_T_83) == 33'sh0; // @[Parameters.scala 137:67:freechips.rocketchip.system.DefaultRV32Config.fir@9453.8]
  assign _T_85 = io_in_a_bits_address ^ 32'h3000; // @[Parameters.scala 137:31:freechips.rocketchip.system.DefaultRV32Config.fir@9454.8]
  assign _T_86 = {1'b0,$signed(_T_85)}; // @[Parameters.scala 137:49:freechips.rocketchip.system.DefaultRV32Config.fir@9455.8]
  assign _T_88 = $signed(_T_86) & -33'sh1000; // @[Parameters.scala 137:52:freechips.rocketchip.system.DefaultRV32Config.fir@9457.8]
  assign _T_89 = $signed(_T_88) == 33'sh0; // @[Parameters.scala 137:67:freechips.rocketchip.system.DefaultRV32Config.fir@9458.8]
  assign _T_90 = io_in_a_bits_address ^ 32'h10000; // @[Parameters.scala 137:31:freechips.rocketchip.system.DefaultRV32Config.fir@9459.8]
  assign _T_91 = {1'b0,$signed(_T_90)}; // @[Parameters.scala 137:49:freechips.rocketchip.system.DefaultRV32Config.fir@9460.8]
  assign _T_93 = $signed(_T_91) & -33'sh10000; // @[Parameters.scala 137:52:freechips.rocketchip.system.DefaultRV32Config.fir@9462.8]
  assign _T_94 = $signed(_T_93) == 33'sh0; // @[Parameters.scala 137:67:freechips.rocketchip.system.DefaultRV32Config.fir@9463.8]
  assign _T_95 = io_in_a_bits_address ^ 32'h2000000; // @[Parameters.scala 137:31:freechips.rocketchip.system.DefaultRV32Config.fir@9464.8]
  assign _T_96 = {1'b0,$signed(_T_95)}; // @[Parameters.scala 137:49:freechips.rocketchip.system.DefaultRV32Config.fir@9465.8]
  assign _T_98 = $signed(_T_96) & -33'sh10000; // @[Parameters.scala 137:52:freechips.rocketchip.system.DefaultRV32Config.fir@9467.8]
  assign _T_99 = $signed(_T_98) == 33'sh0; // @[Parameters.scala 137:67:freechips.rocketchip.system.DefaultRV32Config.fir@9468.8]
  assign _T_100 = io_in_a_bits_address ^ 32'hc000000; // @[Parameters.scala 137:31:freechips.rocketchip.system.DefaultRV32Config.fir@9469.8]
  assign _T_101 = {1'b0,$signed(_T_100)}; // @[Parameters.scala 137:49:freechips.rocketchip.system.DefaultRV32Config.fir@9470.8]
  assign _T_103 = $signed(_T_101) & -33'sh4000000; // @[Parameters.scala 137:52:freechips.rocketchip.system.DefaultRV32Config.fir@9472.8]
  assign _T_104 = $signed(_T_103) == 33'sh0; // @[Parameters.scala 137:67:freechips.rocketchip.system.DefaultRV32Config.fir@9473.8]
  assign _T_105 = io_in_a_bits_address ^ 32'h60000000; // @[Parameters.scala 137:31:freechips.rocketchip.system.DefaultRV32Config.fir@9474.8]
  assign _T_106 = {1'b0,$signed(_T_105)}; // @[Parameters.scala 137:49:freechips.rocketchip.system.DefaultRV32Config.fir@9475.8]
  assign _T_108 = $signed(_T_106) & -33'sh20000000; // @[Parameters.scala 137:52:freechips.rocketchip.system.DefaultRV32Config.fir@9477.8]
  assign _T_109 = $signed(_T_108) == 33'sh0; // @[Parameters.scala 137:67:freechips.rocketchip.system.DefaultRV32Config.fir@9478.8]
  assign _T_110 = _T_84 | _T_89; // @[Parameters.scala 552:42:freechips.rocketchip.system.DefaultRV32Config.fir@9479.8]
  assign _T_117 = io_in_a_bits_size <= 4'h6; // @[Parameters.scala 93:42:freechips.rocketchip.system.DefaultRV32Config.fir@9486.8]
  assign _T_120 = io_in_a_bits_address ^ 32'h80000000; // @[Parameters.scala 137:31:freechips.rocketchip.system.DefaultRV32Config.fir@9489.8]
  assign _T_121 = {1'b0,$signed(_T_120)}; // @[Parameters.scala 137:49:freechips.rocketchip.system.DefaultRV32Config.fir@9490.8]
  assign _T_123 = $signed(_T_121) & -33'sh10000000; // @[Parameters.scala 137:52:freechips.rocketchip.system.DefaultRV32Config.fir@9492.8]
  assign _T_124 = $signed(_T_123) == 33'sh0; // @[Parameters.scala 137:67:freechips.rocketchip.system.DefaultRV32Config.fir@9493.8]
  assign _T_125 = _T_117 & _T_124; // @[Parameters.scala 551:56:freechips.rocketchip.system.DefaultRV32Config.fir@9494.8]
  assign _T_129 = _T_125 | reset; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@9498.8]
  assign _T_130 = ~_T_129; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@9499.8]
  assign _T_135 = 4'h6 == io_in_a_bits_size; // @[Parameters.scala 92:48:freechips.rocketchip.system.DefaultRV32Config.fir@9512.8]
  assign _T_136 = _T_4 & _T_135; // @[Mux.scala 27:72:freechips.rocketchip.system.DefaultRV32Config.fir@9513.8]
  assign _T_143 = _T_136 | reset; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@9521.8]
  assign _T_144 = ~_T_143; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@9522.8]
  assign _T_146 = _T_9 | reset; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@9528.8]
  assign _T_147 = ~_T_146; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@9529.8]
  assign _T_150 = _T_21 | reset; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@9536.8]
  assign _T_151 = ~_T_150; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@9537.8]
  assign _T_153 = _T_15 | reset; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@9543.8]
  assign _T_154 = ~_T_153; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@9544.8]
  assign _T_155 = io_in_a_bits_param <= 3'h2; // @[Bundles.scala 110:27:freechips.rocketchip.system.DefaultRV32Config.fir@9549.8]
  assign _T_157 = _T_155 | reset; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@9551.8]
  assign _T_158 = ~_T_157; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@9552.8]
  assign _T_159 = ~io_in_a_bits_mask; // @[Monitor.scala 86:18:freechips.rocketchip.system.DefaultRV32Config.fir@9557.8]
  assign _T_160 = _T_159 == 4'h0; // @[Monitor.scala 86:31:freechips.rocketchip.system.DefaultRV32Config.fir@9558.8]
  assign _T_162 = _T_160 | reset; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@9560.8]
  assign _T_163 = ~_T_162; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@9561.8]
  assign _T_164 = ~io_in_a_bits_corrupt; // @[Monitor.scala 87:18:freechips.rocketchip.system.DefaultRV32Config.fir@9566.8]
  assign _T_166 = _T_164 | reset; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@9568.8]
  assign _T_167 = ~_T_166; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@9569.8]
  assign _T_168 = io_in_a_bits_opcode == 3'h7; // @[Monitor.scala 90:25:freechips.rocketchip.system.DefaultRV32Config.fir@9575.6]
  assign _T_249 = io_in_a_bits_param != 3'h0; // @[Monitor.scala 97:31:freechips.rocketchip.system.DefaultRV32Config.fir@9686.8]
  assign _T_251 = _T_249 | reset; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@9688.8]
  assign _T_252 = ~_T_251; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@9689.8]
  assign _T_262 = io_in_a_bits_opcode == 3'h4; // @[Monitor.scala 102:25:freechips.rocketchip.system.DefaultRV32Config.fir@9712.6]
  assign _T_264 = io_in_a_bits_size <= 4'hc; // @[Parameters.scala 93:42:freechips.rocketchip.system.DefaultRV32Config.fir@9715.8]
  assign _T_272 = _T_264 & _T_89; // @[Parameters.scala 551:56:freechips.rocketchip.system.DefaultRV32Config.fir@9723.8]
  assign _T_307 = _T_84 | _T_94; // @[Parameters.scala 552:42:freechips.rocketchip.system.DefaultRV32Config.fir@9758.8]
  assign _T_308 = _T_307 | _T_99; // @[Parameters.scala 552:42:freechips.rocketchip.system.DefaultRV32Config.fir@9759.8]
  assign _T_309 = _T_308 | _T_104; // @[Parameters.scala 552:42:freechips.rocketchip.system.DefaultRV32Config.fir@9760.8]
  assign _T_310 = _T_309 | _T_109; // @[Parameters.scala 552:42:freechips.rocketchip.system.DefaultRV32Config.fir@9761.8]
  assign _T_311 = _T_310 | _T_124; // @[Parameters.scala 552:42:freechips.rocketchip.system.DefaultRV32Config.fir@9762.8]
  assign _T_312 = _T_117 & _T_311; // @[Parameters.scala 551:56:freechips.rocketchip.system.DefaultRV32Config.fir@9763.8]
  assign _T_314 = _T_272 | _T_312; // @[Parameters.scala 553:30:freechips.rocketchip.system.DefaultRV32Config.fir@9765.8]
  assign _T_316 = _T_314 | reset; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@9767.8]
  assign _T_317 = ~_T_316; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@9768.8]
  assign _T_324 = io_in_a_bits_param == 3'h0; // @[Monitor.scala 106:31:freechips.rocketchip.system.DefaultRV32Config.fir@9787.8]
  assign _T_326 = _T_324 | reset; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@9789.8]
  assign _T_327 = ~_T_326; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@9790.8]
  assign _T_328 = io_in_a_bits_mask == _T_48; // @[Monitor.scala 107:30:freechips.rocketchip.system.DefaultRV32Config.fir@9795.8]
  assign _T_330 = _T_328 | reset; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@9797.8]
  assign _T_331 = ~_T_330; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@9798.8]
  assign _T_336 = io_in_a_bits_opcode == 3'h0; // @[Monitor.scala 111:25:freechips.rocketchip.system.DefaultRV32Config.fir@9812.6]
  assign _T_371 = _T_84 | _T_99; // @[Parameters.scala 552:42:freechips.rocketchip.system.DefaultRV32Config.fir@9848.8]
  assign _T_372 = _T_371 | _T_104; // @[Parameters.scala 552:42:freechips.rocketchip.system.DefaultRV32Config.fir@9849.8]
  assign _T_373 = _T_372 | _T_124; // @[Parameters.scala 552:42:freechips.rocketchip.system.DefaultRV32Config.fir@9850.8]
  assign _T_374 = _T_117 & _T_373; // @[Parameters.scala 551:56:freechips.rocketchip.system.DefaultRV32Config.fir@9851.8]
  assign _T_383 = io_in_a_bits_size <= 4'h8; // @[Parameters.scala 93:42:freechips.rocketchip.system.DefaultRV32Config.fir@9860.8]
  assign _T_391 = _T_383 & _T_109; // @[Parameters.scala 551:56:freechips.rocketchip.system.DefaultRV32Config.fir@9868.8]
  assign _T_393 = _T_272 | _T_374; // @[Parameters.scala 553:30:freechips.rocketchip.system.DefaultRV32Config.fir@9870.8]
  assign _T_395 = _T_393 | _T_391; // @[Parameters.scala 553:30:freechips.rocketchip.system.DefaultRV32Config.fir@9872.8]
  assign _T_397 = _T_395 | reset; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@9874.8]
  assign _T_398 = ~_T_397; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@9875.8]
  assign _T_413 = io_in_a_bits_opcode == 3'h1; // @[Monitor.scala 119:25:freechips.rocketchip.system.DefaultRV32Config.fir@9911.6]
  assign _T_486 = ~_T_48; // @[Monitor.scala 124:33:freechips.rocketchip.system.DefaultRV32Config.fir@10001.8]
  assign _T_487 = io_in_a_bits_mask & _T_486; // @[Monitor.scala 124:31:freechips.rocketchip.system.DefaultRV32Config.fir@10002.8]
  assign _T_488 = _T_487 == 4'h0; // @[Monitor.scala 124:40:freechips.rocketchip.system.DefaultRV32Config.fir@10003.8]
  assign _T_490 = _T_488 | reset; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@10005.8]
  assign _T_491 = ~_T_490; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@10006.8]
  assign _T_492 = io_in_a_bits_opcode == 3'h2; // @[Monitor.scala 127:25:freechips.rocketchip.system.DefaultRV32Config.fir@10012.6]
  assign _T_494 = io_in_a_bits_size <= 4'h2; // @[Parameters.scala 93:42:freechips.rocketchip.system.DefaultRV32Config.fir@10015.8]
  assign _T_518 = _T_110 | _T_99; // @[Parameters.scala 552:42:freechips.rocketchip.system.DefaultRV32Config.fir@10039.8]
  assign _T_519 = _T_518 | _T_104; // @[Parameters.scala 552:42:freechips.rocketchip.system.DefaultRV32Config.fir@10040.8]
  assign _T_520 = _T_494 & _T_519; // @[Parameters.scala 551:56:freechips.rocketchip.system.DefaultRV32Config.fir@10041.8]
  assign _T_543 = _T_520 | reset; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@10064.8]
  assign _T_544 = ~_T_543; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@10065.8]
  assign _T_551 = io_in_a_bits_param <= 3'h4; // @[Bundles.scala 140:33:freechips.rocketchip.system.DefaultRV32Config.fir@10084.8]
  assign _T_553 = _T_551 | reset; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@10086.8]
  assign _T_554 = ~_T_553; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@10087.8]
  assign _T_559 = io_in_a_bits_opcode == 3'h3; // @[Monitor.scala 135:25:freechips.rocketchip.system.DefaultRV32Config.fir@10101.6]
  assign _T_618 = io_in_a_bits_param <= 3'h3; // @[Bundles.scala 147:30:freechips.rocketchip.system.DefaultRV32Config.fir@10173.8]
  assign _T_620 = _T_618 | reset; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@10175.8]
  assign _T_621 = ~_T_620; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@10176.8]
  assign _T_626 = io_in_a_bits_opcode == 3'h5; // @[Monitor.scala 143:25:freechips.rocketchip.system.DefaultRV32Config.fir@10190.6]
  assign _T_677 = _T_272 | reset; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@10242.8]
  assign _T_678 = ~_T_677; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@10243.8]
  assign _T_685 = io_in_a_bits_param <= 3'h1; // @[Bundles.scala 160:28:freechips.rocketchip.system.DefaultRV32Config.fir@10262.8]
  assign _T_687 = _T_685 | reset; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@10264.8]
  assign _T_688 = ~_T_687; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@10265.8]
  assign _T_697 = io_in_d_bits_opcode <= 3'h6; // @[Bundles.scala 44:24:freechips.rocketchip.system.DefaultRV32Config.fir@10289.6]
  assign _T_699 = _T_697 | reset; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@10291.6]
  assign _T_700 = ~_T_699; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@10292.6]
  assign _T_701 = io_in_d_bits_source == 2'h0; // @[Parameters.scala 47:9:freechips.rocketchip.system.DefaultRV32Config.fir@10297.6]
  assign _T_702 = io_in_d_bits_source == 2'h1; // @[Parameters.scala 47:9:freechips.rocketchip.system.DefaultRV32Config.fir@10298.6]
  assign _T_703 = io_in_d_bits_source == 2'h2; // @[Parameters.scala 47:9:freechips.rocketchip.system.DefaultRV32Config.fir@10299.6]
  assign _T_705 = _T_701 | _T_702; // @[Parameters.scala 924:46:freechips.rocketchip.system.DefaultRV32Config.fir@10305.6]
  assign _T_706 = _T_705 | _T_703; // @[Parameters.scala 924:46:freechips.rocketchip.system.DefaultRV32Config.fir@10306.6]
  assign _T_708 = io_in_d_bits_opcode == 3'h6; // @[Monitor.scala 307:25:freechips.rocketchip.system.DefaultRV32Config.fir@10308.6]
  assign _T_710 = _T_706 | reset; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@10311.8]
  assign _T_711 = ~_T_710; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@10312.8]
  assign _T_712 = io_in_d_bits_size >= 4'h2; // @[Monitor.scala 309:27:freechips.rocketchip.system.DefaultRV32Config.fir@10317.8]
  assign _T_714 = _T_712 | reset; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@10319.8]
  assign _T_715 = ~_T_714; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@10320.8]
  assign _T_716 = io_in_d_bits_param == 2'h0; // @[Monitor.scala 310:28:freechips.rocketchip.system.DefaultRV32Config.fir@10325.8]
  assign _T_718 = _T_716 | reset; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@10327.8]
  assign _T_719 = ~_T_718; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@10328.8]
  assign _T_720 = ~io_in_d_bits_corrupt; // @[Monitor.scala 311:15:freechips.rocketchip.system.DefaultRV32Config.fir@10333.8]
  assign _T_722 = _T_720 | reset; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@10335.8]
  assign _T_723 = ~_T_722; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@10336.8]
  assign _T_724 = ~io_in_d_bits_denied; // @[Monitor.scala 312:15:freechips.rocketchip.system.DefaultRV32Config.fir@10341.8]
  assign _T_726 = _T_724 | reset; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@10343.8]
  assign _T_727 = ~_T_726; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@10344.8]
  assign _T_728 = io_in_d_bits_opcode == 3'h4; // @[Monitor.scala 315:25:freechips.rocketchip.system.DefaultRV32Config.fir@10350.6]
  assign _T_739 = io_in_d_bits_param <= 2'h2; // @[Bundles.scala 104:26:freechips.rocketchip.system.DefaultRV32Config.fir@10374.8]
  assign _T_741 = _T_739 | reset; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@10376.8]
  assign _T_742 = ~_T_741; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@10377.8]
  assign _T_743 = io_in_d_bits_param != 2'h2; // @[Monitor.scala 320:28:freechips.rocketchip.system.DefaultRV32Config.fir@10382.8]
  assign _T_745 = _T_743 | reset; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@10384.8]
  assign _T_746 = ~_T_745; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@10385.8]
  assign _T_756 = io_in_d_bits_opcode == 3'h5; // @[Monitor.scala 325:25:freechips.rocketchip.system.DefaultRV32Config.fir@10408.6]
  assign _T_776 = _T_724 | io_in_d_bits_corrupt; // @[Monitor.scala 331:30:freechips.rocketchip.system.DefaultRV32Config.fir@10449.8]
  assign _T_778 = _T_776 | reset; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@10451.8]
  assign _T_779 = ~_T_778; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@10452.8]
  assign _T_785 = io_in_d_bits_opcode == 3'h0; // @[Monitor.scala 335:25:freechips.rocketchip.system.DefaultRV32Config.fir@10467.6]
  assign _T_802 = io_in_d_bits_opcode == 3'h1; // @[Monitor.scala 343:25:freechips.rocketchip.system.DefaultRV32Config.fir@10502.6]
  assign _T_820 = io_in_d_bits_opcode == 3'h2; // @[Monitor.scala 351:25:freechips.rocketchip.system.DefaultRV32Config.fir@10538.6]
  assign _T_844 = {1'b0,$signed(io_in_b_bits_address)}; // @[Parameters.scala 137:49:freechips.rocketchip.system.DefaultRV32Config.fir@10586.6]
  assign _T_870 = io_in_b_bits_address ^ 32'h3000; // @[Parameters.scala 137:31:freechips.rocketchip.system.DefaultRV32Config.fir@10616.6]
  assign _T_871 = {1'b0,$signed(_T_870)}; // @[Parameters.scala 137:49:freechips.rocketchip.system.DefaultRV32Config.fir@10617.6]
  assign _T_873 = $signed(_T_871) & -33'sh1000; // @[Parameters.scala 137:52:freechips.rocketchip.system.DefaultRV32Config.fir@10619.6]
  assign _T_874 = $signed(_T_873) == 33'sh0; // @[Parameters.scala 137:67:freechips.rocketchip.system.DefaultRV32Config.fir@10620.6]
  assign _T_875 = io_in_b_bits_address ^ 32'hc000000; // @[Parameters.scala 137:31:freechips.rocketchip.system.DefaultRV32Config.fir@10621.6]
  assign _T_876 = {1'b0,$signed(_T_875)}; // @[Parameters.scala 137:49:freechips.rocketchip.system.DefaultRV32Config.fir@10622.6]
  assign _T_878 = $signed(_T_876) & -33'sh4000000; // @[Parameters.scala 137:52:freechips.rocketchip.system.DefaultRV32Config.fir@10624.6]
  assign _T_879 = $signed(_T_878) == 33'sh0; // @[Parameters.scala 137:67:freechips.rocketchip.system.DefaultRV32Config.fir@10625.6]
  assign _T_880 = io_in_b_bits_address ^ 32'h2000000; // @[Parameters.scala 137:31:freechips.rocketchip.system.DefaultRV32Config.fir@10626.6]
  assign _T_881 = {1'b0,$signed(_T_880)}; // @[Parameters.scala 137:49:freechips.rocketchip.system.DefaultRV32Config.fir@10627.6]
  assign _T_883 = $signed(_T_881) & -33'sh10000; // @[Parameters.scala 137:52:freechips.rocketchip.system.DefaultRV32Config.fir@10629.6]
  assign _T_884 = $signed(_T_883) == 33'sh0; // @[Parameters.scala 137:67:freechips.rocketchip.system.DefaultRV32Config.fir@10630.6]
  assign _T_888 = $signed(_T_844) & -33'sh1000; // @[Parameters.scala 137:52:freechips.rocketchip.system.DefaultRV32Config.fir@10634.6]
  assign _T_889 = $signed(_T_888) == 33'sh0; // @[Parameters.scala 137:67:freechips.rocketchip.system.DefaultRV32Config.fir@10635.6]
  assign _T_890 = io_in_b_bits_address ^ 32'h10000; // @[Parameters.scala 137:31:freechips.rocketchip.system.DefaultRV32Config.fir@10636.6]
  assign _T_891 = {1'b0,$signed(_T_890)}; // @[Parameters.scala 137:49:freechips.rocketchip.system.DefaultRV32Config.fir@10637.6]
  assign _T_893 = $signed(_T_891) & -33'sh10000; // @[Parameters.scala 137:52:freechips.rocketchip.system.DefaultRV32Config.fir@10639.6]
  assign _T_894 = $signed(_T_893) == 33'sh0; // @[Parameters.scala 137:67:freechips.rocketchip.system.DefaultRV32Config.fir@10640.6]
  assign _T_895 = io_in_b_bits_address ^ 32'h80000000; // @[Parameters.scala 137:31:freechips.rocketchip.system.DefaultRV32Config.fir@10641.6]
  assign _T_896 = {1'b0,$signed(_T_895)}; // @[Parameters.scala 137:49:freechips.rocketchip.system.DefaultRV32Config.fir@10642.6]
  assign _T_898 = $signed(_T_896) & -33'sh10000000; // @[Parameters.scala 137:52:freechips.rocketchip.system.DefaultRV32Config.fir@10644.6]
  assign _T_899 = $signed(_T_898) == 33'sh0; // @[Parameters.scala 137:67:freechips.rocketchip.system.DefaultRV32Config.fir@10645.6]
  assign _T_900 = io_in_b_bits_address ^ 32'h60000000; // @[Parameters.scala 137:31:freechips.rocketchip.system.DefaultRV32Config.fir@10646.6]
  assign _T_901 = {1'b0,$signed(_T_900)}; // @[Parameters.scala 137:49:freechips.rocketchip.system.DefaultRV32Config.fir@10647.6]
  assign _T_903 = $signed(_T_901) & -33'sh20000000; // @[Parameters.scala 137:52:freechips.rocketchip.system.DefaultRV32Config.fir@10649.6]
  assign _T_904 = $signed(_T_903) == 33'sh0; // @[Parameters.scala 137:67:freechips.rocketchip.system.DefaultRV32Config.fir@10650.6]
  assign _T_906 = _T_874 | _T_879; // @[Parameters.scala 535:64:freechips.rocketchip.system.DefaultRV32Config.fir@10660.6]
  assign _T_907 = _T_906 | _T_884; // @[Parameters.scala 535:64:freechips.rocketchip.system.DefaultRV32Config.fir@10661.6]
  assign _T_908 = _T_907 | _T_889; // @[Parameters.scala 535:64:freechips.rocketchip.system.DefaultRV32Config.fir@10662.6]
  assign _T_909 = _T_908 | _T_894; // @[Parameters.scala 535:64:freechips.rocketchip.system.DefaultRV32Config.fir@10663.6]
  assign _T_910 = _T_909 | _T_899; // @[Parameters.scala 535:64:freechips.rocketchip.system.DefaultRV32Config.fir@10664.6]
  assign _T_911 = _T_910 | _T_904; // @[Parameters.scala 535:64:freechips.rocketchip.system.DefaultRV32Config.fir@10665.6]
  assign _T_916 = io_in_b_bits_address & 32'h3f; // @[Edges.scala 22:16:freechips.rocketchip.system.DefaultRV32Config.fir@10670.6]
  assign _T_917 = _T_916 == 32'h0; // @[Edges.scala 22:24:freechips.rocketchip.system.DefaultRV32Config.fir@10671.6]
  assign _T_978 = _T_911 | reset; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@10747.8]
  assign _T_979 = ~_T_978; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@10748.8]
  assign _T_984 = _T_917 | reset; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@10761.8]
  assign _T_985 = ~_T_984; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@10762.8]
  assign _T_986 = io_in_b_bits_param <= 2'h2; // @[Bundles.scala 104:26:freechips.rocketchip.system.DefaultRV32Config.fir@10767.8]
  assign _T_988 = _T_986 | reset; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@10769.8]
  assign _T_989 = ~_T_988; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@10770.8]
  assign _T_1134 = io_in_c_bits_source == 2'h0; // @[Parameters.scala 47:9:freechips.rocketchip.system.DefaultRV32Config.fir@11094.6]
  assign _T_1135 = io_in_c_bits_source == 2'h1; // @[Parameters.scala 47:9:freechips.rocketchip.system.DefaultRV32Config.fir@11095.6]
  assign _T_1136 = io_in_c_bits_source == 2'h2; // @[Parameters.scala 47:9:freechips.rocketchip.system.DefaultRV32Config.fir@11096.6]
  assign _T_1138 = _T_1134 | _T_1135; // @[Parameters.scala 924:46:freechips.rocketchip.system.DefaultRV32Config.fir@11102.6]
  assign _T_1139 = _T_1138 | _T_1136; // @[Parameters.scala 924:46:freechips.rocketchip.system.DefaultRV32Config.fir@11103.6]
  assign _T_1141 = 27'hfff << io_in_c_bits_size; // @[package.scala 207:77:freechips.rocketchip.system.DefaultRV32Config.fir@11105.6]
  assign _T_1143 = ~_T_1141[11:0]; // @[package.scala 207:46:freechips.rocketchip.system.DefaultRV32Config.fir@11107.6]
  assign _GEN_72 = {{20'd0}, _T_1143}; // @[Edges.scala 22:16:freechips.rocketchip.system.DefaultRV32Config.fir@11108.6]
  assign _T_1144 = io_in_c_bits_address & _GEN_72; // @[Edges.scala 22:16:freechips.rocketchip.system.DefaultRV32Config.fir@11108.6]
  assign _T_1145 = _T_1144 == 32'h0; // @[Edges.scala 22:24:freechips.rocketchip.system.DefaultRV32Config.fir@11109.6]
  assign _T_1146 = io_in_c_bits_address ^ 32'h3000; // @[Parameters.scala 137:31:freechips.rocketchip.system.DefaultRV32Config.fir@11110.6]
  assign _T_1147 = {1'b0,$signed(_T_1146)}; // @[Parameters.scala 137:49:freechips.rocketchip.system.DefaultRV32Config.fir@11111.6]
  assign _T_1149 = $signed(_T_1147) & -33'sh1000; // @[Parameters.scala 137:52:freechips.rocketchip.system.DefaultRV32Config.fir@11113.6]
  assign _T_1150 = $signed(_T_1149) == 33'sh0; // @[Parameters.scala 137:67:freechips.rocketchip.system.DefaultRV32Config.fir@11114.6]
  assign _T_1151 = io_in_c_bits_address ^ 32'hc000000; // @[Parameters.scala 137:31:freechips.rocketchip.system.DefaultRV32Config.fir@11115.6]
  assign _T_1152 = {1'b0,$signed(_T_1151)}; // @[Parameters.scala 137:49:freechips.rocketchip.system.DefaultRV32Config.fir@11116.6]
  assign _T_1154 = $signed(_T_1152) & -33'sh4000000; // @[Parameters.scala 137:52:freechips.rocketchip.system.DefaultRV32Config.fir@11118.6]
  assign _T_1155 = $signed(_T_1154) == 33'sh0; // @[Parameters.scala 137:67:freechips.rocketchip.system.DefaultRV32Config.fir@11119.6]
  assign _T_1156 = io_in_c_bits_address ^ 32'h2000000; // @[Parameters.scala 137:31:freechips.rocketchip.system.DefaultRV32Config.fir@11120.6]
  assign _T_1157 = {1'b0,$signed(_T_1156)}; // @[Parameters.scala 137:49:freechips.rocketchip.system.DefaultRV32Config.fir@11121.6]
  assign _T_1159 = $signed(_T_1157) & -33'sh10000; // @[Parameters.scala 137:52:freechips.rocketchip.system.DefaultRV32Config.fir@11123.6]
  assign _T_1160 = $signed(_T_1159) == 33'sh0; // @[Parameters.scala 137:67:freechips.rocketchip.system.DefaultRV32Config.fir@11124.6]
  assign _T_1162 = {1'b0,$signed(io_in_c_bits_address)}; // @[Parameters.scala 137:49:freechips.rocketchip.system.DefaultRV32Config.fir@11126.6]
  assign _T_1164 = $signed(_T_1162) & -33'sh1000; // @[Parameters.scala 137:52:freechips.rocketchip.system.DefaultRV32Config.fir@11128.6]
  assign _T_1165 = $signed(_T_1164) == 33'sh0; // @[Parameters.scala 137:67:freechips.rocketchip.system.DefaultRV32Config.fir@11129.6]
  assign _T_1166 = io_in_c_bits_address ^ 32'h10000; // @[Parameters.scala 137:31:freechips.rocketchip.system.DefaultRV32Config.fir@11130.6]
  assign _T_1167 = {1'b0,$signed(_T_1166)}; // @[Parameters.scala 137:49:freechips.rocketchip.system.DefaultRV32Config.fir@11131.6]
  assign _T_1169 = $signed(_T_1167) & -33'sh10000; // @[Parameters.scala 137:52:freechips.rocketchip.system.DefaultRV32Config.fir@11133.6]
  assign _T_1170 = $signed(_T_1169) == 33'sh0; // @[Parameters.scala 137:67:freechips.rocketchip.system.DefaultRV32Config.fir@11134.6]
  assign _T_1171 = io_in_c_bits_address ^ 32'h80000000; // @[Parameters.scala 137:31:freechips.rocketchip.system.DefaultRV32Config.fir@11135.6]
  assign _T_1172 = {1'b0,$signed(_T_1171)}; // @[Parameters.scala 137:49:freechips.rocketchip.system.DefaultRV32Config.fir@11136.6]
  assign _T_1174 = $signed(_T_1172) & -33'sh10000000; // @[Parameters.scala 137:52:freechips.rocketchip.system.DefaultRV32Config.fir@11138.6]
  assign _T_1175 = $signed(_T_1174) == 33'sh0; // @[Parameters.scala 137:67:freechips.rocketchip.system.DefaultRV32Config.fir@11139.6]
  assign _T_1176 = io_in_c_bits_address ^ 32'h60000000; // @[Parameters.scala 137:31:freechips.rocketchip.system.DefaultRV32Config.fir@11140.6]
  assign _T_1177 = {1'b0,$signed(_T_1176)}; // @[Parameters.scala 137:49:freechips.rocketchip.system.DefaultRV32Config.fir@11141.6]
  assign _T_1179 = $signed(_T_1177) & -33'sh20000000; // @[Parameters.scala 137:52:freechips.rocketchip.system.DefaultRV32Config.fir@11143.6]
  assign _T_1180 = $signed(_T_1179) == 33'sh0; // @[Parameters.scala 137:67:freechips.rocketchip.system.DefaultRV32Config.fir@11144.6]
  assign _T_1182 = _T_1150 | _T_1155; // @[Parameters.scala 535:64:freechips.rocketchip.system.DefaultRV32Config.fir@11154.6]
  assign _T_1183 = _T_1182 | _T_1160; // @[Parameters.scala 535:64:freechips.rocketchip.system.DefaultRV32Config.fir@11155.6]
  assign _T_1184 = _T_1183 | _T_1165; // @[Parameters.scala 535:64:freechips.rocketchip.system.DefaultRV32Config.fir@11156.6]
  assign _T_1185 = _T_1184 | _T_1170; // @[Parameters.scala 535:64:freechips.rocketchip.system.DefaultRV32Config.fir@11157.6]
  assign _T_1186 = _T_1185 | _T_1175; // @[Parameters.scala 535:64:freechips.rocketchip.system.DefaultRV32Config.fir@11158.6]
  assign _T_1187 = _T_1186 | _T_1180; // @[Parameters.scala 535:64:freechips.rocketchip.system.DefaultRV32Config.fir@11159.6]
  assign _T_1217 = io_in_c_bits_opcode == 3'h4; // @[Monitor.scala 239:25:freechips.rocketchip.system.DefaultRV32Config.fir@11193.6]
  assign _T_1219 = _T_1187 | reset; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@11196.8]
  assign _T_1220 = ~_T_1219; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@11197.8]
  assign _T_1222 = _T_1139 | reset; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@11203.8]
  assign _T_1223 = ~_T_1222; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@11204.8]
  assign _T_1224 = io_in_c_bits_size >= 4'h2; // @[Monitor.scala 242:30:freechips.rocketchip.system.DefaultRV32Config.fir@11209.8]
  assign _T_1226 = _T_1224 | reset; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@11211.8]
  assign _T_1227 = ~_T_1226; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@11212.8]
  assign _T_1229 = _T_1145 | reset; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@11218.8]
  assign _T_1230 = ~_T_1229; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@11219.8]
  assign _T_1231 = io_in_c_bits_param <= 3'h5; // @[Bundles.scala 122:29:freechips.rocketchip.system.DefaultRV32Config.fir@11224.8]
  assign _T_1233 = _T_1231 | reset; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@11226.8]
  assign _T_1234 = ~_T_1233; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@11227.8]
  assign _T_1235 = ~io_in_c_bits_corrupt; // @[Monitor.scala 245:18:freechips.rocketchip.system.DefaultRV32Config.fir@11232.8]
  assign _T_1237 = _T_1235 | reset; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@11234.8]
  assign _T_1238 = ~_T_1237; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@11235.8]
  assign _T_1239 = io_in_c_bits_opcode == 3'h5; // @[Monitor.scala 248:25:freechips.rocketchip.system.DefaultRV32Config.fir@11241.6]
  assign _T_1257 = io_in_c_bits_opcode == 3'h6; // @[Monitor.scala 256:25:freechips.rocketchip.system.DefaultRV32Config.fir@11281.6]
  assign _T_1296 = io_in_c_bits_size <= 4'h6; // @[Parameters.scala 93:42:freechips.rocketchip.system.DefaultRV32Config.fir@11321.8]
  assign _T_1304 = _T_1296 & _T_1175; // @[Parameters.scala 551:56:freechips.rocketchip.system.DefaultRV32Config.fir@11329.8]
  assign _T_1308 = _T_1304 | reset; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@11333.8]
  assign _T_1309 = ~_T_1308; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@11334.8]
  assign _T_1314 = 4'h6 == io_in_c_bits_size; // @[Parameters.scala 92:48:freechips.rocketchip.system.DefaultRV32Config.fir@11347.8]
  assign _T_1315 = _T_1134 & _T_1314; // @[Mux.scala 27:72:freechips.rocketchip.system.DefaultRV32Config.fir@11348.8]
  assign _T_1322 = _T_1315 | reset; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@11356.8]
  assign _T_1323 = ~_T_1322; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@11357.8]
  assign _T_1334 = io_in_c_bits_param <= 3'h2; // @[Bundles.scala 116:29:freechips.rocketchip.system.DefaultRV32Config.fir@11384.8]
  assign _T_1336 = _T_1334 | reset; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@11386.8]
  assign _T_1337 = ~_T_1336; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@11387.8]
  assign _T_1342 = io_in_c_bits_opcode == 3'h7; // @[Monitor.scala 266:25:freechips.rocketchip.system.DefaultRV32Config.fir@11401.6]
  assign _T_1423 = io_in_c_bits_opcode == 3'h0; // @[Monitor.scala 275:25:freechips.rocketchip.system.DefaultRV32Config.fir@11513.6]
  assign _T_1433 = io_in_c_bits_param == 3'h0; // @[Monitor.scala 279:31:freechips.rocketchip.system.DefaultRV32Config.fir@11536.8]
  assign _T_1435 = _T_1433 | reset; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@11538.8]
  assign _T_1436 = ~_T_1435; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@11539.8]
  assign _T_1441 = io_in_c_bits_opcode == 3'h1; // @[Monitor.scala 283:25:freechips.rocketchip.system.DefaultRV32Config.fir@11553.6]
  assign _T_1455 = io_in_c_bits_opcode == 3'h2; // @[Monitor.scala 290:25:freechips.rocketchip.system.DefaultRV32Config.fir@11585.6]
  assign _T_1477 = io_in_a_ready & io_in_a_valid; // @[Decoupled.scala 40:37:freechips.rocketchip.system.DefaultRV32Config.fir@11636.4]
  assign _T_1484 = ~io_in_a_bits_opcode[2]; // @[Edges.scala 93:28:freechips.rocketchip.system.DefaultRV32Config.fir@11643.4]
  assign _T_1488 = _T_1486 - 10'h1; // @[Edges.scala 231:28:freechips.rocketchip.system.DefaultRV32Config.fir@11647.4]
  assign _T_1489 = _T_1486 == 10'h0; // @[Edges.scala 232:25:freechips.rocketchip.system.DefaultRV32Config.fir@11648.4]
  assign _T_1502 = ~_T_1489; // @[Monitor.scala 386:22:freechips.rocketchip.system.DefaultRV32Config.fir@11664.4]
  assign _T_1503 = io_in_a_valid & _T_1502; // @[Monitor.scala 386:19:freechips.rocketchip.system.DefaultRV32Config.fir@11665.4]
  assign _T_1504 = io_in_a_bits_opcode == _T_1497; // @[Monitor.scala 387:32:freechips.rocketchip.system.DefaultRV32Config.fir@11667.6]
  assign _T_1506 = _T_1504 | reset; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@11669.6]
  assign _T_1507 = ~_T_1506; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@11670.6]
  assign _T_1508 = io_in_a_bits_param == _T_1498; // @[Monitor.scala 388:32:freechips.rocketchip.system.DefaultRV32Config.fir@11675.6]
  assign _T_1510 = _T_1508 | reset; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@11677.6]
  assign _T_1511 = ~_T_1510; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@11678.6]
  assign _T_1512 = io_in_a_bits_size == _T_1499; // @[Monitor.scala 389:32:freechips.rocketchip.system.DefaultRV32Config.fir@11683.6]
  assign _T_1514 = _T_1512 | reset; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@11685.6]
  assign _T_1515 = ~_T_1514; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@11686.6]
  assign _T_1516 = io_in_a_bits_source == _T_1500; // @[Monitor.scala 390:32:freechips.rocketchip.system.DefaultRV32Config.fir@11691.6]
  assign _T_1518 = _T_1516 | reset; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@11693.6]
  assign _T_1519 = ~_T_1518; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@11694.6]
  assign _T_1520 = io_in_a_bits_address == _T_1501; // @[Monitor.scala 391:32:freechips.rocketchip.system.DefaultRV32Config.fir@11699.6]
  assign _T_1522 = _T_1520 | reset; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@11701.6]
  assign _T_1523 = ~_T_1522; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@11702.6]
  assign _T_1525 = _T_1477 & _T_1489; // @[Monitor.scala 393:20:freechips.rocketchip.system.DefaultRV32Config.fir@11709.4]
  assign _T_1526 = io_in_d_ready & io_in_d_valid; // @[Decoupled.scala 40:37:freechips.rocketchip.system.DefaultRV32Config.fir@11717.4]
  assign _T_1528 = 27'hfff << io_in_d_bits_size; // @[package.scala 207:77:freechips.rocketchip.system.DefaultRV32Config.fir@11719.4]
  assign _T_1530 = ~_T_1528[11:0]; // @[package.scala 207:46:freechips.rocketchip.system.DefaultRV32Config.fir@11721.4]
  assign _T_1536 = _T_1534 - 10'h1; // @[Edges.scala 231:28:freechips.rocketchip.system.DefaultRV32Config.fir@11727.4]
  assign _T_1537 = _T_1534 == 10'h0; // @[Edges.scala 232:25:freechips.rocketchip.system.DefaultRV32Config.fir@11728.4]
  assign _T_1551 = ~_T_1537; // @[Monitor.scala 538:22:freechips.rocketchip.system.DefaultRV32Config.fir@11745.4]
  assign _T_1552 = io_in_d_valid & _T_1551; // @[Monitor.scala 538:19:freechips.rocketchip.system.DefaultRV32Config.fir@11746.4]
  assign _T_1553 = io_in_d_bits_opcode == _T_1545; // @[Monitor.scala 539:29:freechips.rocketchip.system.DefaultRV32Config.fir@11748.6]
  assign _T_1555 = _T_1553 | reset; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@11750.6]
  assign _T_1556 = ~_T_1555; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@11751.6]
  assign _T_1557 = io_in_d_bits_param == _T_1546; // @[Monitor.scala 540:29:freechips.rocketchip.system.DefaultRV32Config.fir@11756.6]
  assign _T_1559 = _T_1557 | reset; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@11758.6]
  assign _T_1560 = ~_T_1559; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@11759.6]
  assign _T_1561 = io_in_d_bits_size == _T_1547; // @[Monitor.scala 541:29:freechips.rocketchip.system.DefaultRV32Config.fir@11764.6]
  assign _T_1563 = _T_1561 | reset; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@11766.6]
  assign _T_1564 = ~_T_1563; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@11767.6]
  assign _T_1565 = io_in_d_bits_source == _T_1548; // @[Monitor.scala 542:29:freechips.rocketchip.system.DefaultRV32Config.fir@11772.6]
  assign _T_1567 = _T_1565 | reset; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@11774.6]
  assign _T_1568 = ~_T_1567; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@11775.6]
  assign _T_1569 = io_in_d_bits_sink == _T_1549; // @[Monitor.scala 543:29:freechips.rocketchip.system.DefaultRV32Config.fir@11780.6]
  assign _T_1571 = _T_1569 | reset; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@11782.6]
  assign _T_1572 = ~_T_1571; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@11783.6]
  assign _T_1573 = io_in_d_bits_denied == _T_1550; // @[Monitor.scala 544:29:freechips.rocketchip.system.DefaultRV32Config.fir@11788.6]
  assign _T_1575 = _T_1573 | reset; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@11790.6]
  assign _T_1576 = ~_T_1575; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@11791.6]
  assign _T_1578 = _T_1526 & _T_1537; // @[Monitor.scala 546:20:freechips.rocketchip.system.DefaultRV32Config.fir@11798.4]
  assign _T_1579 = io_in_b_ready & io_in_b_valid; // @[Decoupled.scala 40:37:freechips.rocketchip.system.DefaultRV32Config.fir@11807.4]
  assign _T_1590 = _T_1588 - 10'h1; // @[Edges.scala 231:28:freechips.rocketchip.system.DefaultRV32Config.fir@11818.4]
  assign _T_1591 = _T_1588 == 10'h0; // @[Edges.scala 232:25:freechips.rocketchip.system.DefaultRV32Config.fir@11819.4]
  assign _T_1604 = ~_T_1591; // @[Monitor.scala 409:22:freechips.rocketchip.system.DefaultRV32Config.fir@11835.4]
  assign _T_1605 = io_in_b_valid & _T_1604; // @[Monitor.scala 409:19:freechips.rocketchip.system.DefaultRV32Config.fir@11836.4]
  assign _T_1610 = io_in_b_bits_param == _T_1600; // @[Monitor.scala 411:32:freechips.rocketchip.system.DefaultRV32Config.fir@11846.6]
  assign _T_1612 = _T_1610 | reset; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@11848.6]
  assign _T_1613 = ~_T_1612; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@11849.6]
  assign _T_1622 = io_in_b_bits_address == _T_1603; // @[Monitor.scala 414:32:freechips.rocketchip.system.DefaultRV32Config.fir@11870.6]
  assign _T_1624 = _T_1622 | reset; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@11872.6]
  assign _T_1625 = ~_T_1624; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@11873.6]
  assign _T_1627 = _T_1579 & _T_1591; // @[Monitor.scala 416:20:freechips.rocketchip.system.DefaultRV32Config.fir@11880.4]
  assign _T_1628 = io_in_c_ready & io_in_c_valid; // @[Decoupled.scala 40:37:freechips.rocketchip.system.DefaultRV32Config.fir@11888.4]
  assign _T_1638 = _T_1636 - 10'h1; // @[Edges.scala 231:28:freechips.rocketchip.system.DefaultRV32Config.fir@11898.4]
  assign _T_1639 = _T_1636 == 10'h0; // @[Edges.scala 232:25:freechips.rocketchip.system.DefaultRV32Config.fir@11899.4]
  assign _T_1652 = ~_T_1639; // @[Monitor.scala 514:22:freechips.rocketchip.system.DefaultRV32Config.fir@11915.4]
  assign _T_1653 = io_in_c_valid & _T_1652; // @[Monitor.scala 514:19:freechips.rocketchip.system.DefaultRV32Config.fir@11916.4]
  assign _T_1654 = io_in_c_bits_opcode == _T_1647; // @[Monitor.scala 515:32:freechips.rocketchip.system.DefaultRV32Config.fir@11918.6]
  assign _T_1656 = _T_1654 | reset; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@11920.6]
  assign _T_1657 = ~_T_1656; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@11921.6]
  assign _T_1658 = io_in_c_bits_param == _T_1648; // @[Monitor.scala 516:32:freechips.rocketchip.system.DefaultRV32Config.fir@11926.6]
  assign _T_1660 = _T_1658 | reset; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@11928.6]
  assign _T_1661 = ~_T_1660; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@11929.6]
  assign _T_1662 = io_in_c_bits_size == _T_1649; // @[Monitor.scala 517:32:freechips.rocketchip.system.DefaultRV32Config.fir@11934.6]
  assign _T_1664 = _T_1662 | reset; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@11936.6]
  assign _T_1665 = ~_T_1664; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@11937.6]
  assign _T_1666 = io_in_c_bits_source == _T_1650; // @[Monitor.scala 518:32:freechips.rocketchip.system.DefaultRV32Config.fir@11942.6]
  assign _T_1668 = _T_1666 | reset; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@11944.6]
  assign _T_1669 = ~_T_1668; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@11945.6]
  assign _T_1670 = io_in_c_bits_address == _T_1651; // @[Monitor.scala 519:32:freechips.rocketchip.system.DefaultRV32Config.fir@11950.6]
  assign _T_1672 = _T_1670 | reset; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@11952.6]
  assign _T_1673 = ~_T_1672; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@11953.6]
  assign _T_1675 = _T_1628 & _T_1639; // @[Monitor.scala 521:20:freechips.rocketchip.system.DefaultRV32Config.fir@11960.4]
  assign _T_1687 = _T_1685 - 10'h1; // @[Edges.scala 231:28:freechips.rocketchip.system.DefaultRV32Config.fir@11982.4]
  assign a_first = _T_1685 == 10'h0; // @[Edges.scala 232:25:freechips.rocketchip.system.DefaultRV32Config.fir@11983.4]
  assign _T_1705 = _T_1703 - 10'h1; // @[Edges.scala 231:28:freechips.rocketchip.system.DefaultRV32Config.fir@12004.4]
  assign d_first = _T_1703 == 10'h0; // @[Edges.scala 232:25:freechips.rocketchip.system.DefaultRV32Config.fir@12005.4]
  assign _GEN_73 = {io_in_d_bits_source, 2'h0}; // @[Monitor.scala 629:69:freechips.rocketchip.system.DefaultRV32Config.fir@12024.4]
  assign _T_1713 = {{1'd0}, _GEN_73}; // @[Monitor.scala 629:69:freechips.rocketchip.system.DefaultRV32Config.fir@12024.4]
  assign _T_1714 = inflight_opcodes >> _T_1713; // @[Monitor.scala 629:44:freechips.rocketchip.system.DefaultRV32Config.fir@12025.4]
  assign _T_1718 = 16'h10 - 16'h1; // @[Monitor.scala 606:57:freechips.rocketchip.system.DefaultRV32Config.fir@12029.4]
  assign _GEN_74 = {{4'd0}, _T_1714}; // @[Monitor.scala 629:97:freechips.rocketchip.system.DefaultRV32Config.fir@12030.4]
  assign _T_1719 = _GEN_74 & _T_1718; // @[Monitor.scala 629:97:freechips.rocketchip.system.DefaultRV32Config.fir@12030.4]
  assign _T_1720 = {{1'd0}, _T_1719[15:1]}; // @[Monitor.scala 629:152:freechips.rocketchip.system.DefaultRV32Config.fir@12031.4]
  assign _T_1721 = {io_in_d_bits_source, 3'h0}; // @[Monitor.scala 633:65:freechips.rocketchip.system.DefaultRV32Config.fir@12035.4]
  assign _T_1722 = inflight_sizes >> _T_1721; // @[Monitor.scala 633:40:freechips.rocketchip.system.DefaultRV32Config.fir@12036.4]
  assign _T_1726 = 16'h100 - 16'h1; // @[Monitor.scala 606:57:freechips.rocketchip.system.DefaultRV32Config.fir@12040.4]
  assign _GEN_76 = {{8'd0}, _T_1726}; // @[Monitor.scala 633:91:freechips.rocketchip.system.DefaultRV32Config.fir@12041.4]
  assign _T_1727 = _T_1722 & _GEN_76; // @[Monitor.scala 633:91:freechips.rocketchip.system.DefaultRV32Config.fir@12041.4]
  assign _T_1728 = {{1'd0}, _T_1727[23:1]}; // @[Monitor.scala 633:144:freechips.rocketchip.system.DefaultRV32Config.fir@12042.4]
  assign _T_1732 = _T_1477 & a_first; // @[Monitor.scala 643:27:freechips.rocketchip.system.DefaultRV32Config.fir@12067.4]
  assign _T_1734 = 4'h1 << io_in_a_bits_source; // @[OneHot.scala 58:35:freechips.rocketchip.system.DefaultRV32Config.fir@12070.6]
  assign _T_1735 = {io_in_a_bits_opcode, 1'h0}; // @[Monitor.scala 645:53:freechips.rocketchip.system.DefaultRV32Config.fir@12072.6]
  assign _T_1736 = _T_1735 | 4'h1; // @[Monitor.scala 645:61:freechips.rocketchip.system.DefaultRV32Config.fir@12073.6]
  assign _T_1737 = {io_in_a_bits_size, 1'h0}; // @[Monitor.scala 646:49:freechips.rocketchip.system.DefaultRV32Config.fir@12075.6]
  assign _T_1738 = _T_1737 | 5'h1; // @[Monitor.scala 646:57:freechips.rocketchip.system.DefaultRV32Config.fir@12076.6]
  assign _GEN_78 = {io_in_a_bits_source, 2'h0}; // @[Monitor.scala 647:72:freechips.rocketchip.system.DefaultRV32Config.fir@12078.6]
  assign _T_1739 = {{1'd0}, _GEN_78}; // @[Monitor.scala 647:72:freechips.rocketchip.system.DefaultRV32Config.fir@12078.6]
  assign a_opcodes_set_interm = _T_1732 ? _T_1736 : 4'h0; // @[Monitor.scala 643:72:freechips.rocketchip.system.DefaultRV32Config.fir@12069.4]
  assign _GEN_79 = {{31'd0}, a_opcodes_set_interm}; // @[Monitor.scala 647:47:freechips.rocketchip.system.DefaultRV32Config.fir@12079.6]
  assign _T_1740 = _GEN_79 << _T_1739; // @[Monitor.scala 647:47:freechips.rocketchip.system.DefaultRV32Config.fir@12079.6]
  assign _T_1741 = {io_in_a_bits_source, 3'h0}; // @[Monitor.scala 648:68:freechips.rocketchip.system.DefaultRV32Config.fir@12081.6]
  assign a_sizes_set_interm = _T_1732 ? _T_1738 : 5'h0; // @[Monitor.scala 643:72:freechips.rocketchip.system.DefaultRV32Config.fir@12069.4]
  assign _GEN_80 = {{31'd0}, a_sizes_set_interm}; // @[Monitor.scala 648:43:freechips.rocketchip.system.DefaultRV32Config.fir@12082.6]
  assign _T_1742 = _GEN_80 << _T_1741; // @[Monitor.scala 648:43:freechips.rocketchip.system.DefaultRV32Config.fir@12082.6]
  assign _T_1743 = inflight >> io_in_a_bits_source; // @[Monitor.scala 649:26:freechips.rocketchip.system.DefaultRV32Config.fir@12084.6]
  assign _T_1745 = ~_T_1743[0]; // @[Monitor.scala 649:17:freechips.rocketchip.system.DefaultRV32Config.fir@12086.6]
  assign _T_1747 = _T_1745 | reset; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@12088.6]
  assign _T_1748 = ~_T_1747; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@12089.6]
  assign _GEN_27 = _T_1732 ? _T_1734 : 4'h0; // @[Monitor.scala 643:72:freechips.rocketchip.system.DefaultRV32Config.fir@12069.4]
  assign _GEN_30 = _T_1732 ? _T_1740 : 35'h0; // @[Monitor.scala 643:72:freechips.rocketchip.system.DefaultRV32Config.fir@12069.4]
  assign _GEN_31 = _T_1732 ? _T_1742 : 36'h0; // @[Monitor.scala 643:72:freechips.rocketchip.system.DefaultRV32Config.fir@12069.4]
  assign _T_1751 = _T_1526 & d_first; // @[Monitor.scala 660:27:freechips.rocketchip.system.DefaultRV32Config.fir@12103.4]
  assign _T_1753 = ~_T_708; // @[Monitor.scala 660:75:freechips.rocketchip.system.DefaultRV32Config.fir@12105.4]
  assign _T_1754 = _T_1751 & _T_1753; // @[Monitor.scala 660:72:freechips.rocketchip.system.DefaultRV32Config.fir@12106.4]
  assign _T_1755 = 4'h1 << io_in_d_bits_source; // @[OneHot.scala 58:35:freechips.rocketchip.system.DefaultRV32Config.fir@12108.6]
  assign _GEN_82 = {{31'd0}, _T_1718}; // @[Monitor.scala 662:76:freechips.rocketchip.system.DefaultRV32Config.fir@12115.6]
  assign _T_1761 = _GEN_82 << _T_1713; // @[Monitor.scala 662:76:freechips.rocketchip.system.DefaultRV32Config.fir@12115.6]
  assign _GEN_83 = {{31'd0}, _T_1726}; // @[Monitor.scala 663:72:freechips.rocketchip.system.DefaultRV32Config.fir@12122.6]
  assign _T_1767 = _GEN_83 << _T_1721; // @[Monitor.scala 663:72:freechips.rocketchip.system.DefaultRV32Config.fir@12122.6]
  assign _GEN_32 = _T_1754 ? _T_1755 : 4'h0; // @[Monitor.scala 660:91:freechips.rocketchip.system.DefaultRV32Config.fir@12107.4]
  assign _GEN_33 = _T_1754 ? _T_1761 : 47'h0; // @[Monitor.scala 660:91:freechips.rocketchip.system.DefaultRV32Config.fir@12107.4]
  assign _GEN_34 = _T_1754 ? _T_1767 : 47'h0; // @[Monitor.scala 660:91:freechips.rocketchip.system.DefaultRV32Config.fir@12107.4]
  assign _T_1768 = io_in_d_valid & d_first; // @[Monitor.scala 665:26:freechips.rocketchip.system.DefaultRV32Config.fir@12125.4]
  assign _T_1771 = _T_1768 & _T_1753; // @[Monitor.scala 665:71:freechips.rocketchip.system.DefaultRV32Config.fir@12128.4]
  assign _T_1772 = inflight >> io_in_d_bits_source; // @[Monitor.scala 666:25:freechips.rocketchip.system.DefaultRV32Config.fir@12130.6]
  assign _T_1774 = io_in_a_bits_source == io_in_d_bits_source; // @[Monitor.scala 666:93:freechips.rocketchip.system.DefaultRV32Config.fir@12132.6]
  assign _T_1775 = io_in_a_valid & _T_1774; // @[Monitor.scala 666:68:freechips.rocketchip.system.DefaultRV32Config.fir@12133.6]
  assign _T_1776 = io_in_a_bits_size == io_in_d_bits_size; // @[Monitor.scala 666:142:freechips.rocketchip.system.DefaultRV32Config.fir@12134.6]
  assign _T_1777 = _T_1775 & _T_1776; // @[Monitor.scala 666:119:freechips.rocketchip.system.DefaultRV32Config.fir@12135.6]
  assign _T_1778 = _T_1777 & a_first; // @[Monitor.scala 666:166:freechips.rocketchip.system.DefaultRV32Config.fir@12136.6]
  assign _T_1779 = _T_1772[0] | _T_1778; // @[Monitor.scala 666:49:freechips.rocketchip.system.DefaultRV32Config.fir@12137.6]
  assign _T_1781 = _T_1779 | reset; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@12139.6]
  assign _T_1782 = ~_T_1781; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@12140.6]
  assign a_opcode_lookup = _T_1720[3:0]; // @[:freechips.rocketchip.system.DefaultRV32Config.fir@12022.4 :freechips.rocketchip.system.DefaultRV32Config.fir@12023.4 Monitor.scala 629:21:freechips.rocketchip.system.DefaultRV32Config.fir@12032.4]
  assign _GEN_37 = 3'h2 == a_opcode_lookup[2:0] ? 3'h1 : 3'h0; // @[Monitor.scala 667:37:freechips.rocketchip.system.DefaultRV32Config.fir@12146.6]
  assign _GEN_38 = 3'h3 == a_opcode_lookup[2:0] ? 3'h1 : _GEN_37; // @[Monitor.scala 667:37:freechips.rocketchip.system.DefaultRV32Config.fir@12146.6]
  assign _GEN_39 = 3'h4 == a_opcode_lookup[2:0] ? 3'h1 : _GEN_38; // @[Monitor.scala 667:37:freechips.rocketchip.system.DefaultRV32Config.fir@12146.6]
  assign _GEN_40 = 3'h5 == a_opcode_lookup[2:0] ? 3'h2 : _GEN_39; // @[Monitor.scala 667:37:freechips.rocketchip.system.DefaultRV32Config.fir@12146.6]
  assign _GEN_41 = 3'h6 == a_opcode_lookup[2:0] ? 3'h4 : _GEN_40; // @[Monitor.scala 667:37:freechips.rocketchip.system.DefaultRV32Config.fir@12146.6]
  assign _GEN_42 = 3'h7 == a_opcode_lookup[2:0] ? 3'h4 : _GEN_41; // @[Monitor.scala 667:37:freechips.rocketchip.system.DefaultRV32Config.fir@12146.6]
  assign _T_1784 = io_in_d_bits_opcode == _GEN_42; // @[Monitor.scala 667:37:freechips.rocketchip.system.DefaultRV32Config.fir@12146.6]
  assign _GEN_49 = 3'h6 == a_opcode_lookup[2:0] ? 3'h5 : _GEN_40; // @[Monitor.scala 667:96:freechips.rocketchip.system.DefaultRV32Config.fir@12148.6]
  assign _GEN_50 = 3'h7 == a_opcode_lookup[2:0] ? 3'h4 : _GEN_49; // @[Monitor.scala 667:96:freechips.rocketchip.system.DefaultRV32Config.fir@12148.6]
  assign _T_1786 = io_in_d_bits_opcode == _GEN_50; // @[Monitor.scala 667:96:freechips.rocketchip.system.DefaultRV32Config.fir@12148.6]
  assign _T_1787 = _T_1784 | _T_1786; // @[Monitor.scala 667:71:freechips.rocketchip.system.DefaultRV32Config.fir@12149.6]
  assign _GEN_53 = 3'h2 == io_in_a_bits_opcode ? 3'h1 : 3'h0; // @[Monitor.scala 668:60:freechips.rocketchip.system.DefaultRV32Config.fir@12150.6]
  assign _GEN_54 = 3'h3 == io_in_a_bits_opcode ? 3'h1 : _GEN_53; // @[Monitor.scala 668:60:freechips.rocketchip.system.DefaultRV32Config.fir@12150.6]
  assign _GEN_55 = 3'h4 == io_in_a_bits_opcode ? 3'h1 : _GEN_54; // @[Monitor.scala 668:60:freechips.rocketchip.system.DefaultRV32Config.fir@12150.6]
  assign _GEN_56 = 3'h5 == io_in_a_bits_opcode ? 3'h2 : _GEN_55; // @[Monitor.scala 668:60:freechips.rocketchip.system.DefaultRV32Config.fir@12150.6]
  assign _GEN_57 = 3'h6 == io_in_a_bits_opcode ? 3'h4 : _GEN_56; // @[Monitor.scala 668:60:freechips.rocketchip.system.DefaultRV32Config.fir@12150.6]
  assign _GEN_58 = 3'h7 == io_in_a_bits_opcode ? 3'h4 : _GEN_57; // @[Monitor.scala 668:60:freechips.rocketchip.system.DefaultRV32Config.fir@12150.6]
  assign _T_1788 = io_in_d_bits_opcode == _GEN_58; // @[Monitor.scala 668:60:freechips.rocketchip.system.DefaultRV32Config.fir@12150.6]
  assign _GEN_65 = 3'h6 == io_in_a_bits_opcode ? 3'h5 : _GEN_56; // @[Monitor.scala 668:124:freechips.rocketchip.system.DefaultRV32Config.fir@12151.6]
  assign _GEN_66 = 3'h7 == io_in_a_bits_opcode ? 3'h4 : _GEN_65; // @[Monitor.scala 668:124:freechips.rocketchip.system.DefaultRV32Config.fir@12151.6]
  assign _T_1789 = io_in_d_bits_opcode == _GEN_66; // @[Monitor.scala 668:124:freechips.rocketchip.system.DefaultRV32Config.fir@12151.6]
  assign _T_1790 = _T_1788 | _T_1789; // @[Monitor.scala 668:99:freechips.rocketchip.system.DefaultRV32Config.fir@12152.6]
  assign _T_1791 = io_in_a_valid & _T_1790; // @[Monitor.scala 668:34:freechips.rocketchip.system.DefaultRV32Config.fir@12153.6]
  assign _T_1792 = _T_1787 | _T_1791; // @[Monitor.scala 668:15:freechips.rocketchip.system.DefaultRV32Config.fir@12154.6]
  assign _T_1794 = _T_1792 | reset; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@12156.6]
  assign _T_1795 = ~_T_1794; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@12157.6]
  assign a_size_lookup = _T_1728[7:0]; // @[:freechips.rocketchip.system.DefaultRV32Config.fir@12033.4 :freechips.rocketchip.system.DefaultRV32Config.fir@12034.4 Monitor.scala 633:19:freechips.rocketchip.system.DefaultRV32Config.fir@12043.4]
  assign _GEN_84 = {{4'd0}, io_in_d_bits_size}; // @[Monitor.scala 670:34:freechips.rocketchip.system.DefaultRV32Config.fir@12162.6]
  assign _T_1796 = _GEN_84 == a_size_lookup; // @[Monitor.scala 670:34:freechips.rocketchip.system.DefaultRV32Config.fir@12162.6]
  assign _T_1798 = io_in_a_valid & _T_1776; // @[Monitor.scala 670:72:freechips.rocketchip.system.DefaultRV32Config.fir@12164.6]
  assign _T_1799 = _T_1796 | _T_1798; // @[Monitor.scala 670:53:freechips.rocketchip.system.DefaultRV32Config.fir@12165.6]
  assign _T_1801 = _T_1799 | reset; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@12167.6]
  assign _T_1802 = ~_T_1801; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@12168.6]
  assign _T_1804 = _T_1768 & a_first; // @[Monitor.scala 672:36:freechips.rocketchip.system.DefaultRV32Config.fir@12175.4]
  assign _T_1805 = _T_1804 & io_in_a_valid; // @[Monitor.scala 672:47:freechips.rocketchip.system.DefaultRV32Config.fir@12176.4]
  assign _T_1807 = _T_1805 & _T_1774; // @[Monitor.scala 672:65:freechips.rocketchip.system.DefaultRV32Config.fir@12178.4]
  assign _T_1809 = _T_1807 & _T_1753; // @[Monitor.scala 672:116:freechips.rocketchip.system.DefaultRV32Config.fir@12180.4]
  assign _T_1810 = ~io_in_d_ready; // @[Monitor.scala 673:15:freechips.rocketchip.system.DefaultRV32Config.fir@12182.6]
  assign _T_1811 = _T_1810 | io_in_a_ready; // @[Monitor.scala 673:32:freechips.rocketchip.system.DefaultRV32Config.fir@12183.6]
  assign _T_1813 = _T_1811 | reset; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@12185.6]
  assign _T_1814 = ~_T_1813; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@12186.6]
  assign a_set = _GEN_27[2:0]; // @[:freechips.rocketchip.system.DefaultRV32Config.fir@12016.4 :freechips.rocketchip.system.DefaultRV32Config.fir@12017.4 Monitor.scala 644:13:freechips.rocketchip.system.DefaultRV32Config.fir@12071.6]
  assign d_clr = _GEN_32[2:0]; // @[:freechips.rocketchip.system.DefaultRV32Config.fir@12095.4 :freechips.rocketchip.system.DefaultRV32Config.fir@12096.4 Monitor.scala 661:13:freechips.rocketchip.system.DefaultRV32Config.fir@12109.6]
  assign _T_1815 = a_set != d_clr; // @[Monitor.scala 677:20:freechips.rocketchip.system.DefaultRV32Config.fir@12192.4]
  assign _T_1816 = |a_set; // @[Monitor.scala 677:40:freechips.rocketchip.system.DefaultRV32Config.fir@12193.4]
  assign _T_1817 = ~_T_1816; // @[Monitor.scala 677:33:freechips.rocketchip.system.DefaultRV32Config.fir@12194.4]
  assign _T_1818 = _T_1815 | _T_1817; // @[Monitor.scala 677:30:freechips.rocketchip.system.DefaultRV32Config.fir@12195.4]
  assign _T_1820 = _T_1818 | reset; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@12197.4]
  assign _T_1821 = ~_T_1820; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@12198.4]
  assign _T_1822 = inflight | a_set; // @[Monitor.scala 680:27:freechips.rocketchip.system.DefaultRV32Config.fir@12203.4]
  assign _T_1823 = ~d_clr; // @[Monitor.scala 680:38:freechips.rocketchip.system.DefaultRV32Config.fir@12204.4]
  assign _T_1824 = _T_1822 & _T_1823; // @[Monitor.scala 680:36:freechips.rocketchip.system.DefaultRV32Config.fir@12205.4]
  assign a_opcodes_set = _GEN_30[11:0]; // @[:freechips.rocketchip.system.DefaultRV32Config.fir@12018.4 :freechips.rocketchip.system.DefaultRV32Config.fir@12019.4 Monitor.scala 647:21:freechips.rocketchip.system.DefaultRV32Config.fir@12080.6]
  assign _T_1825 = inflight_opcodes | a_opcodes_set; // @[Monitor.scala 681:43:freechips.rocketchip.system.DefaultRV32Config.fir@12207.4]
  assign d_opcodes_clr = _GEN_33[11:0]; // @[:freechips.rocketchip.system.DefaultRV32Config.fir@12097.4 :freechips.rocketchip.system.DefaultRV32Config.fir@12098.4 Monitor.scala 662:21:freechips.rocketchip.system.DefaultRV32Config.fir@12116.6]
  assign _T_1826 = ~d_opcodes_clr; // @[Monitor.scala 681:62:freechips.rocketchip.system.DefaultRV32Config.fir@12208.4]
  assign _T_1827 = _T_1825 & _T_1826; // @[Monitor.scala 681:60:freechips.rocketchip.system.DefaultRV32Config.fir@12209.4]
  assign a_sizes_set = _GEN_31[23:0]; // @[:freechips.rocketchip.system.DefaultRV32Config.fir@12020.4 :freechips.rocketchip.system.DefaultRV32Config.fir@12021.4 Monitor.scala 648:19:freechips.rocketchip.system.DefaultRV32Config.fir@12083.6]
  assign _T_1828 = inflight_sizes | a_sizes_set; // @[Monitor.scala 682:39:freechips.rocketchip.system.DefaultRV32Config.fir@12211.4]
  assign d_sizes_clr = _GEN_34[23:0]; // @[:freechips.rocketchip.system.DefaultRV32Config.fir@12099.4 :freechips.rocketchip.system.DefaultRV32Config.fir@12100.4 Monitor.scala 663:19:freechips.rocketchip.system.DefaultRV32Config.fir@12123.6]
  assign _T_1829 = ~d_sizes_clr; // @[Monitor.scala 682:56:freechips.rocketchip.system.DefaultRV32Config.fir@12212.4]
  assign _T_1830 = _T_1828 & _T_1829; // @[Monitor.scala 682:54:freechips.rocketchip.system.DefaultRV32Config.fir@12213.4]
  assign _T_1832 = |inflight; // @[Monitor.scala 687:26:freechips.rocketchip.system.DefaultRV32Config.fir@12218.4]
  assign _T_1833 = ~_T_1832; // @[Monitor.scala 687:16:freechips.rocketchip.system.DefaultRV32Config.fir@12219.4]
  assign _T_1834 = plusarg_reader_out == 32'h0; // @[Monitor.scala 687:39:freechips.rocketchip.system.DefaultRV32Config.fir@12220.4]
  assign _T_1835 = _T_1833 | _T_1834; // @[Monitor.scala 687:30:freechips.rocketchip.system.DefaultRV32Config.fir@12221.4]
  assign _T_1836 = _T_1831 < plusarg_reader_out; // @[Monitor.scala 687:59:freechips.rocketchip.system.DefaultRV32Config.fir@12222.4]
  assign _T_1837 = _T_1835 | _T_1836; // @[Monitor.scala 687:47:freechips.rocketchip.system.DefaultRV32Config.fir@12223.4]
  assign _T_1839 = _T_1837 | reset; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@12225.4]
  assign _T_1840 = ~_T_1839; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@12226.4]
  assign _T_1842 = _T_1831 + 32'h1; // @[Monitor.scala 689:26:freechips.rocketchip.system.DefaultRV32Config.fir@12232.4]
  assign _T_1845 = _T_1477 | _T_1526; // @[Monitor.scala 690:27:freechips.rocketchip.system.DefaultRV32Config.fir@12236.4]
  assign _T_1857 = _T_1855 - 10'h1; // @[Edges.scala 231:28:freechips.rocketchip.system.DefaultRV32Config.fir@12251.4]
  assign _T_1858 = _T_1855 == 10'h0; // @[Edges.scala 232:25:freechips.rocketchip.system.DefaultRV32Config.fir@12252.4]
  assign _T_1868 = _T_1526 & _T_1858; // @[Monitor.scala 700:27:freechips.rocketchip.system.DefaultRV32Config.fir@12266.4]
  assign _T_1871 = ~io_in_d_bits_opcode[1]; // @[Edges.scala 72:43:freechips.rocketchip.system.DefaultRV32Config.fir@12269.4]
  assign _T_1872 = io_in_d_bits_opcode[2] & _T_1871; // @[Edges.scala 72:40:freechips.rocketchip.system.DefaultRV32Config.fir@12270.4]
  assign _T_1873 = _T_1868 & _T_1872; // @[Monitor.scala 700:38:freechips.rocketchip.system.DefaultRV32Config.fir@12271.4]
  assign _T_1874 = 4'h1 << io_in_d_bits_sink; // @[OneHot.scala 58:35:freechips.rocketchip.system.DefaultRV32Config.fir@12273.6]
  assign _T_1875 = _T_1846 >> io_in_d_bits_sink; // @[Monitor.scala 702:23:freechips.rocketchip.system.DefaultRV32Config.fir@12275.6]
  assign _T_1877 = ~_T_1875[0]; // @[Monitor.scala 702:14:freechips.rocketchip.system.DefaultRV32Config.fir@12277.6]
  assign _T_1879 = _T_1877 | reset; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@12279.6]
  assign _T_1880 = ~_T_1879; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@12280.6]
  assign _GEN_69 = _T_1873 ? _T_1874 : 4'h0; // @[Monitor.scala 700:72:freechips.rocketchip.system.DefaultRV32Config.fir@12272.4]
  assign _T_1885 = 4'h1 << io_in_e_bits_sink; // @[OneHot.scala 58:35:freechips.rocketchip.system.DefaultRV32Config.fir@12292.6]
  assign _T_1886 = _GEN_69 | _T_1846; // @[Monitor.scala 708:24:freechips.rocketchip.system.DefaultRV32Config.fir@12294.6]
  assign _T_1887 = _T_1886 >> io_in_e_bits_sink; // @[Monitor.scala 708:35:freechips.rocketchip.system.DefaultRV32Config.fir@12295.6]
  assign _T_1890 = _T_1887[0] | reset; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@12298.6]
  assign _T_1891 = ~_T_1890; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@12299.6]
  assign _GEN_70 = io_in_e_valid ? _T_1885 : 4'h0; // @[Monitor.scala 706:73:freechips.rocketchip.system.DefaultRV32Config.fir@12291.4]
  assign _T_1892 = _T_1846 | _GEN_69; // @[Monitor.scala 713:27:freechips.rocketchip.system.DefaultRV32Config.fir@12305.4]
  assign _T_1893 = ~_GEN_70; // @[Monitor.scala 713:38:freechips.rocketchip.system.DefaultRV32Config.fir@12306.4]
  assign _T_1894 = _T_1892 & _T_1893; // @[Monitor.scala 713:36:freechips.rocketchip.system.DefaultRV32Config.fir@12307.4]
  assign _GEN_85 = io_in_a_valid & _T_78; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@9501.10]
  assign _GEN_101 = io_in_a_valid & _T_168; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@9630.10]
  assign _GEN_119 = io_in_a_valid & _T_262; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@9770.10]
  assign _GEN_131 = io_in_a_valid & _T_336; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@9877.10]
  assign _GEN_141 = io_in_a_valid & _T_413; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@9976.10]
  assign _GEN_151 = io_in_a_valid & _T_492; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@10067.10]
  assign _GEN_161 = io_in_a_valid & _T_559; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@10156.10]
  assign _GEN_171 = io_in_a_valid & _T_626; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@10245.10]
  assign _GEN_183 = io_in_d_valid & _T_708; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@10314.10]
  assign _GEN_193 = io_in_d_valid & _T_728; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@10356.10]
  assign _GEN_203 = io_in_d_valid & _T_756; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@10414.10]
  assign _GEN_213 = io_in_d_valid & _T_785; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@10473.10]
  assign _GEN_219 = io_in_d_valid & _T_802; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@10508.10]
  assign _GEN_225 = io_in_d_valid & _T_820; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@10544.10]
  assign _GEN_231 = io_in_c_valid & _T_1217; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@11199.10]
  assign _GEN_243 = io_in_c_valid & _T_1239; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@11247.10]
  assign _GEN_253 = io_in_c_valid & _T_1257; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@11336.10]
  assign _GEN_267 = io_in_c_valid & _T_1342; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@11456.10]
  assign _GEN_279 = io_in_c_valid & _T_1423; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@11519.10]
  assign _GEN_289 = io_in_c_valid & _T_1441; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@11559.10]
  assign _GEN_297 = io_in_c_valid & _T_1455; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@11591.10]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_1486 = _RAND_0[9:0];
  _RAND_1 = {1{`RANDOM}};
  _T_1497 = _RAND_1[2:0];
  _RAND_2 = {1{`RANDOM}};
  _T_1498 = _RAND_2[2:0];
  _RAND_3 = {1{`RANDOM}};
  _T_1499 = _RAND_3[3:0];
  _RAND_4 = {1{`RANDOM}};
  _T_1500 = _RAND_4[1:0];
  _RAND_5 = {1{`RANDOM}};
  _T_1501 = _RAND_5[31:0];
  _RAND_6 = {1{`RANDOM}};
  _T_1534 = _RAND_6[9:0];
  _RAND_7 = {1{`RANDOM}};
  _T_1545 = _RAND_7[2:0];
  _RAND_8 = {1{`RANDOM}};
  _T_1546 = _RAND_8[1:0];
  _RAND_9 = {1{`RANDOM}};
  _T_1547 = _RAND_9[3:0];
  _RAND_10 = {1{`RANDOM}};
  _T_1548 = _RAND_10[1:0];
  _RAND_11 = {1{`RANDOM}};
  _T_1549 = _RAND_11[1:0];
  _RAND_12 = {1{`RANDOM}};
  _T_1550 = _RAND_12[0:0];
  _RAND_13 = {1{`RANDOM}};
  _T_1588 = _RAND_13[9:0];
  _RAND_14 = {1{`RANDOM}};
  _T_1600 = _RAND_14[1:0];
  _RAND_15 = {1{`RANDOM}};
  _T_1603 = _RAND_15[31:0];
  _RAND_16 = {1{`RANDOM}};
  _T_1636 = _RAND_16[9:0];
  _RAND_17 = {1{`RANDOM}};
  _T_1647 = _RAND_17[2:0];
  _RAND_18 = {1{`RANDOM}};
  _T_1648 = _RAND_18[2:0];
  _RAND_19 = {1{`RANDOM}};
  _T_1649 = _RAND_19[3:0];
  _RAND_20 = {1{`RANDOM}};
  _T_1650 = _RAND_20[1:0];
  _RAND_21 = {1{`RANDOM}};
  _T_1651 = _RAND_21[31:0];
  _RAND_22 = {1{`RANDOM}};
  inflight = _RAND_22[2:0];
  _RAND_23 = {1{`RANDOM}};
  inflight_opcodes = _RAND_23[11:0];
  _RAND_24 = {1{`RANDOM}};
  inflight_sizes = _RAND_24[23:0];
  _RAND_25 = {1{`RANDOM}};
  _T_1685 = _RAND_25[9:0];
  _RAND_26 = {1{`RANDOM}};
  _T_1703 = _RAND_26[9:0];
  _RAND_27 = {1{`RANDOM}};
  _T_1831 = _RAND_27[31:0];
  _RAND_28 = {1{`RANDOM}};
  _T_1846 = _RAND_28[3:0];
  _RAND_29 = {1{`RANDOM}};
  _T_1855 = _RAND_29[9:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      _T_1486 <= 10'h0;
    end else if (_T_1477) begin
      if (_T_1489) begin
        if (_T_1484) begin
          _T_1486 <= _T_13[11:2];
        end else begin
          _T_1486 <= 10'h0;
        end
      end else begin
        _T_1486 <= _T_1488;
      end
    end
    if (_T_1525) begin
      _T_1497 <= io_in_a_bits_opcode;
    end
    if (_T_1525) begin
      _T_1498 <= io_in_a_bits_param;
    end
    if (_T_1525) begin
      _T_1499 <= io_in_a_bits_size;
    end
    if (_T_1525) begin
      _T_1500 <= io_in_a_bits_source;
    end
    if (_T_1525) begin
      _T_1501 <= io_in_a_bits_address;
    end
    if (reset) begin
      _T_1534 <= 10'h0;
    end else if (_T_1526) begin
      if (_T_1537) begin
        if (io_in_d_bits_opcode[0]) begin
          _T_1534 <= _T_1530[11:2];
        end else begin
          _T_1534 <= 10'h0;
        end
      end else begin
        _T_1534 <= _T_1536;
      end
    end
    if (_T_1578) begin
      _T_1545 <= io_in_d_bits_opcode;
    end
    if (_T_1578) begin
      _T_1546 <= io_in_d_bits_param;
    end
    if (_T_1578) begin
      _T_1547 <= io_in_d_bits_size;
    end
    if (_T_1578) begin
      _T_1548 <= io_in_d_bits_source;
    end
    if (_T_1578) begin
      _T_1549 <= io_in_d_bits_sink;
    end
    if (_T_1578) begin
      _T_1550 <= io_in_d_bits_denied;
    end
    if (reset) begin
      _T_1588 <= 10'h0;
    end else if (_T_1579) begin
      if (_T_1591) begin
        _T_1588 <= 10'h0;
      end else begin
        _T_1588 <= _T_1590;
      end
    end
    if (_T_1627) begin
      _T_1600 <= io_in_b_bits_param;
    end
    if (_T_1627) begin
      _T_1603 <= io_in_b_bits_address;
    end
    if (reset) begin
      _T_1636 <= 10'h0;
    end else if (_T_1628) begin
      if (_T_1639) begin
        if (io_in_c_bits_opcode[0]) begin
          _T_1636 <= _T_1143[11:2];
        end else begin
          _T_1636 <= 10'h0;
        end
      end else begin
        _T_1636 <= _T_1638;
      end
    end
    if (_T_1675) begin
      _T_1647 <= io_in_c_bits_opcode;
    end
    if (_T_1675) begin
      _T_1648 <= io_in_c_bits_param;
    end
    if (_T_1675) begin
      _T_1649 <= io_in_c_bits_size;
    end
    if (_T_1675) begin
      _T_1650 <= io_in_c_bits_source;
    end
    if (_T_1675) begin
      _T_1651 <= io_in_c_bits_address;
    end
    if (reset) begin
      inflight <= 3'h0;
    end else begin
      inflight <= _T_1824;
    end
    if (reset) begin
      inflight_opcodes <= 12'h0;
    end else begin
      inflight_opcodes <= _T_1827;
    end
    if (reset) begin
      inflight_sizes <= 24'h0;
    end else begin
      inflight_sizes <= _T_1830;
    end
    if (reset) begin
      _T_1685 <= 10'h0;
    end else if (_T_1477) begin
      if (a_first) begin
        if (_T_1484) begin
          _T_1685 <= _T_13[11:2];
        end else begin
          _T_1685 <= 10'h0;
        end
      end else begin
        _T_1685 <= _T_1687;
      end
    end
    if (reset) begin
      _T_1703 <= 10'h0;
    end else if (_T_1526) begin
      if (d_first) begin
        if (io_in_d_bits_opcode[0]) begin
          _T_1703 <= _T_1530[11:2];
        end else begin
          _T_1703 <= 10'h0;
        end
      end else begin
        _T_1703 <= _T_1705;
      end
    end
    if (reset) begin
      _T_1831 <= 32'h0;
    end else if (_T_1845) begin
      _T_1831 <= 32'h0;
    end else begin
      _T_1831 <= _T_1842;
    end
    if (reset) begin
      _T_1846 <= 4'h0;
    end else begin
      _T_1846 <= _T_1894;
    end
    if (reset) begin
      _T_1855 <= 10'h0;
    end else if (_T_1526) begin
      if (_T_1858) begin
        if (io_in_d_bits_opcode[0]) begin
          _T_1855 <= _T_1530[11:2];
        end else begin
          _T_1855 <= 10'h0;
        end
      end else begin
        _T_1855 <= _T_1857;
      end
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_85 & _T_130) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel carries AcquireBlock type unsupported by manager (connected at SystemBus.scala:39:96)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@9501.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_85 & _T_130) begin
          $fatal; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@9502.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_85 & _T_144) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel carries AcquireBlock from a client which does not support Probe (connected at SystemBus.scala:39:96)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@9524.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_85 & _T_144) begin
          $fatal; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@9525.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_85 & _T_147) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel AcquireBlock carries invalid source ID (connected at SystemBus.scala:39:96)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@9531.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_85 & _T_147) begin
          $fatal; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@9532.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_85 & _T_151) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel AcquireBlock smaller than a beat (connected at SystemBus.scala:39:96)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@9539.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_85 & _T_151) begin
          $fatal; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@9540.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_85 & _T_154) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel AcquireBlock address not aligned to size (connected at SystemBus.scala:39:96)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@9546.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_85 & _T_154) begin
          $fatal; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@9547.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_85 & _T_158) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel AcquireBlock carries invalid grow param (connected at SystemBus.scala:39:96)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@9554.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_85 & _T_158) begin
          $fatal; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@9555.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_85 & _T_163) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel AcquireBlock contains invalid mask (connected at SystemBus.scala:39:96)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@9563.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_85 & _T_163) begin
          $fatal; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@9564.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_85 & _T_167) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel AcquireBlock is corrupt (connected at SystemBus.scala:39:96)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@9571.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_85 & _T_167) begin
          $fatal; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@9572.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_101 & _T_130) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel carries AcquirePerm type unsupported by manager (connected at SystemBus.scala:39:96)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@9630.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_101 & _T_130) begin
          $fatal; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@9631.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_101 & _T_144) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel carries AcquirePerm from a client which does not support Probe (connected at SystemBus.scala:39:96)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@9653.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_101 & _T_144) begin
          $fatal; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@9654.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_101 & _T_147) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel AcquirePerm carries invalid source ID (connected at SystemBus.scala:39:96)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@9660.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_101 & _T_147) begin
          $fatal; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@9661.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_101 & _T_151) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel AcquirePerm smaller than a beat (connected at SystemBus.scala:39:96)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@9668.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_101 & _T_151) begin
          $fatal; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@9669.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_101 & _T_154) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel AcquirePerm address not aligned to size (connected at SystemBus.scala:39:96)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@9675.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_101 & _T_154) begin
          $fatal; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@9676.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_101 & _T_158) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel AcquirePerm carries invalid grow param (connected at SystemBus.scala:39:96)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@9683.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_101 & _T_158) begin
          $fatal; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@9684.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_101 & _T_252) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel AcquirePerm requests NtoB (connected at SystemBus.scala:39:96)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@9691.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_101 & _T_252) begin
          $fatal; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@9692.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_101 & _T_163) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel AcquirePerm contains invalid mask (connected at SystemBus.scala:39:96)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@9700.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_101 & _T_163) begin
          $fatal; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@9701.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_101 & _T_167) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel AcquirePerm is corrupt (connected at SystemBus.scala:39:96)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@9708.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_101 & _T_167) begin
          $fatal; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@9709.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_119 & _T_317) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel carries Get type unsupported by manager (connected at SystemBus.scala:39:96)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@9770.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_119 & _T_317) begin
          $fatal; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@9771.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_119 & _T_147) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel Get carries invalid source ID (connected at SystemBus.scala:39:96)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@9777.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_119 & _T_147) begin
          $fatal; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@9778.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_119 & _T_154) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel Get address not aligned to size (connected at SystemBus.scala:39:96)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@9784.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_119 & _T_154) begin
          $fatal; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@9785.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_119 & _T_327) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel Get carries invalid param (connected at SystemBus.scala:39:96)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@9792.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_119 & _T_327) begin
          $fatal; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@9793.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_119 & _T_331) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel Get contains invalid mask (connected at SystemBus.scala:39:96)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@9800.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_119 & _T_331) begin
          $fatal; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@9801.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_119 & _T_167) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel Get is corrupt (connected at SystemBus.scala:39:96)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@9808.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_119 & _T_167) begin
          $fatal; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@9809.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_131 & _T_398) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel carries PutFull type unsupported by manager (connected at SystemBus.scala:39:96)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@9877.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_131 & _T_398) begin
          $fatal; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@9878.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_131 & _T_147) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel PutFull carries invalid source ID (connected at SystemBus.scala:39:96)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@9884.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_131 & _T_147) begin
          $fatal; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@9885.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_131 & _T_154) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel PutFull address not aligned to size (connected at SystemBus.scala:39:96)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@9891.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_131 & _T_154) begin
          $fatal; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@9892.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_131 & _T_327) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel PutFull carries invalid param (connected at SystemBus.scala:39:96)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@9899.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_131 & _T_327) begin
          $fatal; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@9900.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_131 & _T_331) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel PutFull contains invalid mask (connected at SystemBus.scala:39:96)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@9907.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_131 & _T_331) begin
          $fatal; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@9908.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_141 & _T_398) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel carries PutPartial type unsupported by manager (connected at SystemBus.scala:39:96)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@9976.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_141 & _T_398) begin
          $fatal; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@9977.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_141 & _T_147) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel PutPartial carries invalid source ID (connected at SystemBus.scala:39:96)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@9983.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_141 & _T_147) begin
          $fatal; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@9984.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_141 & _T_154) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel PutPartial address not aligned to size (connected at SystemBus.scala:39:96)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@9990.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_141 & _T_154) begin
          $fatal; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@9991.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_141 & _T_327) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel PutPartial carries invalid param (connected at SystemBus.scala:39:96)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@9998.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_141 & _T_327) begin
          $fatal; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@9999.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_141 & _T_491) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel PutPartial contains invalid mask (connected at SystemBus.scala:39:96)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@10008.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_141 & _T_491) begin
          $fatal; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@10009.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_151 & _T_544) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel carries Arithmetic type unsupported by manager (connected at SystemBus.scala:39:96)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@10067.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_151 & _T_544) begin
          $fatal; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@10068.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_151 & _T_147) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel Arithmetic carries invalid source ID (connected at SystemBus.scala:39:96)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@10074.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_151 & _T_147) begin
          $fatal; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@10075.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_151 & _T_154) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel Arithmetic address not aligned to size (connected at SystemBus.scala:39:96)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@10081.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_151 & _T_154) begin
          $fatal; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@10082.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_151 & _T_554) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel Arithmetic carries invalid opcode param (connected at SystemBus.scala:39:96)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@10089.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_151 & _T_554) begin
          $fatal; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@10090.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_151 & _T_331) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel Arithmetic contains invalid mask (connected at SystemBus.scala:39:96)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@10097.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_151 & _T_331) begin
          $fatal; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@10098.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_161 & _T_544) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel carries Logical type unsupported by manager (connected at SystemBus.scala:39:96)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@10156.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_161 & _T_544) begin
          $fatal; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@10157.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_161 & _T_147) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel Logical carries invalid source ID (connected at SystemBus.scala:39:96)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@10163.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_161 & _T_147) begin
          $fatal; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@10164.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_161 & _T_154) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel Logical address not aligned to size (connected at SystemBus.scala:39:96)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@10170.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_161 & _T_154) begin
          $fatal; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@10171.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_161 & _T_621) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel Logical carries invalid opcode param (connected at SystemBus.scala:39:96)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@10178.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_161 & _T_621) begin
          $fatal; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@10179.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_161 & _T_331) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel Logical contains invalid mask (connected at SystemBus.scala:39:96)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@10186.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_161 & _T_331) begin
          $fatal; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@10187.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_171 & _T_678) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel carries Hint type unsupported by manager (connected at SystemBus.scala:39:96)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@10245.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_171 & _T_678) begin
          $fatal; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@10246.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_171 & _T_147) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel Hint carries invalid source ID (connected at SystemBus.scala:39:96)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@10252.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_171 & _T_147) begin
          $fatal; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@10253.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_171 & _T_154) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel Hint address not aligned to size (connected at SystemBus.scala:39:96)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@10259.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_171 & _T_154) begin
          $fatal; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@10260.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_171 & _T_688) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel Hint carries invalid opcode param (connected at SystemBus.scala:39:96)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@10267.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_171 & _T_688) begin
          $fatal; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@10268.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_171 & _T_331) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel Hint contains invalid mask (connected at SystemBus.scala:39:96)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@10275.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_171 & _T_331) begin
          $fatal; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@10276.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_171 & _T_167) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel Hint is corrupt (connected at SystemBus.scala:39:96)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@10283.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_171 & _T_167) begin
          $fatal; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@10284.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_d_valid & _T_700) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel has invalid opcode (connected at SystemBus.scala:39:96)\n    at Monitor.scala:51 assert(cond, message)\n"); // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@10294.8]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_d_valid & _T_700) begin
          $fatal; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@10295.8]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_183 & _T_711) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel ReleaseAck carries invalid source ID (connected at SystemBus.scala:39:96)\n    at Monitor.scala:51 assert(cond, message)\n"); // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@10314.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_183 & _T_711) begin
          $fatal; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@10315.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_183 & _T_715) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel ReleaseAck smaller than a beat (connected at SystemBus.scala:39:96)\n    at Monitor.scala:51 assert(cond, message)\n"); // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@10322.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_183 & _T_715) begin
          $fatal; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@10323.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_183 & _T_719) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel ReleaseeAck carries invalid param (connected at SystemBus.scala:39:96)\n    at Monitor.scala:51 assert(cond, message)\n"); // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@10330.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_183 & _T_719) begin
          $fatal; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@10331.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_183 & _T_723) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel ReleaseAck is corrupt (connected at SystemBus.scala:39:96)\n    at Monitor.scala:51 assert(cond, message)\n"); // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@10338.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_183 & _T_723) begin
          $fatal; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@10339.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_183 & _T_727) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel ReleaseAck is denied (connected at SystemBus.scala:39:96)\n    at Monitor.scala:51 assert(cond, message)\n"); // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@10346.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_183 & _T_727) begin
          $fatal; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@10347.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_193 & _T_711) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel Grant carries invalid source ID (connected at SystemBus.scala:39:96)\n    at Monitor.scala:51 assert(cond, message)\n"); // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@10356.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_193 & _T_711) begin
          $fatal; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@10357.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_193 & _T_715) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel Grant smaller than a beat (connected at SystemBus.scala:39:96)\n    at Monitor.scala:51 assert(cond, message)\n"); // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@10371.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_193 & _T_715) begin
          $fatal; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@10372.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_193 & _T_742) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel Grant carries invalid cap param (connected at SystemBus.scala:39:96)\n    at Monitor.scala:51 assert(cond, message)\n"); // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@10379.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_193 & _T_742) begin
          $fatal; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@10380.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_193 & _T_746) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel Grant carries toN param (connected at SystemBus.scala:39:96)\n    at Monitor.scala:51 assert(cond, message)\n"); // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@10387.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_193 & _T_746) begin
          $fatal; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@10388.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_193 & _T_723) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel Grant is corrupt (connected at SystemBus.scala:39:96)\n    at Monitor.scala:51 assert(cond, message)\n"); // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@10395.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_193 & _T_723) begin
          $fatal; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@10396.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_203 & _T_711) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel GrantData carries invalid source ID (connected at SystemBus.scala:39:96)\n    at Monitor.scala:51 assert(cond, message)\n"); // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@10414.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_203 & _T_711) begin
          $fatal; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@10415.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_203 & _T_715) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel GrantData smaller than a beat (connected at SystemBus.scala:39:96)\n    at Monitor.scala:51 assert(cond, message)\n"); // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@10429.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_203 & _T_715) begin
          $fatal; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@10430.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_203 & _T_742) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel GrantData carries invalid cap param (connected at SystemBus.scala:39:96)\n    at Monitor.scala:51 assert(cond, message)\n"); // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@10437.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_203 & _T_742) begin
          $fatal; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@10438.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_203 & _T_746) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel GrantData carries toN param (connected at SystemBus.scala:39:96)\n    at Monitor.scala:51 assert(cond, message)\n"); // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@10445.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_203 & _T_746) begin
          $fatal; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@10446.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_203 & _T_779) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel GrantData is denied but not corrupt (connected at SystemBus.scala:39:96)\n    at Monitor.scala:51 assert(cond, message)\n"); // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@10454.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_203 & _T_779) begin
          $fatal; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@10455.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_213 & _T_711) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel AccessAck carries invalid source ID (connected at SystemBus.scala:39:96)\n    at Monitor.scala:51 assert(cond, message)\n"); // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@10473.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_213 & _T_711) begin
          $fatal; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@10474.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_213 & _T_719) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel AccessAck carries invalid param (connected at SystemBus.scala:39:96)\n    at Monitor.scala:51 assert(cond, message)\n"); // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@10481.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_213 & _T_719) begin
          $fatal; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@10482.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_213 & _T_723) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel AccessAck is corrupt (connected at SystemBus.scala:39:96)\n    at Monitor.scala:51 assert(cond, message)\n"); // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@10489.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_213 & _T_723) begin
          $fatal; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@10490.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_219 & _T_711) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel AccessAckData carries invalid source ID (connected at SystemBus.scala:39:96)\n    at Monitor.scala:51 assert(cond, message)\n"); // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@10508.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_219 & _T_711) begin
          $fatal; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@10509.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_219 & _T_719) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel AccessAckData carries invalid param (connected at SystemBus.scala:39:96)\n    at Monitor.scala:51 assert(cond, message)\n"); // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@10516.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_219 & _T_719) begin
          $fatal; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@10517.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_219 & _T_779) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel AccessAckData is denied but not corrupt (connected at SystemBus.scala:39:96)\n    at Monitor.scala:51 assert(cond, message)\n"); // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@10525.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_219 & _T_779) begin
          $fatal; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@10526.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_225 & _T_711) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel HintAck carries invalid source ID (connected at SystemBus.scala:39:96)\n    at Monitor.scala:51 assert(cond, message)\n"); // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@10544.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_225 & _T_711) begin
          $fatal; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@10545.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_225 & _T_719) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel HintAck carries invalid param (connected at SystemBus.scala:39:96)\n    at Monitor.scala:51 assert(cond, message)\n"); // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@10552.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_225 & _T_719) begin
          $fatal; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@10553.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_225 & _T_723) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel HintAck is corrupt (connected at SystemBus.scala:39:96)\n    at Monitor.scala:51 assert(cond, message)\n"); // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@10560.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_225 & _T_723) begin
          $fatal; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@10561.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_b_valid & _T_979) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel Probe carries unmanaged address (connected at SystemBus.scala:39:96)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@10750.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_b_valid & _T_979) begin
          $fatal; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@10751.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_b_valid & _T_985) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel Probe address not aligned to size (connected at SystemBus.scala:39:96)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@10764.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_b_valid & _T_985) begin
          $fatal; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@10765.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_b_valid & _T_989) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel Probe carries invalid cap param (connected at SystemBus.scala:39:96)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@10772.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_b_valid & _T_989) begin
          $fatal; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@10773.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_231 & _T_1220) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel ProbeAck carries unmanaged address (connected at SystemBus.scala:39:96)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@11199.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_231 & _T_1220) begin
          $fatal; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@11200.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_231 & _T_1223) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel ProbeAck carries invalid source ID (connected at SystemBus.scala:39:96)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@11206.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_231 & _T_1223) begin
          $fatal; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@11207.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_231 & _T_1227) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel ProbeAck smaller than a beat (connected at SystemBus.scala:39:96)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@11214.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_231 & _T_1227) begin
          $fatal; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@11215.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_231 & _T_1230) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel ProbeAck address not aligned to size (connected at SystemBus.scala:39:96)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@11221.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_231 & _T_1230) begin
          $fatal; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@11222.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_231 & _T_1234) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel ProbeAck carries invalid report param (connected at SystemBus.scala:39:96)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@11229.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_231 & _T_1234) begin
          $fatal; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@11230.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_231 & _T_1238) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel ProbeAck is corrupt (connected at SystemBus.scala:39:96)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@11237.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_231 & _T_1238) begin
          $fatal; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@11238.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_243 & _T_1220) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel ProbeAckData carries unmanaged address (connected at SystemBus.scala:39:96)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@11247.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_243 & _T_1220) begin
          $fatal; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@11248.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_243 & _T_1223) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel ProbeAckData carries invalid source ID (connected at SystemBus.scala:39:96)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@11254.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_243 & _T_1223) begin
          $fatal; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@11255.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_243 & _T_1227) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel ProbeAckData smaller than a beat (connected at SystemBus.scala:39:96)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@11262.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_243 & _T_1227) begin
          $fatal; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@11263.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_243 & _T_1230) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel ProbeAckData address not aligned to size (connected at SystemBus.scala:39:96)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@11269.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_243 & _T_1230) begin
          $fatal; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@11270.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_243 & _T_1234) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel ProbeAckData carries invalid report param (connected at SystemBus.scala:39:96)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@11277.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_243 & _T_1234) begin
          $fatal; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@11278.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_253 & _T_1309) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel carries Release type unsupported by manager (connected at SystemBus.scala:39:96)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@11336.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_253 & _T_1309) begin
          $fatal; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@11337.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_253 & _T_1323) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel carries Release from a client which does not support Probe (connected at SystemBus.scala:39:96)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@11359.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_253 & _T_1323) begin
          $fatal; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@11360.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_253 & _T_1223) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel Release carries invalid source ID (connected at SystemBus.scala:39:96)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@11366.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_253 & _T_1223) begin
          $fatal; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@11367.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_253 & _T_1227) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel Release smaller than a beat (connected at SystemBus.scala:39:96)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@11374.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_253 & _T_1227) begin
          $fatal; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@11375.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_253 & _T_1230) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel Release address not aligned to size (connected at SystemBus.scala:39:96)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@11381.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_253 & _T_1230) begin
          $fatal; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@11382.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_253 & _T_1337) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel Release carries invalid shrink param (connected at SystemBus.scala:39:96)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@11389.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_253 & _T_1337) begin
          $fatal; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@11390.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_253 & _T_1238) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel Release is corrupt (connected at SystemBus.scala:39:96)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@11397.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_253 & _T_1238) begin
          $fatal; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@11398.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_267 & _T_1309) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel carries ReleaseData type unsupported by manager (connected at SystemBus.scala:39:96)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@11456.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_267 & _T_1309) begin
          $fatal; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@11457.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_267 & _T_1323) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel carries Release from a client which does not support Probe (connected at SystemBus.scala:39:96)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@11479.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_267 & _T_1323) begin
          $fatal; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@11480.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_267 & _T_1223) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel ReleaseData carries invalid source ID (connected at SystemBus.scala:39:96)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@11486.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_267 & _T_1223) begin
          $fatal; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@11487.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_267 & _T_1227) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel ReleaseData smaller than a beat (connected at SystemBus.scala:39:96)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@11494.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_267 & _T_1227) begin
          $fatal; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@11495.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_267 & _T_1230) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel ReleaseData address not aligned to size (connected at SystemBus.scala:39:96)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@11501.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_267 & _T_1230) begin
          $fatal; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@11502.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_267 & _T_1337) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel ReleaseData carries invalid shrink param (connected at SystemBus.scala:39:96)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@11509.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_267 & _T_1337) begin
          $fatal; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@11510.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_279 & _T_1220) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel AccessAck carries unmanaged address (connected at SystemBus.scala:39:96)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@11519.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_279 & _T_1220) begin
          $fatal; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@11520.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_279 & _T_1223) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel AccessAck carries invalid source ID (connected at SystemBus.scala:39:96)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@11526.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_279 & _T_1223) begin
          $fatal; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@11527.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_279 & _T_1230) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel AccessAck address not aligned to size (connected at SystemBus.scala:39:96)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@11533.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_279 & _T_1230) begin
          $fatal; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@11534.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_279 & _T_1436) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel AccessAck carries invalid param (connected at SystemBus.scala:39:96)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@11541.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_279 & _T_1436) begin
          $fatal; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@11542.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_279 & _T_1238) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel AccessAck is corrupt (connected at SystemBus.scala:39:96)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@11549.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_279 & _T_1238) begin
          $fatal; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@11550.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_289 & _T_1220) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel AccessAckData carries unmanaged address (connected at SystemBus.scala:39:96)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@11559.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_289 & _T_1220) begin
          $fatal; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@11560.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_289 & _T_1223) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel AccessAckData carries invalid source ID (connected at SystemBus.scala:39:96)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@11566.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_289 & _T_1223) begin
          $fatal; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@11567.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_289 & _T_1230) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel AccessAckData address not aligned to size (connected at SystemBus.scala:39:96)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@11573.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_289 & _T_1230) begin
          $fatal; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@11574.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_289 & _T_1436) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel AccessAckData carries invalid param (connected at SystemBus.scala:39:96)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@11581.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_289 & _T_1436) begin
          $fatal; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@11582.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_297 & _T_1220) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel HintAck carries unmanaged address (connected at SystemBus.scala:39:96)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@11591.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_297 & _T_1220) begin
          $fatal; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@11592.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_297 & _T_1223) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel HintAck carries invalid source ID (connected at SystemBus.scala:39:96)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@11598.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_297 & _T_1223) begin
          $fatal; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@11599.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_297 & _T_1230) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel HintAck address not aligned to size (connected at SystemBus.scala:39:96)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@11605.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_297 & _T_1230) begin
          $fatal; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@11606.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_297 & _T_1436) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel HintAck carries invalid param (connected at SystemBus.scala:39:96)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@11613.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_297 & _T_1436) begin
          $fatal; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@11614.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_297 & _T_1238) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel HintAck is corrupt (connected at SystemBus.scala:39:96)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@11621.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_297 & _T_1238) begin
          $fatal; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@11622.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1503 & _T_1507) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel opcode changed within multibeat operation (connected at SystemBus.scala:39:96)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@11672.8]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_1503 & _T_1507) begin
          $fatal; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@11673.8]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1503 & _T_1511) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel param changed within multibeat operation (connected at SystemBus.scala:39:96)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@11680.8]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_1503 & _T_1511) begin
          $fatal; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@11681.8]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1503 & _T_1515) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel size changed within multibeat operation (connected at SystemBus.scala:39:96)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@11688.8]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_1503 & _T_1515) begin
          $fatal; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@11689.8]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1503 & _T_1519) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel source changed within multibeat operation (connected at SystemBus.scala:39:96)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@11696.8]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_1503 & _T_1519) begin
          $fatal; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@11697.8]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1503 & _T_1523) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel address changed with multibeat operation (connected at SystemBus.scala:39:96)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@11704.8]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_1503 & _T_1523) begin
          $fatal; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@11705.8]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1552 & _T_1556) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel opcode changed within multibeat operation (connected at SystemBus.scala:39:96)\n    at Monitor.scala:51 assert(cond, message)\n"); // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@11753.8]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_1552 & _T_1556) begin
          $fatal; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@11754.8]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1552 & _T_1560) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel param changed within multibeat operation (connected at SystemBus.scala:39:96)\n    at Monitor.scala:51 assert(cond, message)\n"); // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@11761.8]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_1552 & _T_1560) begin
          $fatal; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@11762.8]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1552 & _T_1564) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel size changed within multibeat operation (connected at SystemBus.scala:39:96)\n    at Monitor.scala:51 assert(cond, message)\n"); // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@11769.8]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_1552 & _T_1564) begin
          $fatal; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@11770.8]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1552 & _T_1568) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel source changed within multibeat operation (connected at SystemBus.scala:39:96)\n    at Monitor.scala:51 assert(cond, message)\n"); // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@11777.8]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_1552 & _T_1568) begin
          $fatal; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@11778.8]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1552 & _T_1572) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel sink changed with multibeat operation (connected at SystemBus.scala:39:96)\n    at Monitor.scala:51 assert(cond, message)\n"); // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@11785.8]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_1552 & _T_1572) begin
          $fatal; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@11786.8]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1552 & _T_1576) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel denied changed with multibeat operation (connected at SystemBus.scala:39:96)\n    at Monitor.scala:51 assert(cond, message)\n"); // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@11793.8]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_1552 & _T_1576) begin
          $fatal; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@11794.8]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1605 & _T_1613) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel param changed within multibeat operation (connected at SystemBus.scala:39:96)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@11851.8]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_1605 & _T_1613) begin
          $fatal; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@11852.8]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1605 & _T_1625) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel addresss changed with multibeat operation (connected at SystemBus.scala:39:96)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@11875.8]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_1605 & _T_1625) begin
          $fatal; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@11876.8]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1653 & _T_1657) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel opcode changed within multibeat operation (connected at SystemBus.scala:39:96)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@11923.8]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_1653 & _T_1657) begin
          $fatal; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@11924.8]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1653 & _T_1661) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel param changed within multibeat operation (connected at SystemBus.scala:39:96)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@11931.8]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_1653 & _T_1661) begin
          $fatal; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@11932.8]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1653 & _T_1665) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel size changed within multibeat operation (connected at SystemBus.scala:39:96)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@11939.8]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_1653 & _T_1665) begin
          $fatal; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@11940.8]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1653 & _T_1669) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel source changed within multibeat operation (connected at SystemBus.scala:39:96)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@11947.8]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_1653 & _T_1669) begin
          $fatal; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@11948.8]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1653 & _T_1673) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel address changed with multibeat operation (connected at SystemBus.scala:39:96)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@11955.8]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_1653 & _T_1673) begin
          $fatal; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@11956.8]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1732 & _T_1748) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel re-used a source ID (connected at SystemBus.scala:39:96)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@12091.8]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_1732 & _T_1748) begin
          $fatal; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@12092.8]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1771 & _T_1782) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel acknowledged for nothing inflight (connected at SystemBus.scala:39:96)\n    at Monitor.scala:51 assert(cond, message)\n"); // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@12142.8]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_1771 & _T_1782) begin
          $fatal; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@12143.8]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1771 & _T_1795) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel contains improper opcode response (connected at SystemBus.scala:39:96)\n    at Monitor.scala:51 assert(cond, message)\n"); // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@12159.8]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_1771 & _T_1795) begin
          $fatal; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@12160.8]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1771 & _T_1802) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel contains improper response size (connected at SystemBus.scala:39:96)\n    at Monitor.scala:51 assert(cond, message)\n"); // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@12170.8]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_1771 & _T_1802) begin
          $fatal; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@12171.8]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1809 & _T_1814) begin
          $fwrite(32'h80000002,"Assertion failed: ready check\n    at Monitor.scala:51 assert(cond, message)\n"); // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@12188.8]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_1809 & _T_1814) begin
          $fatal; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@12189.8]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1821) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' and 'D' concurrent, despite minlatency 1 (connected at SystemBus.scala:39:96)\n    at Monitor.scala:51 assert(cond, message)\n"); // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@12200.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_1821) begin
          $fatal; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@12201.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1840) begin
          $fwrite(32'h80000002,"Assertion failed: TileLink timeout expired (connected at SystemBus.scala:39:96)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@12228.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_1840) begin
          $fatal; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@12229.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1873 & _T_1880) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel re-used a sink ID (connected at SystemBus.scala:39:96)\n    at Monitor.scala:51 assert(cond, message)\n"); // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@12282.8]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_1873 & _T_1880) begin
          $fatal; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@12283.8]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_e_valid & _T_1891) begin
          $fwrite(32'h80000002,"Assertion failed: 'E' channel acknowledged for nothing inflight (connected at SystemBus.scala:39:96)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@12301.8]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_e_valid & _T_1891) begin
          $fatal; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@12302.8]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
  end
endmodule
